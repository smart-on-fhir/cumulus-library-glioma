#CUI|TUI|TTY|CODE|SAB|STR|PREF
C1370507|T191|SY|0000021045|CHV|cerebellar liponeurocytoma|0000/0
C2347979|T191|ET|HP:0025171|HPO|Rosette-forming glioneuronal tumor of the fourth ventricle|0000/0
C1370507|T191|PN|NOCODE|MTH|Cerebellar Liponeurocytoma|0000/0
C1370507|T191|PT|C6905|NCI|Cerebellar Liponeurocytoma|0000/0
C1370507|T191|SY|C6905|NCI|Lipomatous Medulloblastoma|0000/0
C1513719|T191|PT|C39807|NCI|Mucinous Tubular and Spindle Cell Carcinoma of the Kidney|0000/0
C1337036|T191|PT|C27891|NCI|Renal Cell Carcinoma Associated with Xp11.2 Translocations/TFE3 Gene Fusions|0000/0
C2347979|T191|PT|C67559|NCI|Rosette-Forming Glioneuronal Tumor of the Fourth Ventricle|0000/0
C1337036|T191|SY|C27891|NCI|TFE3-Rearranged Renal Cell Carcinoma|0000/0
C1337036|T191|AB|C27891|NCI|tRCC|0000/0
C1337036|T191|SY|C27891|NCI|Xp11.2 Translocation-Related Renal Cell Carcinoma|0000/0
C1513719|T191|PT|C39807|NCI_CDISC|CARCINOMA, RENAL, TUBULAR, MALIGNANT|0000/0
C1513719|T191|SY|C39807|NCI_CDISC|Mucinous Tubular and Spindle Cell Carcinoma of the Kidney|0000/0
C1337036|T191|DN|C27891|NCI_CTRP|Renal Cell Cancer Associated with Xp11.2 Translocations/TFE3 Gene Fusions|0000/0
C1370507|T191|IS|128858006|SNOMEDCT_US|Cerebellar liponeurocytoma|0000/0
C1370507|T191|PT|734134003|SNOMEDCT_US|Cerebellar liponeurocytoma|0000/0
C1370507|T191|PT|716592003|SNOMEDCT_US|Cerebellar liponeurocytoma|0000/0
C1370507|T191|SY|716592003|SNOMEDCT_US|Liponeurocytoma of cerebellum|0000/0
C0086692|T191|PT|0061294|CCPSS|NEOPLASM BENIGN NOS|8000/0
C0086692|T191|MD|2.16|CCS|Benign neoplasms|8000/0
C0086692|T191|SD|NEO073|CCSR_10|Benign neoplasms|8000/0
C0086692|T191|SY|0000015985|CHV|benign neoplasm|8000/0
C0086692|T191|SY|0000015985|CHV|benign neoplasms|8000/0
C0086692|T191|PT|0000015985|CHV|benign tumor|8000/0
C0086692|T191|SY|0000015985|CHV|benign tumors|8000/0
C0086692|T191|SY|0000015985|CHV|benign tumour|8000/0
C0086692|T191|SY|0000015985|CHV|benign tumours|8000/0
C0086692|T191|SY|0000015985|CHV|nonmalignant tumor|8000/0
C0086692|T191|SY|0000015985|CHV|nonmalignant tumors|8000/0
C0086692|T191|PT|U000008|COSTAR|BENIGN TUMOR|8000/0
C0086692|T191|HT|PATHTUMORBEN|CST|NONMALIGNANT TUMORS|8000/0
C0086692|T191|PT|D36.9|ICD10|Benign neoplasm of unspecified site|8000/0
C0086692|T191|HT|D10-D36.9|ICD10|Benign neoplasms|8000/0
C0086692|T191|AB|D36.9|ICD10CM|Benign neoplasm, unspecified site|8000/0
C0086692|T191|PT|D36.9|ICD10CM|Benign neoplasm, unspecified site|8000/0
C0086692|T191|AB|229.9|ICD9CM|Benign neoplasm NOS|8000/0
C0086692|T191|PT|229.9|ICD9CM|Benign neoplasm of unspecified site|8000/0
C0086692|T191|HT|210-229.99|ICD9CM|BENIGN NEOPLASMS|8000/0
C0086692|T191|PTN|A99018|ICPC2P|benign neoplasm of unspecified site|8000/0
C0086692|T191|PT|A99018|ICPC2P|Neoplasm benign;site unspecifi|8000/0
C0086692|T191|LLT|10060999|MDR|Benign neoplasm|8000/0
C0086692|T191|PT|10060999|MDR|Benign neoplasm|8000/0
C0086692|T191|LLT|10004299|MDR|Benign neoplasm NOS|8000/0
C0086692|T191|LLT|10004417|MDR|Benign neoplasm of unspecified site|8000/0
C0086692|T191|PT|98330|MEDCIN|benign neoplasm|8000/0
C0086692|T191|PT|3585|MEDLINEPLUS|Benign Tumors|8000/0
C0086692|T191|SY|3585|MEDLINEPLUS|Noncancerous tumors|8000/0
C0086692|T191|ET|3585|MEDLINEPLUS|Tumors, Benign|8000/0
C0086692|T191|DEV|D009369|MSH|BENIGN NEOPL|8000/0
C0086692|T191|PM|D009369|MSH|Benign Neoplasm|8000/0
C0086692|T191|PEP|D009369|MSH|Benign Neoplasms|8000/0
C0086692|T191|DEV|D009369|MSH|NEOPL BENIGN|8000/0
C0086692|T191|PM|D009369|MSH|Neoplasm, Benign|8000/0
C0086692|T191|ET|D009369|MSH|Neoplasms, Benign|8000/0
C0086692|T191|PN|NOCODE|MTH|Benign Neoplasm|8000/0
C0086692|T191|PT|C3677|NCI|Benign Neoplasm|8000/0
C0086692|T191|SY|C3677|NCI|Benign Tumor|8000/0
C0086692|T191|SY|C3677|NCI_CDISC|Benign Tumor|8000/0
C0086692|T191|SY|C3677|NCI_CDISC|Benign Unclassifiable Tumor|8000/0
C0086692|T191|PT|C3677|NCI_CDISC|NEOPLASM, BENIGN|8000/0
C0086692|T191|PT|C3677|NCI_CPTAC|Benign Neoplasm|8000/0
C0086692|T191|DN|C3677|NCI_CTRP|Benign Neoplasm|8000/0
C0086692|T191|PT|CDR0000046079|NCI_NCI-GLOSS|benign tumor|8000/0
C0086692|T191|SY|CDR0000664287|PDQ|benign neoplasm|8000/0
C0086692|T191|ET|CDR0000664287|PDQ|Benign tumor or blood disorder|8000/0
C0086692|T191|PT|CDR0000664287|PDQ|nonmalignant neoplasm|8000/0
C0086692|T191|PT|05800|PSY|Benign Neoplasms|8000/0
C0086692|T191|SY|B7...|RCD|Benign neoplasm|8000/0
C0086692|T191|OP|B7zz.|RCD|Benign neoplasm NOS|8000/0
C0086692|T191|PT|B7...|RCD|Benign tumour|8000/0
C0086692|T191|PT|BB00.|RCD|Benign tumour morphology|8000/0
C0086692|T191|PT|B7...|RCDAE|Benign tumor|8000/0
C0086692|T191|PT|BB00.|RCDAE|Benign tumor morphology|8000/0
C0086692|T191|OP|ByuG.|RCDSY|Benign neoplasms|8000/0
C0086692|T191|SY|3898006|SNOMEDCT_US|Benign neoplasm|8000/0
C0086692|T191|OF|154633007|SNOMEDCT_US|Benign neoplasm NOS|8000/0
C0086692|T191|OAP|154633007|SNOMEDCT_US|Benign neoplasm NOS|8000/0
C0086692|T191|OAP|189207002|SNOMEDCT_US|Benign neoplasm NOS|8000/0
C0086692|T191|SY|3898006|SNOMEDCT_US|Benign neoplasm, site unspecified|8000/0
C0086692|T191|PT|20376005|SNOMEDCT_US|Benign neoplastic disease|8000/0
C0086692|T191|OAP|154607004|SNOMEDCT_US|Benign tumor|8000/0
C0086692|T191|SY|3898006|SNOMEDCT_US|Benign tumor morphology|8000/0
C0086692|T191|OAP|154607004|SNOMEDCT_US|Benign tumour|8000/0
C0086692|T191|OF|154607004|SNOMEDCT_US|Benign tumour|8000/0
C0086692|T191|SYGB|3898006|SNOMEDCT_US|Benign tumour morphology|8000/0
C0086692|T191|PT|3898006|SNOMEDCT_US|Neoplasm, benign|8000/0
C0086692|T191|SY|3898006|SNOMEDCT_US|Tumor, benign|8000/0
C0086692|T191|SYGB|3898006|SNOMEDCT_US|Tumour, benign|8000/0
C0086692|T191|SY|3898006|SNOMEDCT_US|Unclassified tumor, benign|8000/0
C0086692|T191|SYGB|3898006|SNOMEDCT_US|Unclassified tumour, benign|8000/0
C0677041|T191|SY|0000042588|CHV|borderline malignancy tumor|8000/1
C0677041|T191|PT|0000042588|CHV|uncertain whether benign or malignant neoplasm|8000/1
C0677041|T191|PN|NOCODE|MTH|Neoplasm, uncertain whether benign or malignant|8000/1
C0677041|T191|HD|C65157|NCI|Neoplasm, Uncertain Whether Benign or Malignant|8000/1
C0677041|T191|PT|C65157|NCI|Neoplasm, Uncertain Whether Benign or Malignant|8000/1
C0677041|T191|PT|C65157|NCI_CPTAC|Neoplasm, Uncertain Whether Benign or Malignant|8000/1
C0677041|T191|OA|BB01.|RCDSY|Neoplasm, ?benign or malig|8000/1
C0677041|T191|OP|BB01.|RCDSY|Neoplasm, uncertain whether benign or malignant|8000/1
C1302828|T191|PT|400095002|SNOMEDCT_US|Blood vessel neoplasm, uncertain whether benign or malignant|8000/1
C1533006|T191|PTGB|414389009|SNOMEDCT_US|Haematopoietic neoplasm of uncertain behaviour|8000/1
C1533006|T191|PT|414389009|SNOMEDCT_US|Hematopoietic neoplasm of uncertain behavior|8000/1
C5190876|T191|PT|783219005|SNOMEDCT_US|Melanocytic tumor of uncertain malignant potential|8000/1
C5190876|T191|PTGB|783219005|SNOMEDCT_US|Melanocytic tumour of uncertain malignant potential|8000/1
C5190876|T191|SY|783219005|SNOMEDCT_US|MELTUMP - melanocytic tumor of uncertain malignant potential|8000/1
C5190876|T191|SYGB|783219005|SNOMEDCT_US|MELTUMP - melanocytic tumour of uncertain malignant potential|8000/1
C0677041|T191|PT|86251006|SNOMEDCT_US|Neoplasm, uncertain whether benign or malignant|8000/1
C0677041|T191|SY|86251006|SNOMEDCT_US|Tumor, borderline malignancy|8000/1
C0677041|T191|SY|86251006|SNOMEDCT_US|Tumor, uncertain whether benign or malignant|8000/1
C0677041|T191|SYGB|86251006|SNOMEDCT_US|Tumour, borderline malignancy|8000/1
C0677041|T191|SYGB|86251006|SNOMEDCT_US|Tumour, uncertain whether benign or malignant|8000/1
C0677041|T191|SY|86251006|SNOMEDCT_US|Unclassified tumor, borderline malignancy|8000/1
C0677041|T191|IS|86251006|SNOMEDCT_US|Unclassified tumor, uncertain whether benign or malignant|8000/1
C0677041|T191|SYGB|86251006|SNOMEDCT_US|Unclassified tumour, borderline malignancy|8000/1
C0006826|T191|DE|0000004520|AOD|cancer|8000/3
C0006826|T191|NP|0000023015|AOD|malignant neoplasm|8000/3
C0006826|T191|NP|0000023016|AOD|malignant tumor|8000/3
C0006826|T191|NP|0000023014|AOD|malignant tumoral disease|8000/3
C0006826|T191|PT|BI00731|BI|malignancies|8000/3
C0006826|T191|PT|1001968|CCPSS|CANCER|8000/3
C0006826|T191|PT|1017904|CCPSS|MALIGNANCY|8000/3
C0006826|T191|MD|2.13|CCS|Malignant neoplasm without specification of site|8000/3
C0006826|T191|SD|43|CCS|Malignant neoplasm without specification of site|8000/3
C0006826|T191|PT|0000002337|CHV|cancer|8000/3
C0006826|T191|SY|0000002337|CHV|cancers|8000/3
C0006826|T191|SY|0000002337|CHV|malignancies|8000/3
C0006826|T191|SY|0000002337|CHV|malignant neoplasm|8000/3
C1306459|T191|SY|0000052870|CHV|malignant neoplasm|8000/3
C0006826|T191|SY|0000002337|CHV|malignant neoplasms|8000/3
C0006826|T191|SY|0000002337|CHV|malignant tumor|8000/3
C0006826|T191|SY|0000002337|CHV|malignant tumors|8000/3
C0006826|T191|SY|0000002337|CHV|malignant tumour|8000/3
C0006826|T191|SY|0000002337|CHV|malignant tumours|8000/3
C1306459|T191|PT|0000052870|CHV|primary cancer|8000/3
C0006826|T191|PT|465|COSTAR|MALIGNANCY|8000/3
C0006826|T191|PT|U000036|COSTAR|MALIGNANT TUMOR|8000/3
C0006826|T191|ET|2000-0173|CSP|cancer|8000/3
C0006826|T191|PT|2000-0173|CSP|neoplasm/cancer|8000/3
C0006826|T191|GT|CARCINOMA|CST|CANCER|8000/3
C0006826|T191|HT|PATHMALIGN|CST|MALIGNANCIES|8000/3
C0006826|T191|HT|RETICMALIG|CST|MALIGNANCY|8000/3
C0006826|T191|GT|CARCINOMA|CST|NEOPLASM MALIGNANT|8000/3
C0006826|T191|FI|U000537|DXP|CANCER|8000/3
C0006826|T191|ET|HP:0002664|HPO|Cancer|8000/3
C0006826|T191|PT|C80|ICD10|Malignant neoplasm without specification of site|8000/3
C0006826|T191|HT|C00-C97.9|ICD10|Malignant neoplasms|8000/3
C0006826|T191|ET|C80.1|ICD10CM|Cancer NOS|8000/3
C0006826|T191|AB|C80|ICD10CM|Malignant neoplasm without specification of site|8000/3
C0006826|T191|HT|C80|ICD10CM|Malignant neoplasm without specification of site|8000/3
C0006826|T191|HT|199|ICD9CM|Malignant neoplasm without specification of site|8000/3
C0006826|T191|PT|A79|ICPC2EENG|Malignancy nos|8000/3
C0006826|T191|AB|A79|ICPC2EENG|Malignancy nos|8000/3
C0006826|T191|PT|MTHU077094|ICPC2ICD10ENG|tumor; malignant, unclassified|8000/3
C0006826|T191|PT|MTHU077120|ICPC2ICD10ENG|tumor; unclassified, malignant|8000/3
C0006826|T191|PTN|A79001|ICPC2P|cancer|8000/3
C0006826|T191|PT|A79001|ICPC2P|Cancer|8000/3
C0006826|T191|PT|U006339|LCH|Cancer|8000/3
C0006826|T191|PT|sh85019492|LCH_NW|Cancer|8000/3
C0006826|T191|LPN|LP281735-3|LNC|^Cancer|8000/3
C0006826|T191|CN|MTHU010328|LNC|Cancer|8000/3
C0006826|T191|LPN|LP100805-3|LNC|Cancer|8000/3
C0006826|T191|LPN|LP7106-0|LNC|Cancer|8000/3
C0006826|T191|LA|LA10524-9|LNC|Cancer|8000/3
C0006826|T191|LS|MTHU051589|LNC|Cancer|8000/3
C0006826|T191|CN|MTHU040703|LNC|Malignancy|8000/3
C0006826|T191|LPN|LP20701-6|LNC|Malignancy|8000/3
C0006826|T191|LPN|LP128794-7|LNC|Malignancy|8000/3
C0006826|T191|LA|LA25513-5|LNC|Malignant neoplasm|8000/3
C0006826|T191|LLT|10007050|MDR|Cancer|8000/3
C0006826|T191|LLT|10025691|MDR|Malignant neoplasm NOS|8000/3
C0006826|T191|LLT|10026655|MDR|Malignant neoplasm without specification of site|8000/3
C0006826|T191|LLT|10049516|MDR|Malignant tumor|8000/3
C0006826|T191|LLT|10073835|MDR|Malignant tumour|8000/3
C0006826|T191|LLT|10028997|MDR|Neoplasm malignant|8000/3
C0006826|T191|PT|10028997|MDR|Neoplasm malignant|8000/3
C1306459|T191|LLT|10078954|MDR|Primary malignant neoplasm|8000/3
C0006826|T191|PT|31465|MEDCIN|cancer|8000/3
C0006826|T191|SY|31465|MEDCIN|cancer, NOS|8000/3
C0006826|T191|PT|99725|MEDCIN|malignant neoplasm|8000/3
C1306459|T191|SY|339753|MEDCIN|malignant neoplasm primary|8000/3
C1306459|T191|PT|339753|MEDCIN|Primary malignant neoplasm|8000/3
C0006826|T191|PT|25|MEDLINEPLUS|Cancer|8000/3
C0006826|T191|HT|1|MEDLINEPLUS|Cancers|8000/3
C0006826|T191|ET|25|MEDLINEPLUS|Malignancy|8000/3
C0006826|T191|SY|25|MEDLINEPLUS|Malignancy|8000/3
C0006826|T191|PEP|D009369|MSH|Cancer|8000/3
C0006826|T191|PM|D009369|MSH|Cancers|8000/3
C0006826|T191|PM|D009369|MSH|Malignancies|8000/3
C0006826|T191|ET|D009369|MSH|Malignancy|8000/3
C0006826|T191|PM|D009369|MSH|Malignant Neoplasm|8000/3
C0006826|T191|ET|D009369|MSH|Malignant Neoplasms|8000/3
C0006826|T191|PM|D009369|MSH|Neoplasm, Malignant|8000/3
C0006826|T191|PM|D009369|MSH|Neoplasms, Malignant|8000/3
C0006826|T191|PN|NOCODE|MTH|Malignant Neoplasms|8000/3
C1306459|T191|PN|NOCODE|MTH|Primary malignant neoplasm|8000/3
C0006826|T191|ET|199.1|MTHICD9|Cancer, unspecified site|8000/3
C0006826|T191|ET|199.1|MTHICD9|Malignancy, unspecified site|8000/3
C0006826|T191|RT|01968|NANDA-I|Cancer|8000/3
C0006826|T191|AB|C9305|NCI|CA|8000/3
C0006826|T191|SY|C9305|NCI|Cancer|8000/3
C0006826|T191|SY|C9305|NCI|Malignancy|8000/3
C0006826|T191|SY|NHIS|NCI|Malignant Neoplasm|8000/3
C0006826|T191|PT|C9305|NCI|Malignant Neoplasm|8000/3
C0006826|T191|SY|TCGA|NCI|Malignant Neoplasm|8000/3
C0006826|T191|SY|C9305|NCI|Malignant Tumor|8000/3
C1306459|T191|PT|C84509|NCI|Primary Malignant Neoplasm|8000/3
C0006826|T191|SY|C9305|NCI_CDISC|CA|8000/3
C0006826|T191|SY|C9305|NCI_CDISC|Cancer|8000/3
C0006826|T191|SY|C9305|NCI_CDISC|Malignancy|8000/3
C0006826|T191|SY|C9305|NCI_CDISC|Malignant Tumor|8000/3
C0006826|T191|PT|C9305|NCI_CDISC|NEOPLASM, MALIGNANT|8000/3
C0006826|T191|PT|C9305|NCI_CPTAC|Malignant Neoplasm|8000/3
C1306459|T191|PT|C84509|NCI_CPTAC|Primary Malignant Neoplasm|8000/3
C0006826|T191|DN|C9305|NCI_CTRP|Malignant Neoplasm|8000/3
C0006826|T191|PT|3262|NCI_FDA|Cancer|8000/3
C0006826|T191|SY|3262|NCI_FDA|Malignant Neoplasm|8000/3
C0006826|T191|PT|CDR0000045333|NCI_NCI-GLOSS|cancer|8000/3
C0006826|T191|PT|CDR0000045771|NCI_NCI-GLOSS|malignancy|8000/3
C0006826|T191|PT|C9305|NCI_NICHD|Cancer|8000/3
C0006826|T191|SY|C9305|NCI_NICHD|Malignancy|8000/3
C0006826|T191|SY|C9305|NCI_NICHD|Malignant Growth|8000/3
C0006826|T191|SY|C9305|NCI_NICHD|Malignant Neoplasm|8000/3
C0006826|T191|SY|C9305|NCI_NICHD|Malignant Neoplastic Disease|8000/3
C0006826|T191|AB|CDR0000041060|PDQ|CA|8000/3
C0006826|T191|SY|CDR0000041060|PDQ|Cancer|8000/3
C0006826|T191|SY|CDR0000041060|PDQ|Malignancy|8000/3
C0006826|T191|PT|CDR0000041060|PDQ|malignant neoplasm|8000/3
C0006826|T191|SY|CDR0000041060|PDQ|Malignant Tumor|8000/3
C0006826|T191|ET|07420|PSY|Cancers|8000/3
C0006826|T191|ET|29280|PSY|Malignant Neoplasms|8000/3
C0006826|T191|SY|X78ef|RCD|CA - Cancer|8000/3
C0006826|T191|OP|XE20H|RCD|Ca - unspecified site NOS|8000/3
C0006826|T191|SY|X78ef|RCD|Cancer|8000/3
C1306459|T191|SY|BB02.|RCD|Cancer morphology|8000/3
C0006826|T191|OA|B59..|RCD|Malig neop of unspec site|8000/3
C0006826|T191|OA|B59z.|RCD|Malig neop of unspec site NOS|8000/3
C1306459|T191|SY|BB02.|RCD|Malignancy|8000/3
C0006826|T191|SY|X78ef|RCD|Malignant neoplasm|8000/3
C0006826|T191|OP|B59..|RCD|Malignant neoplasm of unspecified site|8000/3
C0006826|T191|OP|B59z.|RCD|Malignant neoplasm of unspecified site NOS|8000/3
C0006826|T191|PT|X78ef|RCD|Malignant tumour|8000/3
C1306459|T191|PT|BB02.|RCD|Malignant tumour morphology|8000/3
C0006826|T191|PT|X78ef|RCDAE|Malignant tumor|8000/3
C1306459|T191|PT|BB02.|RCDAE|Malignant tumor morphology|8000/3
C0006826|T191|OA|ByuC8|RCDSY|Mal neo w'out specfctn/site|8000/3
C0006826|T191|OP|ByuC8|RCDSY|Malignant neoplasm without specification of site|8000/3
C0006826|T191|SY|363346000|SNOMEDCT_US|CA - Cancer|8000/3
C0006826|T191|OAS|38807002|SNOMEDCT_US|CA - Cancer|8000/3
C0006826|T191|OAS|269623003|SNOMEDCT_US|Ca - unspecified site|8000/3
C0006826|T191|OAP|154577008|SNOMEDCT_US|Ca - unspecified site NOS|8000/3
C0006826|T191|OAP|269626006|SNOMEDCT_US|Ca - unspecified site NOS|8000/3
C0006826|T191|OF|154577008|SNOMEDCT_US|Ca - unspecified site NOS|8000/3
C0006826|T191|OAS|38807002|SNOMEDCT_US|Cancer|8000/3
C0006826|T191|SY|363346000|SNOMEDCT_US|Cancer|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Cancer|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Cancer morphology|8000/3
C0006826|T191|OAS|187597000|SNOMEDCT_US|Cancers|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Malignancy|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Malignant neoplasm|8000/3
C0006826|T191|SY|363346000|SNOMEDCT_US|Malignant neoplasm|8000/3
C0006826|T191|OAS|38807002|SNOMEDCT_US|Malignant neoplasm|8000/3
C0006826|T191|OAS|269634000|SNOMEDCT_US|Malignant neoplasm NOS|8000/3
C0006826|T191|OAP|188475001|SNOMEDCT_US|Malignant neoplasm of unspecified site|8000/3
C0006826|T191|OAP|188482002|SNOMEDCT_US|Malignant neoplasm of unspecified site NOS|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Malignant neoplasm, primary|8000/3
C0006826|T191|OAS|269513004|SNOMEDCT_US|Malignant neoplasms|8000/3
C0006826|T191|OAS|154433003|SNOMEDCT_US|Malignant neoplasms|8000/3
C0006826|T191|IS|38807002|SNOMEDCT_US|Malignant neoplastic disease|8000/3
C0006826|T191|PT|363346000|SNOMEDCT_US|Malignant neoplastic disease|8000/3
C0006826|T191|OAP|154432008|SNOMEDCT_US|Malignant tumor|8000/3
C0006826|T191|SY|363346000|SNOMEDCT_US|Malignant tumor|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Malignant tumor morphology|8000/3
C0006826|T191|SYGB|363346000|SNOMEDCT_US|Malignant tumour|8000/3
C0006826|T191|OAP|154432008|SNOMEDCT_US|Malignant tumour|8000/3
C0006826|T191|OF|154432008|SNOMEDCT_US|Malignant tumour|8000/3
C1306459|T191|SYGB|86049000|SNOMEDCT_US|Malignant tumour morphology|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Neoplasm, malignant|8000/3
C0006826|T191|OAS|269513004|SNOMEDCT_US|Neoplasms - malignant|8000/3
C0006826|T191|OAS|154433003|SNOMEDCT_US|Neoplasms - malignant|8000/3
C1306459|T191|PT|372087000|SNOMEDCT_US|Primary malignant neoplasm|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Tumor, malignant|8000/3
C1306459|T191|IS|86049000|SNOMEDCT_US|Tumor, malignant, NOS|8000/3
C1306459|T191|SYGB|86049000|SNOMEDCT_US|Tumour, malignant|8000/3
C1306459|T191|SY|86049000|SNOMEDCT_US|Unclassified tumor, malignant|8000/3
C1306459|T191|SYGB|86049000|SNOMEDCT_US|Unclassified tumour, malignant|8000/3
C0006826|T191|PT|1345|WHO|NEOPLASM MALIGNANT|8000/3
C2939419|T191|PT|1017407|CCPSS|CANCER METASTATIC|8000/6
C2939420|T191|PT|0025094|CCPSS|METASTATIC DISEASE|8000/6
C2939419|T191|MD|2.12|CCS|Secondary malignancies|8000/6
C2939419|T191|SD|42|CCS|Secondary malignancies|8000/6
C2939419|T191|SD|NEO070|CCSR_10|Secondary malignancies|8000/6
C2939419|T191|SY|0000015723|CHV|secondary neoplasm|8000/6
C2939420|T191|ET|C79.9|ICD10CM|Metastatic cancer NOS|8000/6
C2939420|T191|ET|C79.9|ICD10CM|Metastatic disease NOS|8000/6
C2939419|T191|PT|MTHU040813|ICPC2ICD10ENG|cancer; metastatic|8000/6
C2939419|T191|PT|MTHU049030|ICPC2ICD10ENG|metastatic; cancer or neoplasm|8000/6
C2939419|T191|PT|MTHU052245|ICPC2ICD10ENG|neoplasm; metastatic|8000/6
C2939420|T191|LA|LA28289-9|LNC|Metastatic cancer|8000/6
C2939420|T191|LLT|10027478|MDR|Metastatic disease|8000/6
C2939419|T191|LLT|10061289|MDR|Metastatic neoplasm|8000/6
C2939419|T191|PT|10061289|MDR|Metastatic neoplasm|8000/6
C2939420|T191|PT|31778|MEDCIN|metastasis from malignant neoplasm|8000/6
C2939420|T191|SY|31778|MEDCIN|metastatic cancer|8000/6
C2939420|T191|PN|NOCODE|MTH|Metastatic Neoplasm|8000/6
C2939419|T191|PN|NOCODE|MTH|Secondary Neoplasm|8000/6
C2939419|T191|SY|C36263|NCI|Metastatic Cancer|8000/6
C2939420|T191|SY|C3261|NCI|Metastatic Disease|8000/6
C2939419|T191|PT|C36263|NCI|Metastatic Malignant Neoplasm|8000/6
C2939420|T191|PT|C3261|NCI|Metastatic Neoplasm|8000/6
C2939420|T191|SY|TCGA|NCI|Metastatic Neoplasm|8000/6
C2939420|T191|SY|C3261|NCI|Metastatic Tumor|8000/6
C2939419|T191|PT|C36255|NCI|Secondary Neoplasm|8000/6
C2939419|T191|SY|C36255|NCI|Secondary Tumor|8000/6
C2939419|T191|PT|C36263|NCI_CPTAC|Metastatic Malignant Neoplasm|8000/6
C2939419|T191|DN|C36263|NCI_CTRP|Metastatic Malignant Neoplasm|8000/6
C2939419|T191|PT|CDR0000045951|NCI_NCI-GLOSS|secondary tumor|8000/6
C2939420|T191|SY|CDR0000041702|PDQ|cancer, metastatic|8000/6
C2939420|T191|ET|CDR0000041702|PDQ|Metastatic cancer|8000/6
C2939420|T191|PT|CDR0000041702|PDQ|metastatic cancer|8000/6
C2939420|T191|SY|CDR0000041687|PDQ|metastatic disease|8000/6
C2939420|T191|SY|CDR0000041702|PDQ|Metastatic Malignant Neoplasm|8000/6
C2939420|T191|PSC|CDR0000041687|PDQ|metastatic neoplasm|8000/6
C2939420|T191|SY|CDR0000041687|PDQ|metastatic tumor|8000/6
C2939419|T191|SY|Xa982|RCD|CA - Secondary cancer|8000/6
C2939419|T191|SY|Xa982|RCD|Metastases|8000/6
C2939419|T191|SY|Xa983|RCD|Metastatic cancer|8000/6
C2939419|T191|PT|Xa982|RCD|Metastatic malignant disease|8000/6
C2939419|T191|SY|Xa982|RCD|Metastatic neoplasm|8000/6
C2939419|T191|SY|Xa982|RCD|Secondaries|8000/6
C2939419|T191|OP|XE20B|RCD|Secondary Ca NOS|8000/6
C2939419|T191|SY|Xa982|RCD|Secondary cancer|8000/6
C2939419|T191|SY|Xa982|RCD|Secondary malignant deposit|8000/6
C2939419|T191|SY|XM1GJ|RCD|Secondary neoplasm|8000/6
C2939419|T191|SY|Xa982|RCD|Secondary tumour|8000/6
C2939419|T191|SY|Xa982|RCD|Tumour metastasis|8000/6
C2939419|T191|SY|Xa982|RCDAE|Secondary tumor|8000/6
C2939419|T191|SY|Xa982|RCDAE|Tumor metastasis|8000/6
C2939419|T191|OP|XE1wR|RCDSY|Neoplasm, metastatic|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|CA - Secondary cancer|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Metastases|8000/6
C2939419|T191|OAS|302818005|SNOMEDCT_US|Metastatic cancer|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Metastatic cancer|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Metastatic malignant disease|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Metastatic neoplasm|8000/6
C2939419|T191|PT|14799000|SNOMEDCT_US|Neoplasm, metastatic|8000/6
C2939419|T191|SY|14799000|SNOMEDCT_US|Neoplasm, secondary|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Secondaries|8000/6
C2939419|T191|OF|154574001|SNOMEDCT_US|Secondary Ca NOS|8000/6
C2939419|T191|OAP|154574001|SNOMEDCT_US|Secondary Ca NOS|8000/6
C2939419|T191|OAP|269622008|SNOMEDCT_US|Secondary Ca NOS|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Secondary cancer|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Secondary malignant deposit|8000/6
C2939419|T191|PT|128462008|SNOMEDCT_US|Secondary malignant neoplastic disease|8000/6
C2939419|T191|SY|79282002|SNOMEDCT_US|Secondary neoplasm|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Secondary tumor|8000/6
C2939419|T191|SYGB|128462008|SNOMEDCT_US|Secondary tumour|8000/6
C2939419|T191|SY|128462008|SNOMEDCT_US|Tumor metastasis|8000/6
C2939419|T191|SY|14799000|SNOMEDCT_US|Tumor, metastatic|8000/6
C2939419|T191|SY|14799000|SNOMEDCT_US|Tumor, secondary|8000/6
C2939419|T191|SYGB|128462008|SNOMEDCT_US|Tumour metastasis|8000/6
C2939419|T191|SYGB|14799000|SNOMEDCT_US|Tumour, metastatic|8000/6
C2939419|T191|SYGB|14799000|SNOMEDCT_US|Tumour, secondary|8000/6
C0334224|T191|PT|C65153|NCI|Malignant Neoplasm, Uncertain Whether Primary or Metastatic|8000/9
C0334224|T191|PT|C65153|NCI_CPTAC|Malignant Neoplasm, Uncertain Whether Primary or Metastatic|8000/9
C0334224|T191|AB|BB04.|RCD|Mal tumour-uncert prim/metast|8000/9
C0334224|T191|PT|BB04.|RCD|Malignant tumour - uncertain whether primary or metastatic|8000/9
C0334224|T191|AB|BB04.|RCDAE|Mal tumor-uncert prim/metast|8000/9
C0334224|T191|PT|BB04.|RCDAE|Malignant tumor - uncertain whether primary or metastatic|8000/9
C0334224|T191|SY|6219000|SNOMEDCT_US|Malignant tumor - uncertain whether primary or metastatic|8000/9
C0334224|T191|SYGB|6219000|SNOMEDCT_US|Malignant tumour - uncertain whether primary or metastatic|8000/9
C0334224|T191|PT|6219000|SNOMEDCT_US|Neoplasm, malignant, uncertain whether primary or metastatic|8000/9
C0334224|T191|SY|6219000|SNOMEDCT_US|Unclassified tumor, malignant, uncertain whether primary or metastatic|8000/9
C0334224|T191|SYGB|6219000|SNOMEDCT_US|Unclassified tumour, malignant, uncertain whether primary or metastatic|8000/9
C0334225|T025|SY|0000029939|CHV|benign cells tumor|8001/0
C0334225|T025|PT|0000029939|CHV|benign tumor cells|8001/0
C0334225|T025|SY|0000029939|CHV|cell tumor benign|8001/0
C0334225|T025|PT|BB05.|RCD|Benign tumour cells|8001/0
C0334225|T025|PT|BB05.|RCDAE|Benign tumor cells|8001/0
C0334225|T025|SY|56696000|SNOMEDCT_US|Benign tumor cells|8001/0
C0334225|T025|SYGB|56696000|SNOMEDCT_US|Benign tumour cells|8001/0
C0334225|T025|PT|56696000|SNOMEDCT_US|Tumor cells, benign|8001/0
C0334225|T025|PTGB|56696000|SNOMEDCT_US|Tumour cells, benign|8001/0
C0431085|T025|PT|0000034147|CHV|tumor cell|8001/1
C0431085|T025|SY|0000034147|CHV|tumor cells|8001/1
C0431085|T025|SY|0000034147|CHV|tumour cell|8001/1
C0431085|T025|SY|0000034147|CHV|tumour cells|8001/1
C0431085|T025|PN|NOCODE|MTH|Tumor cells, uncertain whether benign or malignant|8001/1
C0431085|T025|PT|X77mt|RCD|Tumour cells|8001/1
C0431085|T025|PT|X77mt|RCDAE|Tumor cells|8001/1
C0431085|T025|OP|BB06.|RCDSA|Tumor cells, uncertain whether benign or malignant|8001/1
C0431085|T025|OA|BB06.|RCDSA|Tumor cells,?benign/?malig|8001/1
C0431085|T025|OP|BB0z.|RCDSA|Unspecified tumor cell NOS|8001/1
C0431085|T025|OP|BB06.|RCDSY|Tumour cells, uncertain whether benign or malignant|8001/1
C0431085|T025|OA|BB06.|RCDSY|Tumour cells,?benign/?malig|8001/1
C0431085|T025|OP|BB0z.|RCDSY|Unspecified tumour cell NOS|8001/1
C0431085|T025|SY|252987004|SNOMEDCT_US|Tumor cell|8001/1
C0431085|T025|PT|252987004|SNOMEDCT_US|Tumor cells|8001/1
C0431085|T025|SY|39577004|SNOMEDCT_US|Tumor cells|8001/1
C0431085|T025|IS|39577004|SNOMEDCT_US|Tumor cells, NOS|8001/1
C0431085|T025|OAP|189544001|SNOMEDCT_US|Tumor cells, uncertain whether benign or malignant|8001/1
C0431085|T025|PT|39577004|SNOMEDCT_US|Tumor cells, uncertain whether benign or malignant|8001/1
C0431085|T025|SYGB|252987004|SNOMEDCT_US|Tumour cell|8001/1
C0431085|T025|PTGB|252987004|SNOMEDCT_US|Tumour cells|8001/1
C0431085|T025|SYGB|39577004|SNOMEDCT_US|Tumour cells|8001/1
C0431085|T025|IS|39577004|SNOMEDCT_US|Tumour cells, NOS|8001/1
C0431085|T025|PTGB|39577004|SNOMEDCT_US|Tumour cells, uncertain whether benign or malignant|8001/1
C0431085|T025|OAP|189544001|SNOMEDCT_US|Tumour cells, uncertain whether benign or malignant|8001/1
C0334227|T025|PT|0000029940|CHV|cancer cell|8001/3
C0334227|T025|SY|0000029940|CHV|cancer cells|8001/3
C0334227|T025|SY|0000029940|CHV|cancers cell|8001/3
C0334227|T025|SY|0000058033|CHV|cells malignant|8001/3
C0334227|T025|SY|0000058033|CHV|malignant cell|8001/3
C0334227|T025|PT|0000058033|CHV|malignant cells|8001/3
C0334227|T025|ET|2027-2183|CSP|cancer cell|8001/3
C0334227|T025|CN|MTHU015734|LNC|Malignant cells|8001/3
C0334227|T025|LPN|LP31549-6|LNC|Malignant cells|8001/3
C0334227|T025|SY|C12917|NCI|Cancer Cell|8001/3
C0334227|T025|PT|C12917|NCI|Malignant Cell|8001/3
C0334227|T025|SY|TCGA|NCI|Malignant Cell|8001/3
C0334227|T025|PT|BB07.|RCD|Malignant tumour cells|8001/3
C0334227|T025|PT|BB07.|RCDAE|Malignant tumor cells|8001/3
C0334227|T025|SY|88400008|SNOMEDCT_US|Malignant tumor cells|8001/3
C0334227|T025|SYGB|88400008|SNOMEDCT_US|Malignant tumour cells|8001/3
C0334227|T025|PT|88400008|SNOMEDCT_US|Tumor cells, malignant|8001/3
C0334227|T025|PTGB|88400008|SNOMEDCT_US|Tumour cells, malignant|8001/3
C0334228|T191|PT|0046790|CCPSS|SMALL CELL TUMOR MALIGNANT|8002/3
C0334228|T191|OP|C65154|NCI|Malignant Tumor, Small Cell Type|8002/3
C0334228|T191|PT|C65154|NCI|Malignant Tumor, Small Cell Type|8002/3
C0334228|T191|AB|BB08.|RCD|Malignant tumour - small cell|8002/3
C0334228|T191|PT|BB08.|RCD|Malignant tumour - small cell type|8002/3
C0334228|T191|AB|BB08.|RCDAE|Malignant tumor - small cell|8002/3
C0334228|T191|PT|BB08.|RCDAE|Malignant tumor - small cell type|8002/3
C0334228|T191|SY|82267002|SNOMEDCT_US|Malignant tumor - small cell type|8002/3
C0334228|T191|PT|82267002|SNOMEDCT_US|Malignant tumor, small cell type|8002/3
C0334228|T191|SYGB|82267002|SNOMEDCT_US|Malignant tumour - small cell type|8002/3
C0334228|T191|PTGB|82267002|SNOMEDCT_US|Malignant tumour, small cell type|8002/3
C0334229|T191|LLT|10025564|MDR|Malignant giant cell tumor|8003/3
C0334229|T191|LLT|10062857|MDR|Malignant giant cell tumour|8003/3
C0334229|T191|PT|271465|MEDCIN|giant cell type neoplasm|8003/3
C0334229|T191|SY|271465|MEDCIN|malignant giant cell neoplasm|8003/3
C0334229|T191|PT|C4090|NCI|Malignant Giant Cell Neoplasm|8003/3
C0334229|T191|SY|C4090|NCI|Malignant Giant Cell Tumor|8003/3
C0334229|T191|PT|C4090|NCI_CDISC|GIANT CELL TUMOR, MALIGNANT|8003/3
C0334229|T191|SY|C4090|NCI_CDISC|Malignant Giant Cell Tumor|8003/3
C0334229|T191|PT|C4090|NCI_CPTAC|Malignant Giant Cell Neoplasm|8003/3
C0334229|T191|AB|BB09.|RCD|Malignant tumour - giant cell|8003/3
C0334229|T191|PT|BB09.|RCD|Malignant tumour - giant cell type|8003/3
C0334229|T191|AB|BB09.|RCDAE|Malignant tumor - giant cell|8003/3
C0334229|T191|PT|BB09.|RCDAE|Malignant tumor - giant cell type|8003/3
C0334229|T191|SY|83950009|SNOMEDCT_US|Malignant tumor - giant cell type|8003/3
C0334229|T191|PT|83950009|SNOMEDCT_US|Malignant tumor, giant cell type|8003/3
C0334229|T191|SYGB|83950009|SNOMEDCT_US|Malignant tumour - giant cell type|8003/3
C0334229|T191|PTGB|83950009|SNOMEDCT_US|Malignant tumour, giant cell type|8003/3
C0334230|T191|SY|271441|MEDCIN|malignant spindle cell neoplasm|8004/3
C0334230|T191|PT|271441|MEDCIN|spindle cell type neoplasm|8004/3
C0334230|T191|PT|C27091|NCI|Malignant Spindle Cell Neoplasm|8004/3
C0334230|T191|SY|TCGA|NCI|Malignant Spindle Cell Neoplasm|8004/3
C0334230|T191|SY|C27091|NCI|Malignant Spindle Cell Tumor|8004/3
C0334230|T191|SY|C27091|NCI|Spindle Cell Cancer|8004/3
C0334230|T191|PT|CDR0000044506|NCI_NCI-GLOSS|spindle cell cancer|8004/3
C0334230|T191|AB|BB0A.|RCD|Malign tumour - fusiform cell|8004/3
C0334230|T191|AB|BB0A.|RCD|Malign tumour - spindle cell|8004/3
C0334230|T191|PT|BB0A.|RCD|Malignant tumour - fusiform cell type|8004/3
C0334230|T191|SY|BB0A.|RCD|Malignant tumour - spindle cell type|8004/3
C0334230|T191|AB|BB0A.|RCDAE|Malign tumor - fusiform cell|8004/3
C0334230|T191|AB|BB0A.|RCDAE|Malign tumor - spindle cell|8004/3
C0334230|T191|PT|BB0A.|RCDAE|Malignant tumor - fusiform cell type|8004/3
C0334230|T191|SY|BB0A.|RCDAE|Malignant tumor - spindle cell type|8004/3
C0334230|T191|SY|88897007|SNOMEDCT_US|Malignant tumor - fusiform cell type|8004/3
C0334230|T191|SY|88897007|SNOMEDCT_US|Malignant tumor - spindle cell type|8004/3
C0334230|T191|PT|88897007|SNOMEDCT_US|Malignant tumor, fusiform cell type|8004/3
C0334230|T191|SY|88897007|SNOMEDCT_US|Malignant tumor, spindle cell type|8004/3
C0334230|T191|SYGB|88897007|SNOMEDCT_US|Malignant tumour - fusiform cell type|8004/3
C0334230|T191|SYGB|88897007|SNOMEDCT_US|Malignant tumour - spindle cell type|8004/3
C0334230|T191|PTGB|88897007|SNOMEDCT_US|Malignant tumour, fusiform cell type|8004/3
C0334230|T191|SYGB|88897007|SNOMEDCT_US|Malignant tumour, spindle cell type|8004/3
C1265994|T191|SY|0000056674|CHV|cell clear tumors|8005/0
C1265994|T191|PT|0000056674|CHV|clear cell tumor|8005/0
C1265994|T191|OP|C66752|NCI|Clear Cell Neoplasm|8005/0
C1265994|T191|PT|C66752|NCI|Clear Cell Neoplasm|8005/0
C1265994|T191|OP|C66752|NCI|Clear Cell Tumor|8005/0
C1265994|T191|PT|128626003|SNOMEDCT_US|Clear cell tumor|8005/0
C1265994|T191|PTGB|128626003|SNOMEDCT_US|Clear cell tumour|8005/0
C1880101|T191|PT|271393|MEDCIN|clear cell type neoplasm|8005/3
C1880101|T191|SY|271393|MEDCIN|malignant clear cell neoplasm|8005/3
C1880101|T191|PT|C65156|NCI|Clear Cell Malignant Neoplasm|8005/3
C1880101|T191|OP|C65156|NCI|Clear Cell Malignant Neoplasm|8005/3
C1265995|T191|PT|128627007|SNOMEDCT_US|Malignant tumor, clear cell type|8005/3
C1265995|T191|PTGB|128627007|SNOMEDCT_US|Malignant tumour, clear cell type|8005/3
C0302894|T047|SY|0000028017|CHV|keratosis stucco|8010/0
C0302894|T047|PT|0000028017|CHV|stucco keratosis|8010/0
C0302894|T047|LLT|10081864|MDR|Stucco keratosis|8010/0
C0334232|T191|PN|NOCODE|MTH|Benign Epithelioma|8010/0
C1275160|T191|PN|NOCODE|MTH|Eruptive seborrheic keratosis|8010/0
C0334232|T191|PT|C4092|NCI|Benign Epithelial Neoplasm|8010/0
C0334232|T191|SY|C4092|NCI|Benign Epithelial Tumor|8010/0
C0334232|T191|SY|C4092|NCI|Benign Epithelioma|8010/0
C0334232|T191|SY|C4092|NCI|Benign Neoplasm of Epithelium|8010/0
C0334232|T191|SY|C4092|NCI|Benign Neoplasm of the Epithelium|8010/0
C0334232|T191|SY|C4092|NCI|Benign Tumor of Epithelium|8010/0
C0334232|T191|SY|C4092|NCI|Benign Tumor of the Epithelium|8010/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Epithelial Tumor|8010/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Epithelioma|8010/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Neoplasm of Epithelium|8010/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Neoplasm of the Epithelium|8010/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Tumor of Epithelium|8010/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Tumor of the Epithelium|8010/0
C0334232|T191|PT|C4092|NCI_CDISC|EPITHELIOMA, BENIGN|8010/0
C0334232|T191|PT|X77mx|RCD|Benign epithelial tumour|8010/0
C0334232|T191|PT|BB15.|RCD|Benign epithelioma|8010/0
C0334232|T191|PT|X77mx|RCDAE|Benign epithelial tumor|8010/0
C0334232|T191|OP|BB10.|RCDSA|Epithelial tumor, benign|8010/0
C0334232|T191|OP|BB10.|RCDSY|Epithelial tumour, benign|8010/0
C1302886|T191|PT|400207007|SNOMEDCT_US|Benign epithelial neoplasm - category|8010/0
C0334232|T191|SY|42535003|SNOMEDCT_US|Benign epithelial tumor|8010/0
C0334232|T191|SYGB|42535003|SNOMEDCT_US|Benign epithelial tumour|8010/0
C0334232|T191|SY|63823009|SNOMEDCT_US|Benign epithelioma|8010/0
C0334232|T191|PT|42535003|SNOMEDCT_US|Epithelial tumor, benign|8010/0
C0334232|T191|SY|42535003|SNOMEDCT_US|Epithelial tumor, benign, no ICD-O subtype|8010/0
C0334232|T191|SY|42535003|SNOMEDCT_US|Epithelial tumor, benign, no International Classification of Diseases for Oncology subtype|8010/0
C0334232|T191|PTGB|42535003|SNOMEDCT_US|Epithelial tumour, benign|8010/0
C0334232|T191|PT|63823009|SNOMEDCT_US|Epithelioma, benign|8010/0
C1275160|T191|PT|403868009|SNOMEDCT_US|Eruptive basal cell papillomata|8010/0
C1275160|T191|PT|786905007|SNOMEDCT_US|Eruptive seborrheic keratosis|8010/0
C1275160|T191|SY|403868009|SNOMEDCT_US|Eruptive seborrheic keratosis|8010/0
C1275160|T191|PTGB|786905007|SNOMEDCT_US|Eruptive seborrhoeic keratosis|8010/0
C1275160|T191|SYGB|403868009|SNOMEDCT_US|Eruptive seborrhoeic keratosis|8010/0
C1274598|T047|PT|786035003|SNOMEDCT_US|Multiple actinic keratoses|8010/0
C1274598|T047|PT|403202002|SNOMEDCT_US|Multiple actinic keratoses|8010/0
C5192272|T191|PT|786907004|SNOMEDCT_US|Multiple fibroepithelial polyps|8010/0
C1274598|T047|SY|403202002|SNOMEDCT_US|Multiple solar keratoses|8010/0
C0302894|T047|IS|25499005|SNOMEDCT_US|Stucco keratosis|8010/0
C0302894|T047|PT|403869001|SNOMEDCT_US|Stucco keratosis|8010/0
C0302894|T047|PT|103671002|SNOMEDCT_US|Stucco keratosis|8010/0
C0007099|T191|PT|1013022|CCPSS|CARCINOMA IN SITU|8010/2
C0007099|T191|PT|0000002417|CHV|carcinoma in situ|8010/2
C0007099|T191|SY|0000002417|CHV|carcinoma in-situ|8010/2
C0007099|T191|SY|0000002417|CHV|carcinoma situ|8010/2
C0007099|T191|SY|0000002417|CHV|in situ carcinoma|8010/2
C0007099|T191|SY|0000002417|CHV|in-situ carcinoma|8010/2
C0007099|T191|SY|0000002417|CHV|intraepithelial carcinoma|8010/2
C0007099|T191|PT|D09.9|ICD10|Carcinoma in situ, unspecified|8010/2
C0007099|T191|AB|D09.9|ICD10CM|Carcinoma in situ, unspecified|8010/2
C0007099|T191|PT|D09.9|ICD10CM|Carcinoma in situ, unspecified|8010/2
C0007099|T191|AB|234.9|ICD9CM|Ca in situ NOS|8010/2
C0007099|T191|HT|230-234.99|ICD9CM|CARCINOMA IN SITU|8010/2
C0007099|T191|PT|234.9|ICD9CM|Carcinoma in situ, site unspecified|8010/2
C0007099|T191|PT|A79004|ICPC2P|Carcinoma in situ|8010/2
C0007099|T191|PTN|A79004|ICPC2P|carcinoma in situ|8010/2
C0007099|T191|PT|10061450|MDR|Carcinoma in situ|8010/2
C0007099|T191|LLT|10061450|MDR|Carcinoma in situ|8010/2
C0007099|T191|LLT|10007353|MDR|Carcinoma in situ NOS|8010/2
C0007099|T191|LLT|10007402|MDR|Carcinoma in situ, site unspecified|8010/2
C0007099|T191|PT|99806|MEDCIN|carcinoma in situ|8010/2
C0007099|T191|MH|D002278|MSH|Carcinoma in Situ|8010/2
C0007099|T191|ET|D002278|MSH|Carcinoma, Intraepithelial|8010/2
C0007099|T191|ET|D002278|MSH|Carcinoma, Preinvasive|8010/2
C0007099|T191|PM|D002278|MSH|Intraepithelial Carcinoma|8010/2
C0007099|T191|PM|D002278|MSH|Preinvasive Carcinoma|8010/2
C0007099|T191|PN|NOCODE|MTH|Carcinoma in Situ|8010/2
C0007099|T191|ET|234.9|MTHICD9|Carcinoma in situ NOS|8010/2
C0007099|T191|PT|C2917|NCI|Carcinoma In Situ|8010/2
C0007099|T191|AB|C2917|NCI|CIS|8010/2
C0007099|T191|SY|C2917|NCI|Intraepithelial Carcinoma|8010/2
C0007099|T191|SY|C2917|NCI|Non-invasive Carcinoma|8010/2
C0007099|T191|PT|C2917|NCI_CDISC|CARCINOMA, IN SITU, MALIGNANT|8010/2
C0007099|T191|SY|C2917|NCI_CDISC|CIS|8010/2
C0007099|T191|SY|C2917|NCI_CDISC|Epithelial Tumor, In situ, Malignant|8010/2
C0007099|T191|SY|C2917|NCI_CDISC|Intraepithelial Carcinoma|8010/2
C0007099|T191|SY|C2917|NCI_CDISC|Non-invasive Carcinoma|8010/2
C0007099|T191|PT|C2917|NCI_CPTAC|Carcinoma In Situ|8010/2
C0007099|T191|PT|CDR0000046488|NCI_NCI-GLOSS|carcinoma in situ|8010/2
C0007099|T191|PT|CDR0000638178|NCI_NCI-GLOSS|stage 0 disease|8010/2
C0007099|T191|SY|Xa986|RCD|Carcinoma in situ|8010/2
C0007099|T191|SY|XE2xD|RCD|Carcinoma in situ|8010/2
C0007099|T191|PT|Xa986|RCD|Carcinoma in situ morphology|8010/2
C0007099|T191|OP|B8z..|RCD|Carcinoma in situ NOS|8010/2
C0007099|T191|PT|XE2xD|RCD|Carcinoma in situ tumour|8010/2
C0007099|T191|SY|XE2xD|RCD|CIS - Carcinoma in situ|8010/2
C0007099|T191|SY|Xa986|RCD|Intraepithelial carcinoma|8010/2
C0007099|T191|PT|XE2xD|RCDAE|Carcinoma in situ tumor|8010/2
C0007099|T191|OP|BB11.|RCDSY|Carcinoma in situ NOS|8010/2
C0007099|T191|SY|109355002|SNOMEDCT_US|Cancer in situ|8010/2
C0007099|T191|OAS|189208007|SNOMEDCT_US|Carcinoma in situ|8010/2
C0007099|T191|OAS|271528002|SNOMEDCT_US|Carcinoma in situ|8010/2
C0007099|T191|PT|109355002|SNOMEDCT_US|Carcinoma in situ|8010/2
C0007099|T191|PT|68956006|SNOMEDCT_US|Carcinoma in situ|8010/2
C0007099|T191|PT|399919001|SNOMEDCT_US|Carcinoma in situ - category|8010/2
C0007099|T191|SY|68956006|SNOMEDCT_US|Carcinoma in situ morphology|8010/2
C0007099|T191|OAP|154640008|SNOMEDCT_US|Carcinoma in situ NOS|8010/2
C0007099|T191|OAP|189359006|SNOMEDCT_US|Carcinoma in situ NOS|8010/2
C0007099|T191|OF|154640008|SNOMEDCT_US|Carcinoma in situ NOS|8010/2
C0007099|T191|OAP|271528002|SNOMEDCT_US|Carcinoma in situ tumor|8010/2
C0007099|T191|OAP|154635000|SNOMEDCT_US|Carcinoma in situ tumor|8010/2
C0007099|T191|OF|271528002|SNOMEDCT_US|Carcinoma in situ tumour|8010/2
C0007099|T191|OAP|271528002|SNOMEDCT_US|Carcinoma in situ tumour|8010/2
C0007099|T191|OAP|154635000|SNOMEDCT_US|Carcinoma in situ tumour|8010/2
C0007099|T191|OF|154635000|SNOMEDCT_US|Carcinoma in situ tumour|8010/2
C0007099|T191|SY|68956006|SNOMEDCT_US|Carcinoma in situ, no ICD-O subtype|8010/2
C0007099|T191|SY|68956006|SNOMEDCT_US|Carcinoma in situ, no International Classification of Diseases for Oncology subtype|8010/2
C0007099|T191|IS|68956006|SNOMEDCT_US|Carcinoma in situ, NOS|8010/2
C0007099|T191|OAS|271528002|SNOMEDCT_US|CIS - Carcinoma in situ|8010/2
C0007099|T191|SY|68956006|SNOMEDCT_US|Intraepithelial carcinoma|8010/2
C0007099|T191|IS|68956006|SNOMEDCT_US|Intraepithelial carcinoma, NOS|8010/2
C0007099|T191|SY|399919001|SNOMEDCT_US|Non-invasive carcinoma|8010/2
C0007097|T191|DE|0000004525|AOD|carcinoma|8010/3
C0007097|T191|PT|1018250|CCPSS|CARCINOMA|8010/3
C0741899|T191|PT|1017412|CCPSS|CARCINOMA POORLY DIFFERENTIATED|8010/3
C0349561|T191|SY|0000021165|CHV|bartholin's cancer gland|8010/3
C0349561|T191|PT|0000021165|CHV|bartholin's gland cancer|8010/3
C0007097|T191|PT|0000002416|CHV|carcinoma|8010/3
C0741899|T191|PT|0000047325|CHV|carcinoma poorly differentiated|8010/3
C0007097|T191|SY|0000002416|CHV|carcinomas|8010/3
C0007097|T191|SY|0000002416|CHV|epithelioma|8010/3
C0007097|T191|SY|0000002416|CHV|epitheliomas|8010/3
C0741899|T191|SY|0000047325|CHV|poorly differentiated carcinoma|8010/3
C0007097|T191|PT|134|COSTAR|CARCINOMA|8010/3
C0007097|T191|PT|2000-1867|CSP|carcinoma|8010/3
C0007097|T191|PT|CARCINOMA|CST|CARCINOMA|8010/3
C0007097|T191|SY|NOCODE|DXP|CARCINOMA|8010/3
C0349561|T191|PT|HP:0030419|HPO|Bartholin gland carcinoma|8010/3
C0007097|T191|PT|HP:0030731|HPO|Carcinoma|8010/3
C0007097|T191|PT|MTHU014804|ICPC2ICD10ENG|carcinoma; unspecified site, unspecified site|8010/3
C0007097|T191|PT|MTHU053524|ICPC2ICD10ENG|unspecified site; carcinoma, unspecified site|8010/3
C0007097|T191|LA|LA15448-6|LNC|Carcinoma|8010/3
C0007097|T191|LLT|10007284|MDR|Carcinoma|8010/3
C0007097|T191|LLT|10007423|MDR|Carcinoma NOS|8010/3
C0007097|T191|PT|271392|MEDCIN|carcinoma|8010/3
C0349561|T191|PT|352123|MEDCIN|Carcinoma of Bartholin's gland|8010/3
C0349561|T191|SY|352123|MEDCIN|vulvar neoplasm malignant Bartholin's gland carcinoma|8010/3
C0007097|T191|SY|25|MEDLINEPLUS|Carcinoma|8010/3
C0007097|T191|ET|25|MEDLINEPLUS|Carcinoma|8010/3
C0007097|T191|MH|D002277|MSH|Carcinoma|8010/3
C0007097|T191|PM|D002277|MSH|Carcinomas|8010/3
C0007097|T191|DEV|D002277|MSH|EPITHELIAL NEOPL MALIGNANT|8010/3
C0007097|T191|PM|D002277|MSH|Epithelial Neoplasm, Malignant|8010/3
C0007097|T191|ET|D002277|MSH|Epithelial Neoplasms, Malignant|8010/3
C0007097|T191|PM|D002277|MSH|Epithelial Tumor, Malignant|8010/3
C0007097|T191|ET|D002277|MSH|Epithelial Tumors, Malignant|8010/3
C0007097|T191|ET|D002277|MSH|Epithelioma|8010/3
C0007097|T191|PM|D002277|MSH|Epitheliomas|8010/3
C0007097|T191|DEV|D002277|MSH|MALIGNANT EPITHELIAL NEOPL|8010/3
C0007097|T191|PM|D002277|MSH|Malignant Epithelial Neoplasm|8010/3
C0007097|T191|ET|D002277|MSH|Malignant Epithelial Neoplasms|8010/3
C0007097|T191|PM|D002277|MSH|Malignant Epithelial Tumor|8010/3
C0007097|T191|PM|D002277|MSH|Malignant Epithelial Tumors|8010/3
C0007097|T191|DEV|D002277|MSH|NEOPL MALIGNANT EPITHELIAL|8010/3
C0007097|T191|PM|D002277|MSH|Neoplasm, Malignant Epithelial|8010/3
C0007097|T191|ET|D002277|MSH|Neoplasms, Malignant Epithelial|8010/3
C0007097|T191|PM|D002277|MSH|Tumor, Malignant Epithelial|8010/3
C0007097|T191|PN|NOCODE|MTH|Carcinoma|8010/3
C0349561|T191|PT|C9055|NCI|Bartholin Gland Carcinoma|8010/3
C0349561|T191|SY|C9055|NCI|Bartholin's Gland Cancer|8010/3
C0349561|T191|SY|C9055|NCI|Bartholin's Gland Carcinoma|8010/3
C0007097|T191|PT|C2916|NCI|Carcinoma|8010/3
C0007097|T191|SY|TCGA|NCI|Carcinoma|8010/3
C0349561|T191|SY|C9055|NCI|Carcinoma of Bartholin's Gland|8010/3
C0349561|T191|SY|C9055|NCI|Carcinoma of the Bartholin's Gland|8010/3
C0007097|T191|SY|C2916|NCI|Epithelial Carcinoma|8010/3
C0007097|T191|SY|C2916|NCI|Malignant Epithelial Neoplasm|8010/3
C0007097|T191|SY|C2916|NCI|Malignant Epithelial Tumor|8010/3
C0007097|T191|SY|C2916|NCI|Malignant Epithelioma|8010/3
C0007097|T191|PT|C2916|NCI_CDISC|CARCINOMA, MALIGNANT|8010/3
C0007097|T191|SY|C2916|NCI_CDISC|Epithelial Carcinoma|8010/3
C0007097|T191|SY|C2916|NCI_CDISC|Epithelioma Malignant|8010/3
C0007097|T191|SY|C2916|NCI_CDISC|Malignant Epithelial Neoplasm|8010/3
C0007097|T191|SY|C2916|NCI_CDISC|Malignant Epithelial Tumor|8010/3
C0007097|T191|SY|C2916|NCI_CDISC|Malignant Epithelioma|8010/3
C0007097|T191|PT|C2916|NCI_CPTAC|Carcinoma|8010/3
C0007097|T191|PT|10007423|NCI_CTEP-SDC|Carcinoma, NOS|8010/3
C0349561|T191|DN|C9055|NCI_CTRP|Bartholin Gland Cancer|8010/3
C0007097|T191|PT|C2916|NCI_CTRP|Carcinoma|8010/3
C0007097|T191|DN|C2916|NCI_CTRP|Other Carcinoma|8010/3
C0007097|T191|PT|CDR0000045963|NCI_NCI-GLOSS|carcinoma|8010/3
C0007097|T191|PT|CDR0000046422|NCI_NCI-GLOSS|epithelial carcinoma|8010/3
C0007097|T191|ET|07590|PSY|Carcinomas|8010/3
C0007097|T191|PT|Xa987|RCD|Carcinoma|8010/3
C0349561|T191|PT|Xa0Eq|RCD|Carcinoma of Bartholin's gland|8010/3
C0007097|T191|SY|Xa987|RCD|Malignant epithelial tumour|8010/3
C0007097|T191|SY|Xa987|RCDAE|Malignant epithelial tumor|8010/3
C0007097|T191|OP|BB12.|RCDSY|Carcinoma NOS|8010/3
C0349561|T191|SY|399533005|SNOMEDCT_US|Bartholin gland carcinoma|8010/3
C0349561|T191|PT|399533005|SNOMEDCT_US|Bartholin's gland carcinoma|8010/3
C0007097|T191|OAS|269513004|SNOMEDCT_US|Carcinoma|8010/3
C0007097|T191|OAS|154433003|SNOMEDCT_US|Carcinoma|8010/3
C0007097|T191|SY|722688002|SNOMEDCT_US|Carcinoma|8010/3
C0007097|T191|PT|68453008|SNOMEDCT_US|Carcinoma|8010/3
C0349561|T191|SY|276876007|SNOMEDCT_US|Carcinoma of Bartholin gland|8010/3
C0349561|T191|PT|276876007|SNOMEDCT_US|Carcinoma of Bartholin's gland|8010/3
C1273670|T191|PT|384950003|SNOMEDCT_US|Carcinoma with pleomorphic, sarcomatoid or sarcomatous elements|8010/3
C0007097|T191|SY|68453008|SNOMEDCT_US|Carcinoma, no subtype|8010/3
C0007097|T191|IS|68453008|SNOMEDCT_US|Carcinoma, NOS|8010/3
C0007097|T191|SY|68453008|SNOMEDCT_US|Epithelial tumor, malignant|8010/3
C0007097|T191|SYGB|68453008|SNOMEDCT_US|Epithelial tumour, malignant|8010/3
C0007097|T191|PT|722688002|SNOMEDCT_US|Malignant epithelial neoplasm|8010/3
C0007097|T191|SY|68453008|SNOMEDCT_US|Malignant epithelial tumor|8010/3
C0007097|T191|SYGB|68453008|SNOMEDCT_US|Malignant epithelial tumour|8010/3
C0741899|T191|PT|703078002|SNOMEDCT_US|Poorly differentiated carcinoma|8010/3
C0007097|T191|PT|0746|WHO|CARCINOMA|8010/3
C1384494|T191|SY|0000015723|CHV|carcinoma metastatic|8010/6
C1384494|T191|PT|0000015723|CHV|metastatic carcinoma|8010/6
C1384494|T191|PT|U000442|COSTAR|METASTATIC CARCINOMA|8010/6
C1384494|T191|LLT|10027477|MDR|Metastatic carcinoma|8010/6
C1384494|T191|PN|NOCODE|MTH|Metastatic Carcinoma|8010/6
C1384494|T191|PT|C3482|NCI|Metastatic Carcinoma|8010/6
C1384494|T191|DN|C3482|NCI_CTRP|Metastatic Carcinoma|8010/6
C1384494|T191|PT|XM1GJ|RCD|Metastatic carcinoma|8010/6
C1384494|T191|OP|BB13.|RCDSY|Carcinoma, metastatic, NOS|8010/6
C1384494|T191|PT|79282002|SNOMEDCT_US|Carcinoma, metastatic|8010/6
C1384494|T191|IS|79282002|SNOMEDCT_US|Carcinoma, metastatic, NOS|8010/6
C1384494|T191|OAS|269624009|SNOMEDCT_US|Metastatic carcinoma|8010/6
C1384494|T191|OAS|154576004|SNOMEDCT_US|Metastatic carcinoma|8010/6
C0205699|T191|PT|0000020685|CHV|carcinomatosis|8010/9
C0205699|T191|PT|U000013|COSTAR|CARCINOMATOSIS|8010/9
C0205699|T191|ET|C80.0|ICD10CM|Carcinomatosis NOS|8010/9
C0205699|T191|LA|LA9144-2|LNC|Carcinomatosis|8010/9
C0205699|T191|LLT|10007506|MDR|Carcinomatosis|8010/9
C0577731|T191|LLT|10013430|MDR|Disseminated adenocarcinoma|8010/9
C0205699|T191|PM|D002277|MSH|Carcinomatoses|8010/9
C0205699|T191|PEP|D002277|MSH|Carcinomatosis|8010/9
C0205699|T191|PN|NOCODE|MTH|Carcinomatosis|8010/9
C0205699|T191|PT|C3693|NCI|Carcinomatosis|8010/9
C0577731|T191|PT|C27185|NCI|Disseminated Adenocarcinoma|8010/9
C0205699|T191|PT|CDR0000257223|NCI_NCI-GLOSS|carcinomatosis|8010/9
C0205699|T191|PT|CDR0000285963|NCI_NCI-GLOSS|carcinosis|8010/9
C0205699|T191|PT|XaBAn|RCD|Carcinomatosis|8010/9
C0577731|T191|PT|Xa7o3|RCD|Disseminated adenocarcinoma|8010/9
C0205699|T191|SY|XaBAn|RCD|Disseminated carcinomatosis|8010/9
C0205699|T191|PT|BB14.|RCDSY|Carcinomatosis|8010/9
C0205699|T191|OAS|188476000|SNOMEDCT_US|Carcinomatosis|8010/9
C0205699|T191|PT|307593001|SNOMEDCT_US|Carcinomatosis|8010/9
C0205699|T191|OAS|269624009|SNOMEDCT_US|Carcinomatosis|8010/9
C0205699|T191|PT|7010000|SNOMEDCT_US|Carcinomatosis|8010/9
C0205699|T191|OAS|154576004|SNOMEDCT_US|Carcinomatosis|8010/9
C0577731|T191|PT|301036008|SNOMEDCT_US|Disseminated adenocarcinoma|8010/9
C0205699|T191|SY|307593001|SNOMEDCT_US|Disseminated carcinomatosis|8010/9
C0205699|T191|IT|1259|WHO|CARCINOMATOSIS|8010/9
C0346027|T191|SY|0000031042|CHV|carcinomas syringomatous|8011/0
C0346027|T191|PT|0000031042|CHV|microcystic adnexal carcinoma|8011/0
C0346027|T191|LLT|10073091|MDR|Microcystic adnexal carcinoma|8011/0
C0346027|T191|PT|231630|MEDCIN|sclerosing carcinoma of sweat duct|8011/0
C0346027|T191|SY|231630|MEDCIN|sclerosing sweat duct carcinoma|8011/0
C0346027|T191|NM|C000632664|MSH|Microcystic adnexal carcinoma|8011/0
C0334232|T191|PN|NOCODE|MTH|Benign Epithelioma|8011/0
C0334232|T191|PT|C4092|NCI|Benign Epithelial Neoplasm|8011/0
C0334232|T191|SY|C4092|NCI|Benign Epithelial Tumor|8011/0
C0334232|T191|SY|C4092|NCI|Benign Epithelioma|8011/0
C0334232|T191|SY|C4092|NCI|Benign Neoplasm of Epithelium|8011/0
C0334232|T191|SY|C4092|NCI|Benign Neoplasm of the Epithelium|8011/0
C0334232|T191|SY|C4092|NCI|Benign Tumor of Epithelium|8011/0
C0334232|T191|SY|C4092|NCI|Benign Tumor of the Epithelium|8011/0
C0346027|T191|SY|C7581|NCI|Eccrine Epithelioma|8011/0
C0346027|T191|PT|C7581|NCI|Microcystic Adnexal Carcinoma|8011/0
C0346027|T191|SY|C7581|NCI|Syringomatous Carcinoma|8011/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Epithelial Tumor|8011/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Epithelioma|8011/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Neoplasm of Epithelium|8011/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Neoplasm of the Epithelium|8011/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Tumor of Epithelium|8011/0
C0334232|T191|SY|C4092|NCI_CDISC|Benign Tumor of the Epithelium|8011/0
C0334232|T191|PT|C4092|NCI_CDISC|EPITHELIOMA, BENIGN|8011/0
C0334232|T191|PT|X77mx|RCD|Benign epithelial tumour|8011/0
C0334232|T191|PT|BB15.|RCD|Benign epithelioma|8011/0
C0346027|T191|PT|X78Sx|RCD|Eccrine epithelioma|8011/0
C0346027|T191|SY|X78Si|RCD|Malignant syringoma|8011/0
C0346027|T191|PT|X78Si|RCD|Microcystic adnexal carcinoma|8011/0
C0346027|T191|AB|X78Si|RCD|Sclerosing sweat duct carcinom|8011/0
C0346027|T191|SY|X78Si|RCD|Sclerosing sweat duct carcinoma|8011/0
C0346027|T191|SY|X78Si|RCD|Syringoid eccrine carcinoma|8011/0
C0346027|T191|AB|X78Si|RCD|Syringomat sweat duct carcinom|8011/0
C0346027|T191|SY|X78Si|RCD|Syringomatous sweat duct carcinoma|8011/0
C0334232|T191|PT|X77mx|RCDAE|Benign epithelial tumor|8011/0
C0334232|T191|OP|BB10.|RCDSA|Epithelial tumor, benign|8011/0
C0334232|T191|OP|BB10.|RCDSY|Epithelial tumour, benign|8011/0
C0334232|T191|SY|42535003|SNOMEDCT_US|Benign epithelial tumor|8011/0
C0334232|T191|SYGB|42535003|SNOMEDCT_US|Benign epithelial tumour|8011/0
C0334232|T191|SY|63823009|SNOMEDCT_US|Benign epithelioma|8011/0
C0346027|T191|PT|400135003|SNOMEDCT_US|Eccrine epithelioma|8011/0
C0346027|T191|PT|254722001|SNOMEDCT_US|Eccrine epithelioma|8011/0
C0346027|T191|SY|254722001|SNOMEDCT_US|Eccrine epithelioma of skin|8011/0
C0334232|T191|PT|42535003|SNOMEDCT_US|Epithelial tumor, benign|8011/0
C0334232|T191|SY|42535003|SNOMEDCT_US|Epithelial tumor, benign, no ICD-O subtype|8011/0
C0334232|T191|SY|42535003|SNOMEDCT_US|Epithelial tumor, benign, no International Classification of Diseases for Oncology subtype|8011/0
C0334232|T191|PTGB|42535003|SNOMEDCT_US|Epithelial tumour, benign|8011/0
C0334232|T191|PT|63823009|SNOMEDCT_US|Epithelioma, benign|8011/0
C0346027|T191|SY|254712007|SNOMEDCT_US|Malignant syringoma|8011/0
C0346027|T191|PT|254712007|SNOMEDCT_US|Microcystic adnexal carcinoma|8011/0
C0346027|T191|SY|128896007|SNOMEDCT_US|Microcystic adnexal carcinoma|8011/0
C0346027|T191|SY|254712007|SNOMEDCT_US|Microcystic adnexal carcinoma of skin|8011/0
C0346027|T191|SY|254712007|SNOMEDCT_US|Sclerosing sweat duct carcinoma|8011/0
C0346027|T191|PT|128896007|SNOMEDCT_US|Sclerosing sweat duct carcinoma|8011/0
C0346027|T191|SY|254712007|SNOMEDCT_US|Syringoid eccrine carcinoma|8011/0
C0346027|T191|SY|128896007|SNOMEDCT_US|Syringomatous carcinoma|8011/0
C0346027|T191|SY|254712007|SNOMEDCT_US|Syringomatous sweat duct carcinoma|8011/0
C0007097|T191|DE|0000004525|AOD|carcinoma|8011/3
C0007097|T191|PT|1018250|CCPSS|CARCINOMA|8011/3
C0007097|T191|PT|0000002416|CHV|carcinoma|8011/3
C0007097|T191|SY|0000002416|CHV|carcinomas|8011/3
C0007097|T191|SY|0000002416|CHV|epithelioma|8011/3
C0553707|T191|PT|0000039116|CHV|epithelioma|8011/3
C0007097|T191|SY|0000002416|CHV|epitheliomas|8011/3
C0007097|T191|PT|134|COSTAR|CARCINOMA|8011/3
C0007097|T191|PT|2000-1867|CSP|carcinoma|8011/3
C0007097|T191|PT|CARCINOMA|CST|CARCINOMA|8011/3
C0007097|T191|SY|NOCODE|DXP|CARCINOMA|8011/3
C0007097|T191|PT|HP:0030731|HPO|Carcinoma|8011/3
C0007097|T191|PT|MTHU014804|ICPC2ICD10ENG|carcinoma; unspecified site, unspecified site|8011/3
C0007097|T191|PT|MTHU053524|ICPC2ICD10ENG|unspecified site; carcinoma, unspecified site|8011/3
C0007097|T191|LA|LA15448-6|LNC|Carcinoma|8011/3
C0007097|T191|LLT|10007284|MDR|Carcinoma|8011/3
C0007097|T191|LLT|10007423|MDR|Carcinoma NOS|8011/3
C0007097|T191|PT|271392|MEDCIN|carcinoma|8011/3
C0553707|T191|SY|31726|MEDCIN|epithelioma|8011/3
C0553707|T191|PT|31726|MEDCIN|malignant epithelioma|8011/3
C0007097|T191|SY|25|MEDLINEPLUS|Carcinoma|8011/3
C0007097|T191|ET|25|MEDLINEPLUS|Carcinoma|8011/3
C0007097|T191|MH|D002277|MSH|Carcinoma|8011/3
C0007097|T191|PM|D002277|MSH|Carcinomas|8011/3
C0007097|T191|DEV|D002277|MSH|EPITHELIAL NEOPL MALIGNANT|8011/3
C0007097|T191|PM|D002277|MSH|Epithelial Neoplasm, Malignant|8011/3
C0007097|T191|ET|D002277|MSH|Epithelial Neoplasms, Malignant|8011/3
C0007097|T191|PM|D002277|MSH|Epithelial Tumor, Malignant|8011/3
C0007097|T191|ET|D002277|MSH|Epithelial Tumors, Malignant|8011/3
C0007097|T191|ET|D002277|MSH|Epithelioma|8011/3
C0007097|T191|PM|D002277|MSH|Epitheliomas|8011/3
C0007097|T191|DEV|D002277|MSH|MALIGNANT EPITHELIAL NEOPL|8011/3
C0007097|T191|PM|D002277|MSH|Malignant Epithelial Neoplasm|8011/3
C0007097|T191|ET|D002277|MSH|Malignant Epithelial Neoplasms|8011/3
C0007097|T191|PM|D002277|MSH|Malignant Epithelial Tumor|8011/3
C0007097|T191|PM|D002277|MSH|Malignant Epithelial Tumors|8011/3
C0007097|T191|DEV|D002277|MSH|NEOPL MALIGNANT EPITHELIAL|8011/3
C0007097|T191|PM|D002277|MSH|Neoplasm, Malignant Epithelial|8011/3
C0007097|T191|ET|D002277|MSH|Neoplasms, Malignant Epithelial|8011/3
C0007097|T191|PM|D002277|MSH|Tumor, Malignant Epithelial|8011/3
C0007097|T191|PN|NOCODE|MTH|Carcinoma|8011/3
C0553707|T191|PN|NOCODE|MTH|Malignant epithelioma|8011/3
C0007097|T191|PT|C2916|NCI|Carcinoma|8011/3
C0007097|T191|SY|TCGA|NCI|Carcinoma|8011/3
C0007097|T191|SY|C2916|NCI|Epithelial Carcinoma|8011/3
C0007097|T191|SY|C2916|NCI|Malignant Epithelial Neoplasm|8011/3
C0007097|T191|SY|C2916|NCI|Malignant Epithelial Tumor|8011/3
C0007097|T191|SY|C2916|NCI|Malignant Epithelioma|8011/3
C0007097|T191|PT|C2916|NCI_CDISC|CARCINOMA, MALIGNANT|8011/3
C0007097|T191|SY|C2916|NCI_CDISC|Epithelial Carcinoma|8011/3
C0007097|T191|SY|C2916|NCI_CDISC|Epithelioma Malignant|8011/3
C0007097|T191|SY|C2916|NCI_CDISC|Malignant Epithelial Neoplasm|8011/3
C0007097|T191|SY|C2916|NCI_CDISC|Malignant Epithelial Tumor|8011/3
C0007097|T191|SY|C2916|NCI_CDISC|Malignant Epithelioma|8011/3
C0007097|T191|PT|C2916|NCI_CPTAC|Carcinoma|8011/3
C0007097|T191|PT|10007423|NCI_CTEP-SDC|Carcinoma, NOS|8011/3
C0007097|T191|PT|C2916|NCI_CTRP|Carcinoma|8011/3
C0007097|T191|DN|C2916|NCI_CTRP|Other Carcinoma|8011/3
C0007097|T191|PT|CDR0000045963|NCI_NCI-GLOSS|carcinoma|8011/3
C0007097|T191|PT|CDR0000046422|NCI_NCI-GLOSS|epithelial carcinoma|8011/3
C0007097|T191|ET|07590|PSY|Carcinomas|8011/3
C0007097|T191|PT|Xa987|RCD|Carcinoma|8011/3
C0553707|T191|SY|BB16.|RCD|Epithelioma|8011/3
C0007097|T191|SY|Xa987|RCD|Malignant epithelial tumour|8011/3
C0553707|T191|PT|BB16.|RCD|Malignant epithelioma|8011/3
C0007097|T191|SY|Xa987|RCDAE|Malignant epithelial tumor|8011/3
C0007097|T191|OP|BB12.|RCDSY|Carcinoma NOS|8011/3
C0007097|T191|OAS|269513004|SNOMEDCT_US|Carcinoma|8011/3
C0007097|T191|OAS|154433003|SNOMEDCT_US|Carcinoma|8011/3
C0007097|T191|SY|722688002|SNOMEDCT_US|Carcinoma|8011/3
C0007097|T191|PT|68453008|SNOMEDCT_US|Carcinoma|8011/3
C0007097|T191|SY|68453008|SNOMEDCT_US|Carcinoma, no subtype|8011/3
C0007097|T191|IS|68453008|SNOMEDCT_US|Carcinoma, NOS|8011/3
C0007097|T191|SY|68453008|SNOMEDCT_US|Epithelial tumor, malignant|8011/3
C0007097|T191|SYGB|68453008|SNOMEDCT_US|Epithelial tumour, malignant|8011/3
C0553707|T191|SY|71298006|SNOMEDCT_US|Epithelioma|8011/3
C0553707|T191|PT|71298006|SNOMEDCT_US|Epithelioma, malignant|8011/3
C0553707|T191|IS|71298006|SNOMEDCT_US|Epithelioma, NOS|8011/3
C0007097|T191|PT|722688002|SNOMEDCT_US|Malignant epithelial neoplasm|8011/3
C0007097|T191|SY|68453008|SNOMEDCT_US|Malignant epithelial tumor|8011/3
C0007097|T191|SYGB|68453008|SNOMEDCT_US|Malignant epithelial tumour|8011/3
C0553707|T191|SY|71298006|SNOMEDCT_US|Malignant epithelioma|8011/3
C0007097|T191|PT|0746|WHO|CARCINOMA|8011/3
C0553707|T191|IT|1798|WHO|EPITHELIOMA|8011/3
C0206704|T191|PT|0010263|CCPSS|LARGE CELL CARCINOMA|8012/3
C0206704|T191|PT|0000021034|CHV|large cell carcinoma|8012/3
C0206704|T191|PT|U000035|COSTAR|LARGE CELL CARCINOMA|8012/3
C0206704|T191|PT|271394|MEDCIN|large cell carcinoma|8012/3
C0206704|T191|MH|D018287|MSH|Carcinoma, Large Cell|8012/3
C0206704|T191|PM|D018287|MSH|Carcinomas, Large Cell|8012/3
C0206704|T191|PM|D018287|MSH|Cell Carcinoma, Large|8012/3
C0206704|T191|PM|D018287|MSH|Cell Carcinomas, Large|8012/3
C0206704|T191|PM|D018287|MSH|Large Cell Carcinoma|8012/3
C0206704|T191|PM|D018287|MSH|Large Cell Carcinomas|8012/3
C0206704|T191|SY|C3780|NCI|Carcinoma, Large Cell|8012/3
C0206704|T191|PT|C3780|NCI|Large Cell Carcinoma|8012/3
C0206704|T191|SY|TCGA|NCI|Large Cell Carcinoma|8012/3
C0206704|T191|PT|C3780|NCI_CPTAC|Large Cell Carcinoma|8012/3
C0206704|T191|PT|CDR0000046316|NCI_NCI-GLOSS|large cell carcinoma|8012/3
C0206704|T191|PT|Xa988|RCD|Large cell carcinoma|8012/3
C0206704|T191|OP|BB17.|RCDSY|Large cell carcinoma NOS|8012/3
C0206704|T191|PT|22687000|SNOMEDCT_US|Large cell carcinoma|8012/3
C0206704|T191|IS|22687000|SNOMEDCT_US|Large cell carcinoma, NOS|8012/3
C1265996|T191|LA|LA26100-0|LNC|Large cell neuroendocrine carcinoma|8013/3
C1265996|T191|PT|271395|MEDCIN|large cell neuroendocrine carcinoma|8013/3
C1265996|T191|SY|C6875|NCI|Large Cell NEC|8013/3
C1265996|T191|PT|C6875|NCI|Large Cell Neuroendocrine Carcinoma|8013/3
C1265996|T191|SY|TCGA|NCI|Large Cell Neuroendocrine Carcinoma|8013/3
C1265996|T191|SY|C6875|NCI|Large-cell neuroendocrine carcinoma|8013/3
C1265996|T191|AB|C6875|NCI|LCNEC|8013/3
C1265996|T191|SY|CDR0000774873|PDQ|large cell NEC|8013/3
C1265996|T191|PT|CDR0000774873|PDQ|large cell neuroendocrine carcinoma|8013/3
C1265996|T191|SY|CDR0000774873|PDQ|large-cell neuroendocrine carcinoma|8013/3
C3163943|T191|PT|448546006|SNOMEDCT_US|Combined large cell neuroendocrine carcinoma|8013/3
C1265996|T191|IS|128628002|SNOMEDCT_US|Large cell neuroendocrine carcinoma|8013/3
C1265996|T191|PT|128628002|SNOMEDCT_US|Large cell neuroendocrine carcinoma|8013/3
C1265997|T191|PT|219566|MEDCIN|large cell carcinoma of lung with rhabdoid phenotype|8014/3
C1265997|T191|PT|271396|MEDCIN|large cell carcinoma with rhabdoid phenotype|8014/3
C1265997|T191|SY|271396|MEDCIN|malignant neoplasm carcinoma large cell with rhabdoid phenotype|8014/3
C1265997|T191|SY|C6876|NCI|Large Cell Carcinoma with Rhabdoid Phenotype|8014/3
C1265997|T191|SY|C6876|NCI|Large Cell Lung Carcinoma with Rhabdoid Phenotype|8014/3
C1265997|T191|PT|C6876|NCI|Lung Large Cell Carcinoma with Rhabdoid Phenotype|8014/3
C1265997|T191|PT|128629005|SNOMEDCT_US|Large cell carcinoma with rhabdoid phenotype|8014/3
C1265998|T191|PT|271397|MEDCIN|glassy cell carcinoma|8015/3
C1265998|T191|PT|C65159|NCI|Glassy Cell Carcinoma|8015/3
C1265998|T191|OP|C65159|NCI|Glassy Cell Carcinoma|8015/3
C1265998|T191|PT|128630000|SNOMEDCT_US|Glassy cell carcinoma|8015/3
C0205698|T191|SY|0000020684|CHV|carcinoma undifferentiated|8020/3
C0205698|T191|PT|0000020684|CHV|undifferentiated carcinoma|8020/3
C0205698|T191|LA|LA15447-8|LNC|Undifferentiated carcinoma|8020/3
C0205698|T191|PT|271398|MEDCIN|undifferentiated carcinoma|8020/3
C0205698|T191|PEP|D002277|MSH|Carcinoma, Undifferentiated|8020/3
C0205698|T191|PM|D002277|MSH|Undifferentiated Carcinoma|8020/3
C0205698|T191|PM|D002277|MSH|Undifferentiated Carcinomas|8020/3
C0205698|T191|PN|NOCODE|MTH|Undifferentiated carcinoma|8020/3
C0205698|T191|SY|C3692|NCI|Anaplastic Carcinoma|8020/3
C0205698|T191|SY|C3692|NCI|Carcinoma, Undifferentiated|8020/3
C0205698|T191|PT|C3692|NCI|Undifferentiated Carcinoma|8020/3
C0205698|T191|SY|TCGA|NCI|Undifferentiated Carcinoma|8020/3
C0205698|T191|SY|C3692|NCI_CDISC|Anaplastic Carcinoma|8020/3
C0205698|T191|SY|C3692|NCI_CDISC|Carcinoma, Undifferentiated|8020/3
C0205698|T191|PT|C3692|NCI_CDISC|CARCINOMA, UNDIFFERENTIATED, MALIGNANT|8020/3
C0205698|T191|PT|C3692|NCI_CPTAC|Undifferentiated Carcinoma|8020/3
C0205698|T191|PT|XM1F6|RCD|Undifferentiated carcinoma|8020/3
C0205698|T191|OA|BB18.|RCDSY|Carcinoma, undiff. type NOS|8020/3
C0205698|T191|OP|BB18.|RCDSY|Carcinoma, undifferentiated type, NOS|8020/3
C0205698|T191|PT|38549000|SNOMEDCT_US|Carcinoma, undifferentiated|8020/3
C0205698|T191|IS|38549000|SNOMEDCT_US|Carcinoma, undifferentiated, NOS|8020/3
C0205698|T191|SY|38549000|SNOMEDCT_US|Undifferentiated carcinoma|8020/3
C0205696|T191|PT|0000020682|CHV|anaplastic carcinoma|8021/3
C0205696|T191|SY|0000020682|CHV|anaplastic carcinomas|8021/3
C0205696|T191|SY|0000020682|CHV|carcinoma anaplastic|8021/3
C0205698|T191|SY|0000020684|CHV|carcinoma undifferentiated|8021/3
C0205698|T191|PT|0000020684|CHV|undifferentiated carcinoma|8021/3
C0205698|T191|LA|LA15447-8|LNC|Undifferentiated carcinoma|8021/3
C0205696|T191|LLT|10072461|MDR|Anaplastic carcinoma|8021/3
C0205696|T191|PT|271399|MEDCIN|anaplastic carcinoma|8021/3
C0205698|T191|PT|271398|MEDCIN|undifferentiated carcinoma|8021/3
C0205696|T191|PM|D002277|MSH|Anaplastic Carcinoma|8021/3
C0205696|T191|PM|D002277|MSH|Anaplastic Carcinomas|8021/3
C0205696|T191|PEP|D002277|MSH|Carcinoma, Anaplastic|8021/3
C0205698|T191|PEP|D002277|MSH|Carcinoma, Undifferentiated|8021/3
C0205698|T191|PM|D002277|MSH|Undifferentiated Carcinoma|8021/3
C0205698|T191|PM|D002277|MSH|Undifferentiated Carcinomas|8021/3
C0205696|T191|PN|NOCODE|MTH|Anaplastic carcinoma|8021/3
C0205698|T191|PN|NOCODE|MTH|Undifferentiated carcinoma|8021/3
C0205698|T191|SY|C3692|NCI|Anaplastic Carcinoma|8021/3
C0205698|T191|SY|C3692|NCI|Carcinoma, Undifferentiated|8021/3
C0205698|T191|PT|C3692|NCI|Undifferentiated Carcinoma|8021/3
C0205698|T191|SY|TCGA|NCI|Undifferentiated Carcinoma|8021/3
C0205698|T191|SY|C3692|NCI_CDISC|Anaplastic Carcinoma|8021/3
C0205698|T191|SY|C3692|NCI_CDISC|Carcinoma, Undifferentiated|8021/3
C0205698|T191|PT|C3692|NCI_CDISC|CARCINOMA, UNDIFFERENTIATED, MALIGNANT|8021/3
C0205698|T191|PT|C3692|NCI_CPTAC|Undifferentiated Carcinoma|8021/3
C0205696|T191|PT|XM1F7|RCD|Anaplastic carcinoma|8021/3
C0205698|T191|PT|XM1F6|RCD|Undifferentiated carcinoma|8021/3
C0205696|T191|OA|BB19.|RCDSY|Carcinoma, anaplastic NOS|8021/3
C0205696|T191|OP|BB19.|RCDSY|Carcinoma, anaplastic type, NOS|8021/3
C0205698|T191|OA|BB18.|RCDSY|Carcinoma, undiff. type NOS|8021/3
C0205698|T191|OP|BB18.|RCDSY|Carcinoma, undifferentiated type, NOS|8021/3
C0205696|T191|SY|58248003|SNOMEDCT_US|Anaplastic carcinoma|8021/3
C0205696|T191|PT|58248003|SNOMEDCT_US|Carcinoma, anaplastic|8021/3
C0205696|T191|IS|58248003|SNOMEDCT_US|Carcinoma, anaplastic, NOS|8021/3
C0205698|T191|PT|38549000|SNOMEDCT_US|Carcinoma, undifferentiated|8021/3
C0205698|T191|IS|38549000|SNOMEDCT_US|Carcinoma, undifferentiated, NOS|8021/3
C0205698|T191|SY|38549000|SNOMEDCT_US|Undifferentiated carcinoma|8021/3
C0334233|T191|PT|271400|MEDCIN|pleomorphic carcinoma|8022/3
C0334233|T191|PT|C4094|NCI|Pleomorphic Carcinoma|8022/3
C0334233|T191|PT|BB1A.|RCD|Pleomorphic carcinoma|8022/3
C0334233|T191|PT|16741004|SNOMEDCT_US|Pleomorphic carcinoma|8022/3
C0334234|T191|PT|271403|MEDCIN|giant cell and spindle cell carcinoma|8030/3
C0334234|T191|OP|C65160|NCI|Giant Cell and Spindle Cell Carcinoma|8030/3
C0334234|T191|PT|C65160|NCI|Giant Cell and Spindle Cell Carcinoma|8030/3
C0334234|T191|AB|BB1B.|RCD|Giant cell & spindle cell ca|8030/3
C0334234|T191|PT|BB1B.|RCD|Giant cell and spindle cell carcinoma|8030/3
C0334234|T191|PT|72969003|SNOMEDCT_US|Giant cell and spindle cell carcinoma|8030/3
C0206703|T191|PT|271401|MEDCIN|giant cell carcinoma|8031/3
C0206703|T191|MH|D018286|MSH|Carcinoma, Giant Cell|8031/3
C0206703|T191|PM|D018286|MSH|Carcinomas, Giant Cell|8031/3
C0206703|T191|PM|D018286|MSH|Cell Carcinoma, Giant|8031/3
C0206703|T191|PM|D018286|MSH|Cell Carcinomas, Giant|8031/3
C0206703|T191|PM|D018286|MSH|Giant Cell Carcinoma|8031/3
C0206703|T191|PM|D018286|MSH|Giant Cell Carcinomas|8031/3
C0206703|T191|SY|C3779|NCI|Carcinoma, Giant Cell|8031/3
C0206703|T191|PT|C3779|NCI|Giant Cell Carcinoma|8031/3
C0206703|T191|PT|BB1C.|RCD|Giant cell carcinoma|8031/3
C0206703|T191|PT|42596004|SNOMEDCT_US|Giant cell carcinoma|8031/3
C0205697|T191|PT|0000029941|CHV|sarcomatoid carcinoma|8032/3
C0205697|T191|PT|0000020683|CHV|spindle cell carcinoma|8032/3
C0205697|T191|SY|0000020683|CHV|spindle-cell carcinoma|8032/3
C0205697|T191|LA|LA26501-9|LNC|Spindle cell carcinoma, NOS|8032/3
C0205697|T191|LLT|10080324|MDR|Sarcomatoid carcinoma|8032/3
C0205697|T191|PT|10080324|MDR|Sarcomatoid carcinoma|8032/3
C0205697|T191|PT|271404|MEDCIN|pseudosarcomatous carcinoma|8032/3
C0205697|T191|PT|271402|MEDCIN|spindle cell carcinoma|8032/3
C0205697|T191|PM|D002277|MSH|Carcinoma, Spindle Cell|8032/3
C0205697|T191|PEP|D002277|MSH|Carcinoma, Spindle-Cell|8032/3
C0205697|T191|PM|D002277|MSH|Spindle-Cell Carcinoma|8032/3
C0205697|T191|PM|D002277|MSH|Spindle-Cell Carcinomas|8032/3
C0205697|T191|SY|C27004|NCI|Pseudosarcomatous Carcinoma|8032/3
C0205697|T191|PT|C27004|NCI|Sarcomatoid Carcinoma|8032/3
C0205697|T191|SY|TCGA|NCI|Sarcomatoid Carcinoma|8032/3
C0205697|T191|SY|C27004|NCI|Spindle Cell Carcinoma|8032/3
C0205697|T191|PT|C27004|NCI_CDISC|CARCINOMA, SPINDLE CELL, MALIGNANT|8032/3
C0205697|T191|SY|C27004|NCI_CDISC|Pseudosarcomatous Carcinoma|8032/3
C0205697|T191|SY|C27004|NCI_CDISC|Spindle Cell Carcinoma|8032/3
C0205697|T191|PT|C27004|NCI_CPTAC|Sarcomatoid Carcinoma|8032/3
C0205697|T191|PT|CDR0000476767|NCI_NCI-GLOSS|sarcomatoid carcinoma|8032/3
C0205697|T191|PT|BB1E.|RCD|Pseudosarcomatous carcinoma|8032/3
C0205697|T191|PT|BB1D.|RCD|Spindle cell carcinoma|8032/3
C0205697|T191|SY|65692009|SNOMEDCT_US|Polypoid squamous cell carcinoma|8032/3
C0205697|T191|PT|23109009|SNOMEDCT_US|Pseudosarcomatous carcinoma|8032/3
C0205697|T191|SY|23109009|SNOMEDCT_US|Sarcomatoid carcinoma|8032/3
C0205697|T191|PT|65692009|SNOMEDCT_US|Spindle cell carcinoma|8032/3
C0205697|T191|PT|0000029941|CHV|sarcomatoid carcinoma|8033/3
C0205697|T191|PT|0000020683|CHV|spindle cell carcinoma|8033/3
C0205697|T191|SY|0000020683|CHV|spindle-cell carcinoma|8033/3
C0205697|T191|LA|LA26501-9|LNC|Spindle cell carcinoma, NOS|8033/3
C0205697|T191|LLT|10080324|MDR|Sarcomatoid carcinoma|8033/3
C0205697|T191|PT|10080324|MDR|Sarcomatoid carcinoma|8033/3
C0205697|T191|PT|271404|MEDCIN|pseudosarcomatous carcinoma|8033/3
C0205697|T191|PT|271402|MEDCIN|spindle cell carcinoma|8033/3
C0205697|T191|PM|D002277|MSH|Carcinoma, Spindle Cell|8033/3
C0205697|T191|PEP|D002277|MSH|Carcinoma, Spindle-Cell|8033/3
C0205697|T191|PM|D002277|MSH|Spindle-Cell Carcinoma|8033/3
C0205697|T191|PM|D002277|MSH|Spindle-Cell Carcinomas|8033/3
C0205697|T191|SY|C27004|NCI|Pseudosarcomatous Carcinoma|8033/3
C0205697|T191|PT|C27004|NCI|Sarcomatoid Carcinoma|8033/3
C0205697|T191|SY|TCGA|NCI|Sarcomatoid Carcinoma|8033/3
C0205697|T191|SY|C27004|NCI|Spindle Cell Carcinoma|8033/3
C0205697|T191|PT|C27004|NCI_CDISC|CARCINOMA, SPINDLE CELL, MALIGNANT|8033/3
C0205697|T191|SY|C27004|NCI_CDISC|Pseudosarcomatous Carcinoma|8033/3
C0205697|T191|SY|C27004|NCI_CDISC|Spindle Cell Carcinoma|8033/3
C0205697|T191|PT|C27004|NCI_CPTAC|Sarcomatoid Carcinoma|8033/3
C0205697|T191|PT|CDR0000476767|NCI_NCI-GLOSS|sarcomatoid carcinoma|8033/3
C0205697|T191|PT|BB1E.|RCD|Pseudosarcomatous carcinoma|8033/3
C0205697|T191|PT|BB1D.|RCD|Spindle cell carcinoma|8033/3
C0205697|T191|SY|65692009|SNOMEDCT_US|Polypoid squamous cell carcinoma|8033/3
C0205697|T191|PT|23109009|SNOMEDCT_US|Pseudosarcomatous carcinoma|8033/3
C0205697|T191|SY|23109009|SNOMEDCT_US|Sarcomatoid carcinoma|8033/3
C0205697|T191|PT|65692009|SNOMEDCT_US|Spindle cell carcinoma|8033/3
C0334236|T191|PT|271405|MEDCIN|polygonal cell carcinoma|8034/3
C0334236|T191|OP|C65161|NCI|Polygonal Cell Carcinoma|8034/3
C0334236|T191|PT|C65161|NCI|Polygonal Cell Carcinoma|8034/3
C0334236|T191|PT|BB1F.|RCD|Polygonal cell carcinoma|8034/3
C0334236|T191|PT|70401000|SNOMEDCT_US|Polygonal cell carcinoma|8034/3
C1266000|T191|PT|271406|MEDCIN|carcinoma with osteoclast-like giant cells|8035/3
C1266000|T191|SY|271406|MEDCIN|malignant neoplasm carcinoma w/ osteoclast-like giant cells|8035/3
C1883424|T191|PT|C63622|NCI|Undifferentiated Carcinoma with Osteoclast-Like Giant Cells|8035/3
C1883424|T191|SY|TCGA|NCI|Undifferentiated Carcinoma with Osteoclast-Like Giant Cells|8035/3
C1266000|T191|PT|128631001|SNOMEDCT_US|Carcinoma with osteoclast-like giant cells|8035/3
C0334237|T191|SY|C65162|NCI|Benign Tumorlet|8040/0
C0334237|T191|PT|C65162|NCI|Tumorlet|8040/0
C0334237|T191|PT|BB1H.|RCD|Tumourlet|8040/0
C0334237|T191|PT|72938002|SNOMEDCT_US|Tumorlet|8040/0
C1266001|T191|PT|128876004|SNOMEDCT_US|Tumorlet, benign|8040/0
C0334237|T191|PTGB|72938002|SNOMEDCT_US|Tumourlet|8040/0
C1266001|T191|PTGB|128876004|SNOMEDCT_US|Tumourlet, benign|8040/0
C0334237|T191|SY|C65162|NCI|Benign Tumorlet|8040/1
C0334237|T191|PT|C65162|NCI|Tumorlet|8040/1
C0334237|T191|PT|BB1H.|RCD|Tumourlet|8040/1
C0334237|T191|PT|72938002|SNOMEDCT_US|Tumorlet|8040/1
C0334237|T191|PTGB|72938002|SNOMEDCT_US|Tumourlet|8040/1
C0262584|T191|PT|0000025445|CHV|oat cell carcinoma|8041/3
C0262584|T191|ET|2017-6589|CSP|oat cell carcinoma|8041/3
C0262584|T191|LA|LA26101-8|LNC|Small cell neuroendocrine carcinoma|8041/3
C0262584|T191|LLT|10029882|MDR|Oat cell carcinoma|8041/3
C0262584|T191|LLT|10041056|MDR|Small cell carcinoma|8041/3
C0262584|T191|PT|10041056|MDR|Small cell carcinoma|8041/3
C1275215|T191|SY|357596|MEDCIN|skin neoplasm malignant adnexa with eccrine differentiation small cell carcinoma|8041/3
C0262584|T191|PT|271407|MEDCIN|small cell carcinoma|8041/3
C1275215|T191|PT|357596|MEDCIN|Small cell eccrine carcinoma of skin|8041/3
C0262584|T191|ET|D018288|MSH|Carcinoma, Oat Cell|8041/3
C0262584|T191|MH|D018288|MSH|Carcinoma, Small Cell|8041/3
C0262584|T191|PM|D018288|MSH|Carcinomas, Oat Cell|8041/3
C0262584|T191|PM|D018288|MSH|Carcinomas, Small Cell|8041/3
C0262584|T191|ET|D018288|MSH|Oat Cell Carcinoma|8041/3
C0262584|T191|PM|D018288|MSH|Oat Cell Carcinomas|8041/3
C0262584|T191|DEV|D018288|MSH|SCLC|8041/3
C0262584|T191|ET|D018288|MSH|Small Cell Carcinoma|8041/3
C0262584|T191|PM|D018288|MSH|Small Cell Carcinomas|8041/3
C0262584|T191|PN|NOCODE|MTH|Carcinoma, Small Cell|8041/3
C0262584|T191|OP|C3915|NCI|Oat Cell Cancer|8041/3
C0262584|T191|OP|C3915|NCI|Oat Cell Carcinoma|8041/3
C0262584|T191|SY|C3915|NCI|Small Cell Cancer|8041/3
C0262584|T191|PT|C3915|NCI|Small Cell Carcinoma|8041/3
C0262584|T191|SY|TCGA|NCI|Small Cell Carcinoma|8041/3
C0262584|T191|SY|C3915|NCI|Small Cell NEC|8041/3
C0262584|T191|SY|C3915|NCI|Small Cell Neuroendocrine Carcinoma|8041/3
C0262584|T191|DN|C3915|NCI_CTRP|Small Cell Carcinoma|8041/3
C0262584|T191|PT|CDR0000046256|NCI_NCI-GLOSS|oat cell cancer|8041/3
C0262584|T191|PT|BB1K.|RCD|Oat cell carcinoma|8041/3
C0262584|T191|SY|Xa989|RCD|Reserve cell carcinoma|8041/3
C0262584|T191|SY|Xa989|RCD|Round cell carcinoma|8041/3
C0262584|T191|SY|Xa989|RCD|SCC - Small cell carcinoma|8041/3
C0262584|T191|PT|Xa989|RCD|Small cell carcinoma|8041/3
C0262584|T191|OP|BB1J.|RCDSY|Small cell carcinoma NOS|8041/3
C0262584|T191|PT|76817009|SNOMEDCT_US|Oat cell carcinoma|8041/3
C0262584|T191|SY|74364000|SNOMEDCT_US|Reserve cell carcinoma|8041/3
C0262584|T191|SY|74364000|SNOMEDCT_US|Round cell carcinoma|8041/3
C0262584|T191|SY|74364000|SNOMEDCT_US|SCC - Small cell carcinoma|8041/3
C0262584|T191|PT|11010461000119101|SNOMEDCT_US|Small cell carcinoma|8041/3
C0262584|T191|PT|74364000|SNOMEDCT_US|Small cell carcinoma|8041/3
C0262584|T191|IS|74364000|SNOMEDCT_US|Small cell carcinoma, NOS|8041/3
C1275215|T191|PT|403944002|SNOMEDCT_US|Small cell eccrine carcinoma|8041/3
C1275215|T191|PT|400134004|SNOMEDCT_US|Small cell eccrine carcinoma|8041/3
C1275215|T191|SY|403944002|SNOMEDCT_US|Small cell eccrine carcinoma of skin|8041/3
C0262584|T191|IS|74364000|SNOMEDCT_US|Small cell neuroendocrine carcinoma|8041/3
C0262584|T191|PT|719105002|SNOMEDCT_US|Small cell neuroendocrine carcinoma|8041/3
C0262584|T191|PT|0000025445|CHV|oat cell carcinoma|8042/3
C0262584|T191|ET|2017-6589|CSP|oat cell carcinoma|8042/3
C0262584|T191|LA|LA26101-8|LNC|Small cell neuroendocrine carcinoma|8042/3
C0262584|T191|LLT|10029882|MDR|Oat cell carcinoma|8042/3
C0262584|T191|LLT|10041056|MDR|Small cell carcinoma|8042/3
C0262584|T191|PT|10041056|MDR|Small cell carcinoma|8042/3
C0262584|T191|PT|271407|MEDCIN|small cell carcinoma|8042/3
C0262584|T191|ET|D018288|MSH|Carcinoma, Oat Cell|8042/3
C0262584|T191|MH|D018288|MSH|Carcinoma, Small Cell|8042/3
C0262584|T191|PM|D018288|MSH|Carcinomas, Oat Cell|8042/3
C0262584|T191|PM|D018288|MSH|Carcinomas, Small Cell|8042/3
C0262584|T191|ET|D018288|MSH|Oat Cell Carcinoma|8042/3
C0262584|T191|PM|D018288|MSH|Oat Cell Carcinomas|8042/3
C0262584|T191|DEV|D018288|MSH|SCLC|8042/3
C0262584|T191|ET|D018288|MSH|Small Cell Carcinoma|8042/3
C0262584|T191|PM|D018288|MSH|Small Cell Carcinomas|8042/3
C0262584|T191|PN|NOCODE|MTH|Carcinoma, Small Cell|8042/3
C0262584|T191|OP|C3915|NCI|Oat Cell Cancer|8042/3
C0262584|T191|OP|C3915|NCI|Oat Cell Carcinoma|8042/3
C0262584|T191|SY|C3915|NCI|Small Cell Cancer|8042/3
C0262584|T191|PT|C3915|NCI|Small Cell Carcinoma|8042/3
C0262584|T191|SY|TCGA|NCI|Small Cell Carcinoma|8042/3
C0262584|T191|SY|C3915|NCI|Small Cell NEC|8042/3
C0262584|T191|SY|C3915|NCI|Small Cell Neuroendocrine Carcinoma|8042/3
C0262584|T191|DN|C3915|NCI_CTRP|Small Cell Carcinoma|8042/3
C0262584|T191|PT|CDR0000046256|NCI_NCI-GLOSS|oat cell cancer|8042/3
C0262584|T191|PT|BB1K.|RCD|Oat cell carcinoma|8042/3
C0262584|T191|SY|Xa989|RCD|Reserve cell carcinoma|8042/3
C0262584|T191|SY|Xa989|RCD|Round cell carcinoma|8042/3
C0262584|T191|SY|Xa989|RCD|SCC - Small cell carcinoma|8042/3
C0262584|T191|PT|Xa989|RCD|Small cell carcinoma|8042/3
C0262584|T191|OP|BB1J.|RCDSY|Small cell carcinoma NOS|8042/3
C0262584|T191|PT|76817009|SNOMEDCT_US|Oat cell carcinoma|8042/3
C0262584|T191|SY|74364000|SNOMEDCT_US|Reserve cell carcinoma|8042/3
C0262584|T191|SY|74364000|SNOMEDCT_US|Round cell carcinoma|8042/3
C0262584|T191|SY|74364000|SNOMEDCT_US|SCC - Small cell carcinoma|8042/3
C0262584|T191|PT|11010461000119101|SNOMEDCT_US|Small cell carcinoma|8042/3
C0262584|T191|PT|74364000|SNOMEDCT_US|Small cell carcinoma|8042/3
C0262584|T191|IS|74364000|SNOMEDCT_US|Small cell carcinoma, NOS|8042/3
C0262584|T191|IS|74364000|SNOMEDCT_US|Small cell neuroendocrine carcinoma|8042/3
C0262584|T191|PT|719105002|SNOMEDCT_US|Small cell neuroendocrine carcinoma|8042/3
C0334238|T191|PT|271408|MEDCIN|fusiform type small cell carcinoma|8043/3
C0334238|T191|SY|271408|MEDCIN|small cell carcinoma, fusiform cell|8043/3
C0334238|T191|OP|C27092|NCI|Small Cell Carcinoma, Fusiform Cell Type|8043/3
C0334238|T191|PT|C27092|NCI|Small Cell Carcinoma, Fusiform Cell Type|8043/3
C0334238|T191|DN|C27092|NCI_CTRP|Small Cell Cancer, Fusiform Cell Type|8043/3
C0334238|T191|SY|CDR0000039857|PDQ|fusiform type SCLC|8043/3
C0334238|T191|PT|CDR0000039857|PDQ|fusiform type small cell lung cancer|8043/3
C0334238|T191|SY|CDR0000039857|PDQ|lung cancer, fusiform type, small cell|8043/3
C0334238|T191|SY|CDR0000039857|PDQ|SCLC, fusiform type|8043/3
C0334238|T191|IS|CDR0000039857|PDQ|Small Cell Carcinoma, Fusiform Cell Type|8043/3
C0334238|T191|SY|CDR0000039857|PDQ|small cell lung cancer, fusiform type|8043/3
C0334238|T191|AB|BB1L.|RCD|Small cell ca - fusiform cell|8043/3
C0334238|T191|PT|BB1L.|RCD|Small cell carcinoma - fusiform cell|8043/3
C0334238|T191|SY|74042001|SNOMEDCT_US|Small cell carcinoma - fusiform cell|8043/3
C0334238|T191|PT|74042001|SNOMEDCT_US|Small cell carcinoma, fusiform cell|8043/3
C0334239|T191|PT|MTHU014783|ICPC2ICD10ENG|carcinoma; small cell, with intermediate cell, unspecified site|8044/3
C0334239|T191|PT|MTHU041503|ICPC2ICD10ENG|small cell; carcinoma, with intermediate cell, unspecified site|8044/3
C0334239|T191|OP|C4099|NCI|Small Cell Carcinoma, Intermediate Cell|8044/3
C0334239|T191|OP|C4099|NCI|Small Cell Intermediate Cell Carcinoma|8044/3
C0334239|T191|PT|C4099|NCI|Small Cell Intermediate Cell Carcinoma|8044/3
C0334239|T191|DN|C4099|NCI_CTRP|Small Cell Cancer, Intermediate Cell Type|8044/3
C0334239|T191|SY|CDR0000039855|PDQ|intermediate type SCLC|8044/3
C0334239|T191|PT|CDR0000039855|PDQ|intermediate type small cell lung cancer|8044/3
C0334239|T191|SY|CDR0000039855|PDQ|lung cancer, intermediate type, small cell|8044/3
C0334239|T191|SY|CDR0000039855|PDQ|SCLC, intermediate type|8044/3
C0334239|T191|SY|CDR0000039855|PDQ|Small Cell Carcinoma, Intermediate Cell|8044/3
C0334239|T191|IS|CDR0000039855|PDQ|Small Cell Intermediate Cell Carcinoma|8044/3
C0334239|T191|SY|CDR0000039855|PDQ|small cell lung cancer, intermediate type|8044/3
C0334239|T191|AB|X77mv|RCD|Small cell ca - intermed cell|8044/3
C0334239|T191|PT|X77mv|RCD|Small cell carcinoma - intermediate cell|8044/3
C0334239|T191|AB|X77mv|RCDSY|Small cell carc, interm cel|8044/3
C0334239|T191|SY|X77mv|RCDSY|Small cell carcinoma, intermediate cell|8044/3
C0334239|T191|OAP|189557009|SNOMEDCT_US|Small cell carcinoma - intermediate cell|8044/3
C0334239|T191|OF|189557009|SNOMEDCT_US|Small cell carcinoma - intermediate cell|8044/3
C3839982|T191|PTGB|703549009|SNOMEDCT_US|Small cell carcinoma, hypercalcaemic type|8044/3
C3839982|T191|PT|703549009|SNOMEDCT_US|Small cell carcinoma, hypercalcemic type|8044/3
C0334239|T191|PT|5958006|SNOMEDCT_US|Small cell carcinoma, intermediate cell|8044/3
C1333125|T191|PT|219590|MEDCIN|combined small cell carcinoma of lung|8045/3
C1333125|T191|PT|C9137|NCI|Combined Lung Small Cell Carcinoma|8045/3
C1333125|T191|SY|C9137|NCI|Combined Small and Large Cell Lung Cancer|8045/3
C1333125|T191|SY|C9137|NCI|Combined Small and Large Cell Lung Carcinoma|8045/3
C1333125|T191|SY|C9137|NCI|Combined Small Cell and Large Cell Lung Carcinoma|8045/3
C1333125|T191|SY|C9137|NCI|Combined Small Cell Carcinoma of Lung|8045/3
C1333125|T191|SY|C9137|NCI|Combined Small Cell Carcinoma of the Lung|8045/3
C1333125|T191|SY|C9137|NCI|Combined Small Cell Lung Carcinoma|8045/3
C1333125|T191|SY|C9137|NCI|Combined Type Small Cell Carcinoma of Lung|8045/3
C1333125|T191|SY|C9137|NCI|Combined Type Small Cell Carcinoma of the Lung|8045/3
C1333125|T191|SY|C9137|NCI|Combined Type Small Cell Lung Carcinoma|8045/3
C1333125|T191|SY|C9137|NCI|Mixed Small Cell and Large Cell Carcinoma of Lung|8045/3
C1333125|T191|SY|C9137|NCI|Mixed Small Cell and Large Cell Carcinoma of the Lung|8045/3
C1333125|T191|SY|C9137|NCI|Mixed Small Cell and Large Cell Lung Carcinoma|8045/3
C1333125|T191|SY|C9137|NCI|Small Cell and Large Cell Carcinoma of Lung|8045/3
C1333125|T191|SY|C9137|NCI|Small Cell and Large Cell Carcinoma of the Lung|8045/3
C1333125|T191|SY|C9137|NCI|Small Cell and Large Cell Lung Carcinoma|8045/3
C1333125|T191|DN|C9137|NCI_CTRP|Combined Small Cell Lung Cancer|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Small and Large Cell Lung Cancer|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Small and Large Cell Lung Carcinoma|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Small Cell and Large Cell Lung Carcinoma|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Small Cell Carcinoma of Lung|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Small Cell Carcinoma of the Lung|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Small Cell Lung Carcinoma|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|combined type SCLC|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Type Small Cell Carcinoma of Lung|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Type Small Cell Carcinoma of the Lung|8045/3
C1333125|T191|PT|CDR0000039858|PDQ|combined type small cell lung cancer|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Combined Type Small Cell Lung Carcinoma|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|lung cancer, combined type, small cell|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Mixed Small Cell and Large Cell Carcinoma of Lung|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Mixed Small Cell and Large Cell Carcinoma of the Lung|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Mixed Small Cell and Large Cell Lung Carcinoma|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|SCLC, combined type|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Small Cell and Large Cell Carcinoma of Lung|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Small Cell and Large Cell Carcinoma of the Lung|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|Small Cell and Large Cell Lung Carcinoma|8045/3
C1333125|T191|SY|CDR0000039858|PDQ|small cell lung cancer, combined type|8045/3
C0334240|T191|AB|X77mw|RCD|Small cell - large cell ca|8045/3
C0334240|T191|PT|X77mw|RCD|Small cell - large cell carcinoma|8045/3
C0334240|T191|AB|X77mw|RCDSY|Small cell-large cell carc|8045/3
C0334240|T191|SY|X77mw|RCDSY|Small cell-large cell carcinoma|8045/3
C0334240|T191|PT|21326004|SNOMEDCT_US|Combined small cell carcinoma|8045/3
C0334240|T191|SY|21326004|SNOMEDCT_US|Combined small cell-adenocarcinoma|8045/3
C0334240|T191|SY|21326004|SNOMEDCT_US|Combined small cell-squamous cell carcinoma|8045/3
C0334240|T191|SY|21326004|SNOMEDCT_US|Mixed small cell carcinoma|8045/3
C4518201|T191|PT|733844008|SNOMEDCT_US|Neuroendocrine type combined small cell carcinoma|8045/3
C0334240|T191|OAP|189558004|SNOMEDCT_US|Small cell - large cell carcinoma|8045/3
C0334240|T191|OF|189558004|SNOMEDCT_US|Small cell - large cell carcinoma|8045/3
C0334240|T191|SY|21326004|SNOMEDCT_US|Small cell-large cell carcinoma|8045/3
C1266002|T191|SY|0000056675|CHV|non small cell carcinoma|8046/3
C1266002|T191|PT|0000056675|CHV|non-small cell carcinoma|8046/3
C1266002|T191|SY|0000056675|CHV|small cell carcinoma non|8046/3
C1266002|T191|PT|C65151|NCI|Non-Small Cell Carcinoma|8046/3
C1266002|T191|SY|TCGA|NCI|Non-Small Cell Carcinoma|8046/3
C1266002|T191|PT|C65151|NCI_CPTAC|Non-Small Cell Carcinoma|8046/3
C1266002|T191|PT|128632008|SNOMEDCT_US|Non-small cell carcinoma|8046/3
C0030354|T191|DE|0000004529|AOD|papilloma|8050/0
C0030354|T191|PT|0044946|CCPSS|PAPILLOMA|8050/0
C0030354|T191|PT|0000009247|CHV|non cancerous skin tumor|8050/0
C0030354|T191|SY|0000009247|CHV|papilloma|8050/0
C0030354|T191|SY|0000009247|CHV|papillomas|8050/0
C0030354|T191|SY|0000009247|CHV|papillomata|8050/0
C0030354|T191|PT|U000505|COSTAR|PAPILLOMA|8050/0
C0030354|T191|FI|U003008|DXP|PAPILLOMA|8050/0
C0030354|T191|PT|HP:0012740|HPO|Papilloma|8050/0
C0030354|T191|PT|U003462|LCH|Papilloma|8050/0
C0030354|T191|PT|sh85097677|LCH_NW|Papilloma|8050/0
C0030354|T191|LLT|10033713|MDR|Papilloma|8050/0
C0030354|T191|PT|10033713|MDR|Papilloma|8050/0
C0030354|T191|LLT|10033715|MDR|Papilloma NOS|8050/0
C0030354|T191|LLT|10033725|MDR|Papillomata|8050/0
C0030354|T191|PT|6231|MEDCIN|papilloma|8050/0
C0030354|T191|MH|D010212|MSH|Papilloma|8050/0
C0030354|T191|PM|D010212|MSH|Papillomas|8050/0
C0030354|T191|PN|NOCODE|MTH|Papilloma|8050/0
C0030354|T191|PT|C7440|NCI|Papilloma|8050/0
C0030354|T191|PT|C7440|NCI_CDISC|PAPILLOMA, BENIGN|8050/0
C0030354|T191|PT|X77n9|RCD|Papilloma|8050/0
C0030354|T191|PT|711329002|SNOMEDCT_US|Papilloma|8050/0
C0030354|T191|SY|23730008|SNOMEDCT_US|Papilloma|8050/0
C0030354|T191|IS|23730008|SNOMEDCT_US|Papilloma, NOS|8050/0
C0030354|T191|PT|1486|WHO|PAPILLOMA|8050/0
C0334242|T191|PT|271380|MEDCIN|papillary carcinoma in situ|8050/2
C0334242|T191|PN|NOCODE|MTH|Papillary carcinoma in situ|8050/2
C0334242|T191|PT|C65163|NCI|Papillary Carcinoma In Situ|8050/2
C0334242|T191|PT|BB21.|RCD|Papillary carcinoma in situ|8050/2
C0334242|T191|PT|10376009|SNOMEDCT_US|Papillary carcinoma in situ|8050/2
C0007133|T191|SY|0000002434|CHV|carcinoma papillary|8050/3
C0007133|T191|PT|0000002434|CHV|papillary carcinoma|8050/3
C0007133|T191|SY|0000002434|CHV|papillary carcinomas|8050/3
C0007133|T191|PT|271409|MEDCIN|papillary carcinoma|8050/3
C0007133|T191|MH|D002291|MSH|Carcinoma, Papillary|8050/3
C0007133|T191|PM|D002291|MSH|Carcinomas, Papillary|8050/3
C0007133|T191|PM|D002291|MSH|Papillary Carcinoma|8050/3
C0007133|T191|PM|D002291|MSH|Papillary Carcinomas|8050/3
C0007133|T191|PT|C2927|NCI|Papillary Carcinoma|8050/3
C0007133|T191|SY|TCGA|NCI|Papillary Carcinoma|8050/3
C0007133|T191|PT|C2927|NCI_CPTAC|Papillary Carcinoma|8050/3
C0007133|T191|PT|Xa98A|RCD|Papillary carcinoma|8050/3
C0007133|T191|OP|BB22.|RCDSY|Papillary carcinoma NOS|8050/3
C0007133|T191|PT|25910003|SNOMEDCT_US|Papillary carcinoma|8050/3
C1720430|T191|PT|421630008|SNOMEDCT_US|Papillary carcinoma, clear cell|8050/3
C1720274|T191|PT|422238009|SNOMEDCT_US|Papillary carcinoma, cribriform-morular|8050/3
C1720126|T191|PT|421414006|SNOMEDCT_US|Papillary carcinoma, macrofollicular|8050/3
C0007133|T191|IS|25910003|SNOMEDCT_US|Papillary carcinoma, NOS|8050/3
C1719884|T191|SYGB|421980000|SNOMEDCT_US|Papillary carcinoma, radiation-induced paediatric variant|8050/3
C1719884|T191|SY|421980000|SNOMEDCT_US|Papillary carcinoma, radiation-induced pediatric variant|8050/3
C1719884|T191|PT|421980000|SNOMEDCT_US|Papillary carcinoma, solid|8050/3
C1720441|T191|PT|421658000|SNOMEDCT_US|Papillary carcinoma, Warthin-like|8050/3
C0302180|T047|PT|0059444|CCPSS|CONDYLOMA|8051/0
C0302180|T047|PT|0000027927|CHV|condyloma|8051/0
C0302180|T047|SY|0000027927|CHV|condylomas|8051/0
C0302180|T047|SY|0000027927|CHV|condylomata|8051/0
C0302180|T047|PT|U000197|COSTAR|CONDYLOMATA|8051/0
C0302180|T047|ET|2020-4312|CSP|condyloma|8051/0
C0302180|T047|PT|MTHU018427|ICPC2ICD10ENG|condyloma|8051/0
C0302180|T047|LLT|10053433|MDR|Condyloma|8051/0
C0302180|T047|PN|NOCODE|MTH|Condyloma|8051/0
C0302180|T047|ET|078.11|MTHICD9|Condyloma NOS|8051/0
C0334243|T191|PT|C4101|NCI|Verrucous Papilloma|8051/0
C0334243|T191|OP|C4101|NCI|Verrucous Papilloma|8051/0
C0334243|T191|PT|BB23.|RCD|Verrucous papilloma|8051/0
C0302180|T047|PT|19672005|SNOMEDCT_US|Condyloma|8051/0
C0302180|T047|IS|19672005|SNOMEDCT_US|Condyloma, NOS|8051/0
C0334243|T191|PT|48218007|SNOMEDCT_US|Verrucous papilloma|8051/0
C0206706|T191|SY|0000021035|CHV|carcinoma verrucous|8051/3
C0206706|T191|PT|0000021035|CHV|verrucous carcinoma|8051/3
C0206706|T191|SY|0000021035|CHV|verrucous carcinomas|8051/3
C0206706|T191|PT|351487|MEDCIN|squamous cell carcinoma verrucous|8051/3
C0206706|T191|PT|271411|MEDCIN|verrucous carcinoma|8051/3
C0206706|T191|MH|D018289|MSH|Carcinoma, Verrucous|8051/3
C0206706|T191|PM|D018289|MSH|Carcinomas, Verrucous|8051/3
C0206706|T191|PM|D018289|MSH|Verrucous Carcinoma|8051/3
C0206706|T191|PM|D018289|MSH|Verrucous Carcinomas|8051/3
C3251817|T191|PN|NOCODE|MTH|Condylomatous carcinoma|8051/3
C0206706|T191|PN|NOCODE|MTH|Verrucous carcinoma|8051/3
C0206706|T191|PT|C3781|NCI|Verrucous Carcinoma|8051/3
C0206706|T191|SY|C3781|NCI|Verrucous Epidermoid Carcinoma|8051/3
C0206706|T191|SY|C3781|NCI|Verrucous Epidermoid Cell Carcinoma|8051/3
C0206706|T191|SY|C3781|NCI|Verrucous Squamous Carcinoma|8051/3
C0206706|T191|SY|C3781|NCI|Verrucous Squamous Cell Carcinoma|8051/3
C0206706|T191|SY|Xa98B|RCD|SCC - Verrucous squamous cell carcinoma|8051/3
C0206706|T191|PT|Xa98B|RCD|Verrucous carcinoma|8051/3
C0206706|T191|SY|Xa98B|RCD|Verrucous epidermoid carcinoma|8051/3
C0206706|T191|AB|Xa98B|RCD|Verrucous SCC|8051/3
C0206706|T191|AB|Xa98B|RCD|Verrucous squamous cell ca|8051/3
C0206706|T191|SY|Xa98B|RCD|Verrucous squamous cell carcinoma|8051/3
C0206706|T191|OP|BB24.|RCDSY|Verrucous carcinoma NOS|8051/3
C0206706|T191|SY|89906000|SNOMEDCT_US|Condylomatous carcinoma|8051/3
C3251817|T191|SY|399408005|SNOMEDCT_US|Condylomatous carcinoma|8051/3
C0206706|T191|SY|89906000|SNOMEDCT_US|SCC - Verrucous squamous cell carcinoma|8051/3
C0206706|T191|PT|89906000|SNOMEDCT_US|Verrucous carcinoma|8051/3
C0206706|T191|IS|89906000|SNOMEDCT_US|Verrucous carcinoma, NOS|8051/3
C0206706|T191|SY|89906000|SNOMEDCT_US|Verrucous epidermoid carcinoma|8051/3
C0206706|T191|SY|403904009|SNOMEDCT_US|Verrucous epidermoid carcinoma|8051/3
C0206706|T191|PT|403904009|SNOMEDCT_US|Verrucous squamous cell carcinoma|8051/3
C0206706|T191|SY|89906000|SNOMEDCT_US|Verrucous squamous cell carcinoma|8051/3
C3251817|T191|SY|399408005|SNOMEDCT_US|Warty carcinoma|8051/3
C0206706|T191|SY|89906000|SNOMEDCT_US|Warty carcinoma|8051/3
C0205874|T191|SY|0000020738|CHV|cells papilloma squamous|8052/0
C0205874|T191|SY|0000020738|CHV|papillomas squamous|8052/0
C0205874|T191|SY|0000020738|CHV|squamous cell papilloma|8052/0
C0205874|T191|PT|0000020738|CHV|squamous papilloma|8052/0
C0205874|T191|PT|HP:0031021|HPO|Squamous Papilloma|8052/0
C0205874|T191|LLT|10081692|MDR|Squamous cell papilloma|8052/0
C0205874|T191|PEP|D010212|MSH|Papilloma, Squamous Cell|8052/0
C0205874|T191|PM|D010212|MSH|Papillomas, Squamous Cell|8052/0
C0205874|T191|PM|D010212|MSH|Squamous Cell Papilloma|8052/0
C0205874|T191|PM|D010212|MSH|Squamous Cell Papillomas|8052/0
C0205874|T191|SY|C3712|NCI|Epidermoid Cell Papilloma|8052/0
C0205874|T191|SY|C3712|NCI|Epidermoid Papilloma|8052/0
C0205874|T191|SY|C3712|NCI|Keratotic Papilloma|8052/0
C0205874|T191|PT|C3712|NCI|Squamous Cell Papilloma|8052/0
C0205874|T191|SY|C3712|NCI|Squamous Papilloma|8052/0
C0205874|T191|SY|C3712|NCI_CDISC|Epidermoid Cell Papilloma|8052/0
C0205874|T191|SY|C3712|NCI_CDISC|Epidermoid Papilloma|8052/0
C0205874|T191|SY|C3712|NCI_CDISC|Keratotic Papilloma|8052/0
C0205874|T191|PT|C3712|NCI_CDISC|PAPILLOMA, SQUAMOUS CELL, BENIGN|8052/0
C0205874|T191|SY|C3712|NCI_CDISC|Squamous Cell Papilloma|8052/0
C0205874|T191|SY|BB25.|RCD|Keratotic papilloma|8052/0
C0205874|T191|PT|BB25.|RCD|Squamous cell papilloma|8052/0
C0205874|T191|SY|BB25.|RCD|Squamous papilloma|8052/0
C0205874|T191|SY|63451008|SNOMEDCT_US|Keratotic papilloma|8052/0
C0205874|T191|PT|63451008|SNOMEDCT_US|Squamous cell papilloma|8052/0
C0205874|T191|SY|63451008|SNOMEDCT_US|Squamous papilloma|8052/0
C1266003|T191|PT|C65164|NCI|Non-Invasive Papillary Squamous Cell Carcinoma|8052/2
C1266003|T191|SY|128647004|SNOMEDCT_US|Papillary squamous cell carcinoma in situ|8052/2
C1266003|T191|PT|128647004|SNOMEDCT_US|Papillary squamous cell carcinoma, non-invasive|8052/2
C0334244|T191|PT|271410|MEDCIN|papillary squamous cell carcinoma|8052/3
C0334244|T191|SY|C4102|NCI|Papillary Epidermoid Carcinoma|8052/3
C0334244|T191|SY|C4102|NCI|Papillary Epidermoid Cell Carcinoma|8052/3
C0334244|T191|SY|C4102|NCI|Papillary Squamous Carcinoma|8052/3
C0334244|T191|PT|C4102|NCI|Papillary Squamous Cell Carcinoma|8052/3
C0334244|T191|SY|TCGA|NCI|Papillary Squamous Cell Carcinoma|8052/3
C0334244|T191|SY|BB26.|RCD|Papillary epidermoid carcinoma|8052/3
C0334244|T191|AB|BB26.|RCD|Papillary squamous cell ca|8052/3
C0334244|T191|PT|BB26.|RCD|Papillary squamous cell carcinoma|8052/3
C0334244|T191|SY|39056008|SNOMEDCT_US|Papillary epidermoid carcinoma|8052/3
C0334244|T191|PT|39056008|SNOMEDCT_US|Papillary squamous cell carcinoma|8052/3
C1881254|T191|PN|NOCODE|MTH|Inverted Squamous Cell Papilloma|8053/0
C1881254|T191|PT|C65165|NCI|Inverted Squamous Cell Papilloma|8053/0
C1881254|T191|SY|90121000|SNOMEDCT_US|Inverted papilloma|8053/0
C1881254|T191|SY|90121000|SNOMEDCT_US|Inverted papilloma, squamous cell|8053/0
C1881254|T191|PT|90121000|SNOMEDCT_US|Squamous cell papilloma, inverted|8053/0
C1378340|T191|PT|C9009|NCI|Squamous Papillomatosis|8060/0
C1378340|T191|SY|82049002|SNOMEDCT_US|Papillomatosis, squamous|8060/0
C1378340|T191|PT|82049002|SNOMEDCT_US|Squamous papillomatosis|8060/0
C0334245|T191|SY|0000029942|CHV|carcinoma squamous cell in situ|8070/2
C0334245|T191|SY|0000029942|CHV|in situ squamous cell carcinoma|8070/2
C0334245|T191|PT|0000029942|CHV|squamous cell carcinoma in situ|8070/2
C0334245|T191|LLT|10022739|MDR|Intra-epidermal carcinoma|8070/2
C0334245|T191|LLT|10022782|MDR|Intraepidermal carcinoma|8070/2
C0334245|T191|PT|271382|MEDCIN|squamous cell carcinoma in situ|8070/2
C0334245|T191|PN|NOCODE|MTH|Intraepithelial Squamous Cell Carcinoma|8070/2
C0334245|T191|SY|C27093|NCI|Epidermoid Carcinoma in situ|8070/2
C0334245|T191|SY|C27093|NCI|Epidermoid Cell Carcinoma in situ|8070/2
C0334245|T191|AB|C27093|NCI|Grade 3 SIN|8070/2
C0334245|T191|SY|C27093|NCI|Grade 3 Squamous Intraepithelial Neoplasia|8070/2
C0334245|T191|AB|C27093|NCI|Grade III SIN|8070/2
C0334245|T191|SY|C27093|NCI|Grade III Squamous Intraepithelial Neoplasia|8070/2
C0334245|T191|SY|C27093|NCI|Intraepithelial Squamous Cell Carcinoma|8070/2
C0334245|T191|SY|C27093|NCI|Squamous Carcinoma in situ|8070/2
C0334245|T191|SY|C27093|NCI|Squamous Cell Carcinoma in situ|8070/2
C0334245|T191|SY|C27093|NCI|Squamous Cell Carcinoma in-situ|8070/2
C0334245|T191|PT|C27093|NCI|Stage 0 Squamous Cell Carcinoma|8070/2
C0334245|T191|PT|C27093|NCI_CDISC|CARCINOMA, SQUAMOUS CELL, IN SITU, MALIGNANT|8070/2
C0334245|T191|SY|C27093|NCI_CDISC|Epidermoid Carcinoma In situ|8070/2
C0334245|T191|SY|C27093|NCI_CDISC|Epidermoid Cell Carcinoma In situ|8070/2
C0334245|T191|SY|C27093|NCI_CDISC|Grade 3 Squamous Intraepithelial Neoplasia|8070/2
C0334245|T191|SY|C27093|NCI_CDISC|Grade III Squamous Intraepithelial Neoplasia|8070/2
C0334245|T191|SY|C27093|NCI_CDISC|Intraepithelial Squamous Cell Carcinoma|8070/2
C0334245|T191|SY|C27093|NCI_CDISC|Squamous Carcinoma In situ|8070/2
C0334245|T191|SY|C27093|NCI_CDISC|Squamous Cell Carcinoma In situ|8070/2
C0334245|T191|SY|Xa98D|RCD|Epidermoid carcinoma in situ|8070/2
C0334245|T191|SY|Xa98D|RCD|IEC - Intraepidermal carcinoma|8070/2
C0334245|T191|SY|Xa98D|RCD|Intraepidermal carcinoma|8070/2
C0334245|T191|AB|Xa98D|RCD|Intraepithel squamous cell ca|8070/2
C0334245|T191|SY|Xa98D|RCD|Intraepithelial squamous cell carcinoma|8070/2
C0334245|T191|PT|X77n1|RCD|Squamous carcinoma in situ|8070/2
C0334245|T191|AB|Xa98D|RCD|Squamous cell ca in situ|8070/2
C0334245|T191|PT|Xa98D|RCD|Squamous cell carcinoma in situ|8070/2
C0334245|T191|AB|Xa98D|RCDSY|Squam cell ca-in-situ NOS|8070/2
C0334245|T191|SY|Xa98D|RCDSY|Squamous cell carcinoma in situ NOS|8070/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Epidermoid carcinoma in situ|8070/2
C0334245|T191|IS|59529006|SNOMEDCT_US|Epidermoid carcinoma in situ, NOS|8070/2
C0334245|T191|SY|59529006|SNOMEDCT_US|IEC - Intraepidermal carcinoma|8070/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Intraepidermal carcinoma|8070/2
C0334245|T191|IS|59529006|SNOMEDCT_US|Intraepidermal carcinoma, NOS|8070/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Intraepithelial squamous cell carcinoma|8070/2
C0334245|T191|PT|400066006|SNOMEDCT_US|Intraepithelial squamous cell carcinoma|8070/2
C0334245|T191|PT|252989001|SNOMEDCT_US|Squamous carcinoma in situ|8070/2
C0334245|T191|SY|252989001|SNOMEDCT_US|Squamous carcinoma in situ - category|8070/2
C0334245|T191|OF|189565007|SNOMEDCT_US|Squamous cell carcinoma in situ|8070/2
C0334245|T191|PT|189565007|SNOMEDCT_US|Squamous cell carcinoma in situ|8070/2
C0334245|T191|PT|59529006|SNOMEDCT_US|Squamous cell carcinoma in situ|8070/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Squamous cell carcinoma in situ, no ICD-O subtype|8070/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Squamous cell carcinoma in situ, no International Classification of Diseases for Oncology subtype|8070/2
C0334245|T191|IS|59529006|SNOMEDCT_US|Squamous cell carcinoma in situ, NOS|8070/2
C0334245|T191|SY|20365006|SNOMEDCT_US|Squamous intraepithelial neoplasia, grade III|8070/2
C0334245|T191|PT|20365006|SNOMEDCT_US|Squamous intraepithelial neoplasia, high grade|8070/2
C0007137|T191|DE|0000004527|AOD|squamous cell carcinoma|8070/3
C0007137|T191|PT|BI00611|BI|squamous cell carcinoma|8070/3
C0007137|T191|PT|1007881|CCPSS|SQUAMOUS CELL CARCINOMA|8070/3
C0007137|T191|SY|0000002437|CHV|epidermoid carcinoma|8070/3
C0007137|T191|SY|0000002437|CHV|squamous carcinoma|8070/3
C0007137|T191|SY|0000002437|CHV|squamous carcinomas|8070/3
C0007137|T191|PT|0000002437|CHV|squamous cell carcinoma|8070/3
C0007137|T191|SY|0000002437|CHV|squamous cell carcinomas|8070/3
C0007137|T191|SY|0000002437|CHV|squamous cell epithelioma|8070/3
C0007137|T191|ET|2000-3145|CSP|epidermoid carcinoma|8070/3
C0007137|T191|PT|2000-3145|CSP|squamous cell carcinoma|8070/3
C0007137|T191|GT|CARCINOMA SKIN|CST|CARCINOMA EPIDERMOID|8070/3
C0007137|T191|PT|HP:0002860|HPO|Squamous cell carcinoma|8070/3
C0007137|T191|PT|S77006|ICPC2P|Squamous cell carcinoma|8070/3
C0007137|T191|PTN|S77006|ICPC2P|squamous cell carcinoma|8070/3
C0007137|T191|PT|sh88005247|LCH_NW|Squamous cell carcinoma|8070/3
C0007137|T191|LA|LA23735-6|LNC|Squamous cell carcinoma|8070/3
C0007137|T191|LPN|LP17968-6|LNC|Squamous cell carcinoma|8070/3
C0007137|T191|LLT|10007349|MDR|Carcinoma epidermoid|8070/3
C0007137|T191|LLT|10007473|MDR|Carcinoma squamous|8070/3
C0007137|T191|LLT|10014987|MDR|Epidermoid carcinoma|8070/3
C0007137|T191|PT|10041823|MDR|Squamous cell carcinoma|8070/3
C0007137|T191|LLT|10041823|MDR|Squamous cell carcinoma|8070/3
C0007137|T191|PT|271412|MEDCIN|squamous cell carcinoma|8070/3
C0007137|T191|ET|D002294|MSH|Carcinoma, Epidermoid|8070/3
C0007137|T191|ET|D002294|MSH|Carcinoma, Planocellular|8070/3
C0007137|T191|ET|D002294|MSH|Carcinoma, Squamous|8070/3
C0007137|T191|MH|D002294|MSH|Carcinoma, Squamous Cell|8070/3
C0007137|T191|PM|D002294|MSH|Carcinomas, Epidermoid|8070/3
C0007137|T191|PM|D002294|MSH|Carcinomas, Planocellular|8070/3
C0007137|T191|PM|D002294|MSH|Carcinomas, Squamous|8070/3
C0007137|T191|PM|D002294|MSH|Carcinomas, Squamous Cell|8070/3
C0007137|T191|PM|D002294|MSH|Epidermoid Carcinoma|8070/3
C0007137|T191|PM|D002294|MSH|Epidermoid Carcinomas|8070/3
C0007137|T191|PM|D002294|MSH|Planocellular Carcinoma|8070/3
C0007137|T191|PM|D002294|MSH|Planocellular Carcinomas|8070/3
C0007137|T191|PM|D002294|MSH|Squamous Carcinoma|8070/3
C0007137|T191|PM|D002294|MSH|Squamous Carcinomas|8070/3
C0007137|T191|ET|D002294|MSH|Squamous Cell Carcinoma|8070/3
C0007137|T191|PM|D002294|MSH|Squamous Cell Carcinomas|8070/3
C0007137|T191|PN|NOCODE|MTH|Squamous cell carcinoma|8070/3
C0577691|T191|PT|C4829|NCI|Disseminated Squamous Cell Carcinoma|8070/3
C0007137|T191|SY|C2929|NCI|Epidermoid Carcinoma|8070/3
C0007137|T191|SY|C2929|NCI|Epidermoid Cell Cancer|8070/3
C0007137|T191|SY|C2929|NCI|Malignant Epidermoid Cell Neoplasm|8070/3
C0007137|T191|SY|C2929|NCI|Malignant Epidermoid Cell Tumor|8070/3
C0007137|T191|SY|C2929|NCI|Malignant Squamous Cell Neoplasm|8070/3
C0007137|T191|SY|C2929|NCI|Malignant Squamous Cell Tumor|8070/3
C0007137|T191|SY|C2929|NCI|Squamous Carcinoma|8070/3
C0007137|T191|SY|C2929|NCI|Squamous Cell Cancer|8070/3
C0007137|T191|PT|C2929|NCI|Squamous Cell Carcinoma|8070/3
C0007137|T191|SY|TCGA|NCI|Squamous Cell Carcinoma|8070/3
C0007137|T191|SY|C2929|NCI|Squamous Cell Carcinoma, NOS|8070/3
C0007137|T191|SY|C2929|NCI|Squamous Cell Carcinoma, Not Otherwise Specified|8070/3
C0007137|T191|SY|C2929|NCI|Squamous Cell Epithelioma|8070/3
C0007137|T191|PT|C2929|NCI_CDISC|CARCINOMA, SQUAMOUS CELL, MALIGNANT|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Epidermoid Carcinoma|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Epidermoid Cell Cancer|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Malignant Epidermoid Cell Neoplasm|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Malignant Epidermoid Cell Tumor|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Malignant Squamous Cell Neoplasm|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Malignant Squamous Cell Tumor|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Squamous Carcinoma|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Squamous Cell Cancer|8070/3
C0007137|T191|SY|C2929|NCI_CDISC|Squamous Cell Epithelioma|8070/3
C0007137|T191|PT|C2929|NCI_CPTAC|Squamous Cell Carcinoma|8070/3
C0007137|T191|PT|CDR0000046419|NCI_NCI-GLOSS|epidermoid carcinoma|8070/3
C0007137|T191|PT|CDR0000046595|NCI_NCI-GLOSS|squamous cell carcinoma|8070/3
C0577691|T191|AB|Xa7n8|RCD|Dissemin squam cell carcinoma|8070/3
C0577691|T191|PT|Xa7n8|RCD|Disseminated squamous cell carcinoma|8070/3
C0007137|T191|SY|Xa98E|RCD|Epidermoid carcinoma|8070/3
C0007137|T191|SY|Xa98E|RCD|SCC - Squamous cell carcinoma|8070/3
C0007137|T191|SY|Xa98E|RCD|Squamous carcinoma|8070/3
C0007137|T191|PT|Xa98E|RCD|Squamous cell carcinoma|8070/3
C0007137|T191|SY|Xa98E|RCD|Squamous cell epithelioma|8070/3
C0007137|T191|OP|BB2A.|RCDSY|Squamous cell carcinoma NOS|8070/3
C1275874|T191|SY|399739006|SNOMEDCT_US|Carcinosarcomatous squamous cell carcinoma|8070/3
C0577691|T191|PT|300987004|SNOMEDCT_US|Disseminated squamous cell carcinoma|8070/3
C0007137|T191|SY|28899001|SNOMEDCT_US|Epidermoid carcinoma|8070/3
C0007137|T191|IS|28899001|SNOMEDCT_US|Epidermoid carcinoma, NOS|8070/3
C5190966|T191|PT|783213006|SNOMEDCT_US|Human papillomavirus negative squamous cell carcinoma|8070/3
C5190967|T191|PT|783212001|SNOMEDCT_US|Human papillomavirus positive squamous cell carcinoma|8070/3
C1275874|T191|PT|399739006|SNOMEDCT_US|Metaplastic squamous cell carcinoma|8070/3
C0007137|T191|SY|28899001|SNOMEDCT_US|SCC - Squamous cell carcinoma|8070/3
C0007137|T191|SY|28899001|SNOMEDCT_US|Squamous carcinoma|8070/3
C0007137|T191|OAP|154605007|SNOMEDCT_US|Squamous cell carcinoma|8070/3
C0007137|T191|PT|28899001|SNOMEDCT_US|Squamous cell carcinoma|8070/3
C0007137|T191|OF|154605007|SNOMEDCT_US|Squamous cell carcinoma|8070/3
C0007137|T191|PT|402815007|SNOMEDCT_US|Squamous cell carcinoma|8070/3
C1302451|T191|PT|399494004|SNOMEDCT_US|Squamous cell carcinoma in post-traumatic skin lesion|8070/3
C0007137|T191|SY|28899001|SNOMEDCT_US|Squamous cell carcinoma, no ICD-O subtype|8070/3
C0007137|T191|SY|28899001|SNOMEDCT_US|Squamous cell carcinoma, no International Classification of Diseases for Oncology subtype|8070/3
C0007137|T191|IS|28899001|SNOMEDCT_US|Squamous cell carcinoma, NOS|8070/3
C0007137|T191|SY|28899001|SNOMEDCT_US|Squamous cell epithelioma|8070/3
C0007137|T191|PT|1798|WHO|CARCINOMA SQUAMOUS|8070/3
C0334246|T191|PT|0011888|CCPSS|SQUAMOUS CELL CARCINOMA METASTATIC|8070/6
C0334246|T191|PT|10063569|MDR|Metastatic squamous cell carcinoma|8070/6
C0334246|T191|LLT|10063569|MDR|Metastatic squamous cell carcinoma|8070/6
C0334246|T191|SY|351486|MEDCIN|squamous cell carcinoma metastatic|8070/6
C0334246|T191|PT|351486|MEDCIN|Squamous cell carcinoma, metastatic|8070/6
C0334246|T191|PT|C4104|NCI|Metastatic Squamous Cell Carcinoma|8070/6
C0334246|T191|AB|X77n0|RCD|Metastatic squamous cell ca|8070/6
C0334246|T191|PT|X77n0|RCD|Metastatic squamous cell carcinoma|8070/6
C0334246|T191|OA|BB2B.|RCDSY|Squamous cell ca.,metastat.|8070/6
C0334246|T191|OP|BB2B.|RCDSY|Squamous cell carcinoma, metastatic NOS|8070/6
C0334246|T191|PT|403906006|SNOMEDCT_US|Metastatic squamous cell carcinoma|8070/6
C0334246|T191|SY|64204000|SNOMEDCT_US|Metastatic squamous cell carcinoma|8070/6
C0334246|T191|PT|64204000|SNOMEDCT_US|Squamous cell carcinoma, metastatic|8070/6
C0334246|T191|IS|64204000|SNOMEDCT_US|Squamous cell carcinoma, metastatic, NOS|8070/6
C0022572|T191|PT|0000007053|CHV|keratoacanthoma|8071/1
C0022572|T191|SY|0000007053|CHV|keratoacanthomas|8071/1
C0022572|T191|PT|NOCODE|COSTAR|Keratoacanthoma|8071/1
C0022572|T191|PT|2020-2121|CSP|keratoacanthoma|8071/1
C0022572|T191|PT|HP:0031525|HPO|Keratoacanthoma|8071/1
C0022572|T191|PT|MTHU041235|ICPC2ICD10ENG|keratoacanthoma|8071/1
C0022572|T191|PT|S99026|ICPC2P|Keratoacanthoma|8071/1
C0022572|T191|PTN|S99026|ICPC2P|keratoacanthoma|8071/1
C0022572|T191|PT|U002570|LCH|Keratoacanthoma|8071/1
C0022572|T191|PT|sh85072036|LCH_NW|Keratoacanthoma|8071/1
C0022572|T191|LLT|10023347|MDR|Keratoacanthoma|8071/1
C0022572|T191|PT|10023347|MDR|Keratoacanthoma|8071/1
C0022572|T191|LLT|10073955|MDR|Squamous cell carcinoma, keratoacanthoma-type|8071/1
C0022572|T191|PT|272917|MEDCIN|keratoacanthoma|8071/1
C0022572|T191|MH|D007636|MSH|Keratoacanthoma|8071/1
C0022572|T191|PM|D007636|MSH|Keratoacanthomas|8071/1
C0022572|T191|PN|NOCODE|MTH|keratoacanthoma|8071/1
C0022572|T191|PT|C3146|NCI|Keratoacanthoma|8071/1
C0022572|T191|PT|CDR0000044253|NCI_NCI-GLOSS|keratoacanthoma|8071/1
C0022572|T191|SY|X78Rc|RCD|KA - Keratoacanthoma|8071/1
C0022572|T191|PT|X78Rc|RCD|Keratoacanthoma|8071/1
C0022572|T191|SY|X78Rc|RCD|Molluscum sebaceum|8071/1
C0022572|T191|SY|254662007|SNOMEDCT_US|KA - Keratoacanthoma|8071/1
C0022572|T191|OAS|156395005|SNOMEDCT_US|Keratoacanthoma|8071/1
C0022572|T191|OAS|267858008|SNOMEDCT_US|Keratoacanthoma|8071/1
C0022572|T191|PT|254662007|SNOMEDCT_US|Keratoacanthoma|8071/1
C0022572|T191|OF|201061007|SNOMEDCT_US|Keratoacanthoma|8071/1
C0022572|T191|OAP|201061007|SNOMEDCT_US|Keratoacanthoma|8071/1
C0022572|T191|OAP|58220003|SNOMEDCT_US|Keratoacanthoma|8071/1
C0022572|T191|OAS|201064004|SNOMEDCT_US|Keratoacanthoma|8071/1
C0022572|T191|IS|58220003|SNOMEDCT_US|Keratoacanthoma, NOS|8071/1
C0022572|T191|SY|254662007|SNOMEDCT_US|Molluscum sebaceum|8071/1
C0022572|T191|IT|0966|WHO|KERATOACANTHOMA|8071/1
C0334247|T191|PT|271413|MEDCIN|keratinizing squamous cell carcinoma|8071/3
C0334247|T191|PN|NOCODE|MTH|Squamous cell carcinoma, keratinizing|8071/3
C0334247|T191|PT|C4105|NCI|Keratinizing Squamous Cell Carcinoma|8071/3
C0334247|T191|SY|TCGA|NCI|Keratinizing Squamous Cell Carcinoma|8071/3
C0334247|T191|AB|Xa98F|RCD|Keratinising epidermoid ca|8071/3
C0334247|T191|SY|Xa98F|RCD|Keratinising epidermoid carcinoma|8071/3
C0334247|T191|AB|Xa98F|RCD|Keratinising SCC - large cell|8071/3
C0334247|T191|AB|Xa98F|RCD|Keratinising squamous cell ca|8071/3
C0334247|T191|PT|Xa98F|RCD|Keratinising squamous cell carcinoma|8071/3
C0334247|T191|SY|Xa98F|RCD|Keratinising squamous cell carcinoma - large cell|8071/3
C0334247|T191|AB|Xa98F|RCDAE|Keratinizing epidermoid ca|8071/3
C0334247|T191|SY|Xa98F|RCDAE|Keratinizing epidermoid carcinoma|8071/3
C0334247|T191|AB|Xa98F|RCDAE|Keratinizing SCC - large cell|8071/3
C0334247|T191|AB|Xa98F|RCDAE|Keratinizing squamous cell ca|8071/3
C0334247|T191|PT|Xa98F|RCDAE|Keratinizing squamous cell carcinoma|8071/3
C0334247|T191|SY|Xa98F|RCDAE|Keratinizing squamous cell carcinoma - large cell|8071/3
C0334247|T191|SY|Xa98F|RCDSA|Squamous cell carcinoma, keratinizing type NOS|8071/3
C0334247|T191|AB|Xa98F|RCDSY|Squamous cell ca keratinis|8071/3
C0334247|T191|SY|Xa98F|RCDSY|Squamous cell carcinoma, keratinising type NOS|8071/3
C0334247|T191|SYGB|18048008|SNOMEDCT_US|Epidermoid carcinoma, keratinising|8071/3
C0334247|T191|SY|18048008|SNOMEDCT_US|Epidermoid carcinoma, keratinizing|8071/3
C0334247|T191|SYGB|18048008|SNOMEDCT_US|Keratinising epidermoid carcinoma|8071/3
C0334247|T191|OAP|189568009|SNOMEDCT_US|Keratinising squamous cell carcinoma|8071/3
C0334247|T191|OF|189568009|SNOMEDCT_US|Keratinising squamous cell carcinoma|8071/3
C0334247|T191|SYGB|18048008|SNOMEDCT_US|Keratinising squamous cell carcinoma - large cell|8071/3
C0334247|T191|SY|18048008|SNOMEDCT_US|Keratinizing epidermoid carcinoma|8071/3
C0334247|T191|OAP|189568009|SNOMEDCT_US|Keratinizing squamous cell carcinoma|8071/3
C0334247|T191|SY|18048008|SNOMEDCT_US|Keratinizing squamous cell carcinoma - large cell|8071/3
C0334247|T191|PTGB|18048008|SNOMEDCT_US|Squamous cell carcinoma, keratinising|8071/3
C0334247|T191|PT|18048008|SNOMEDCT_US|Squamous cell carcinoma, keratinizing|8071/3
C0334247|T191|IS|18048008|SNOMEDCT_US|Squamous cell carcinoma, keratinizing, NOS|8071/3
C0334247|T191|SYGB|18048008|SNOMEDCT_US|Squamous cell carcinoma, large cell, keratinising|8071/3
C0334247|T191|SY|18048008|SNOMEDCT_US|Squamous cell carcinoma, large cell, keratinizing|8071/3
C0334248|T191|SY|271414|MEDCIN|large cell, nonkeratinizing squamous cell carcinoma|8072/3
C0334248|T191|PT|271414|MEDCIN|nonkeratinizing large cell squamous cell carcinoma|8072/3
C0334248|T191|PT|C65173|NCI|Non-Keratinizing Large Cell Squamous Cell Carcinoma|8072/3
C0334248|T191|SY|BB2D.|RCD|Non-keratinising epidermoid carcinoma - large cell|8072/3
C0334248|T191|AB|BB2D.|RCD|Non-keratinising SCC|8072/3
C0334248|T191|SY|BB2D.|RCD|Non-keratinising squamous cell carcinoma|8072/3
C0334248|T191|PT|BB2D.|RCD|Non-keratinising squamous cell carcinoma - large cell|8072/3
C0334248|T191|AB|BB2D.|RCD|Nonkerat epiderm ca-large cell|8072/3
C0334248|T191|AB|BB2D.|RCD|Nonkeratinising SCC-large cell|8072/3
C0334248|T191|SY|BB2D.|RCDAE|Non-keratinizing epidermoid carcinoma - large cell|8072/3
C0334248|T191|AB|BB2D.|RCDAE|Non-keratinizing SCC|8072/3
C0334248|T191|SY|BB2D.|RCDAE|Non-keratinizing squamous cell carcinoma|8072/3
C0334248|T191|PT|BB2D.|RCDAE|Non-keratinizing squamous cell carcinoma - large cell|8072/3
C0334248|T191|SYGB|45490001|SNOMEDCT_US|Epidermoid carcinoma, large cell, nonkeratinising|8072/3
C0334248|T191|SY|45490001|SNOMEDCT_US|Epidermoid carcinoma, large cell, nonkeratinizing|8072/3
C0334248|T191|SYGB|45490001|SNOMEDCT_US|Non-keratinising epidermoid carcinoma - large cell|8072/3
C0334248|T191|SYGB|45490001|SNOMEDCT_US|Non-keratinising squamous cell carcinoma|8072/3
C0334248|T191|SYGB|45490001|SNOMEDCT_US|Non-keratinising squamous cell carcinoma - large cell|8072/3
C0334248|T191|SY|45490001|SNOMEDCT_US|Non-keratinizing epidermoid carcinoma - large cell|8072/3
C0334248|T191|SY|45490001|SNOMEDCT_US|Non-keratinizing squamous cell carcinoma|8072/3
C0334248|T191|SY|45490001|SNOMEDCT_US|Non-keratinizing squamous cell carcinoma - large cell|8072/3
C0334248|T191|PTGB|45490001|SNOMEDCT_US|Squamous cell carcinoma, large cell, nonkeratinising|8072/3
C0334248|T191|PT|45490001|SNOMEDCT_US|Squamous cell carcinoma, large cell, nonkeratinizing|8072/3
C0334248|T191|SYGB|45490001|SNOMEDCT_US|Squamous cell carcinoma, nonkeratinising|8072/3
C1302524|T191|PTGB|399582005|SNOMEDCT_US|Squamous cell carcinoma, nonkeratinising, differentiated|8072/3
C1302619|T191|PTGB|399694008|SNOMEDCT_US|Squamous cell carcinoma, nonkeratinising, mixed differentiated and undifferentiated|8072/3
C0334248|T191|SY|45490001|SNOMEDCT_US|Squamous cell carcinoma, nonkeratinizing|8072/3
C1302524|T191|PT|399582005|SNOMEDCT_US|Squamous cell carcinoma, nonkeratinizing, differentiated|8072/3
C1302619|T191|PT|399694008|SNOMEDCT_US|Squamous cell carcinoma, nonkeratinizing, mixed differentiated and undifferentiated|8072/3
C0334248|T191|IS|45490001|SNOMEDCT_US|Squamous cell carcinoma, nonkeratinizing, NOS|8072/3
C3266067|T191|PT|449778005|SNOMEDCT_US|Undifferentiated nonkeratinizing squamous cell carcinoma|8072/3
C0334249|T191|PT|271415|MEDCIN|nonkeratinizing small cell squamous cell carcinoma|8073/3
C0334249|T191|SY|271415|MEDCIN|small cell, nonkeratinizing squamous cell carcinoma|8073/3
C0334249|T191|PT|C65175|NCI|Non-Keratinizing Small Cell Squamous Cell Carcinoma|8073/3
C0334249|T191|SY|BB2E.|RCD|Non-keratinising epidermoid carcinoma - small cell|8073/3
C0334249|T191|PT|BB2E.|RCD|Non-keratinising squamous cell carcinoma - small cell|8073/3
C0334249|T191|AB|BB2E.|RCD|Nonkerat epiderm ca-small cell|8073/3
C0334249|T191|AB|BB2E.|RCD|Nonkeratinising SCC-small cell|8073/3
C0334249|T191|SY|BB2E.|RCDAE|Non-keratinizing epidermoid carcinoma - small cell|8073/3
C0334249|T191|PT|BB2E.|RCDAE|Non-keratinizing squamous cell carcinoma - small cell|8073/3
C0334249|T191|SYGB|35718007|SNOMEDCT_US|Epidermoid carcinoma, small cell, nonkeratinising|8073/3
C0334249|T191|SY|35718007|SNOMEDCT_US|Epidermoid carcinoma, small cell, nonkeratinizing|8073/3
C0334249|T191|SYGB|35718007|SNOMEDCT_US|Non-keratinising epidermoid carcinoma - small cell|8073/3
C0334249|T191|SYGB|35718007|SNOMEDCT_US|Non-keratinising squamous cell carcinoma - small cell|8073/3
C0334249|T191|SY|35718007|SNOMEDCT_US|Non-keratinizing epidermoid carcinoma - small cell|8073/3
C0334249|T191|SY|35718007|SNOMEDCT_US|Non-keratinizing squamous cell carcinoma - small cell|8073/3
C0334249|T191|PTGB|35718007|SNOMEDCT_US|Squamous cell carcinoma, small cell, nonkeratinising|8073/3
C0334249|T191|PT|35718007|SNOMEDCT_US|Squamous cell carcinoma, small cell, nonkeratinizing|8073/3
C0349656|T191|LLT|10080970|MDR|Sarcomatoid squamous cell carcinoma|8074/3
C0349656|T191|SY|355121|MEDCIN|skin neoplasm carcinoma squamous spindle cell|8074/3
C0349656|T191|PT|355121|MEDCIN|Spindle cell squamous carcinoma of skin|8074/3
C0349656|T191|PT|271416|MEDCIN|spindle cell squamous cell carcinoma|8074/3
C0349656|T191|SY|C27084|NCI|Epidermoid Spindle Cell Carcinoma|8074/3
C0349656|T191|PT|C27084|NCI|Sarcomatoid Squamous Cell Carcinoma|8074/3
C0349656|T191|SY|C4666|NCI|Spindle Cell Squamous Carcinoma of Skin|8074/3
C0349656|T191|SY|C4666|NCI|Spindle Cell Squamous Carcinoma of the Skin|8074/3
C0349656|T191|SY|C27084|NCI|Squamous Cell Carcinoma, Sarcomatoid|8074/3
C0349656|T191|SY|C27084|NCI|Squamous Cell Carcinoma, Spindle Cell|8074/3
C0349656|T191|SY|C27084|NCI|Squamous Cell Spindle Cell Carcinoma|8074/3
C0349656|T191|AB|BB2F.|RCD|Epidermoid ca - spindle cell|8074/3
C0349656|T191|SY|BB2F.|RCD|Epidermoid carcinoma - spindle cell|8074/3
C0349656|T191|SY|X78RT|RCD|Pseudosarcoma of skin|8074/3
C0349656|T191|AB|BB2F.|RCD|SCC - spindle cell|8074/3
C0349656|T191|AB|X78RT|RCD|Spindle cell carcinoma of skin|8074/3
C0349656|T191|PT|X78RT|RCD|Spindle cell squamous carcinoma of skin|8074/3
C0349656|T191|PT|BB2F.|RCD|Squamous cell carcinoma - spindle cell|8074/3
C0349656|T191|SY|10288008|SNOMEDCT_US|Epidermoid carcinoma - spindle cell|8074/3
C0349656|T191|SY|10288008|SNOMEDCT_US|Epidermoid carcinoma, spindle cell|8074/3
C0349656|T191|SY|254653005|SNOMEDCT_US|Pseudosarcoma of skin|8074/3
C0349656|T191|SY|403900000|SNOMEDCT_US|Pseudosarcoma of the skin|8074/3
C0349656|T191|PT|254653005|SNOMEDCT_US|Spindle cell squamous carcinoma of skin|8074/3
C0349656|T191|PT|403900000|SNOMEDCT_US|Spindle cell squamous cell carcinoma|8074/3
C0349656|T191|SY|10288008|SNOMEDCT_US|Squamous cell carcinoma - spindle cell|8074/3
C0349656|T191|SY|10288008|SNOMEDCT_US|Squamous cell carcinoma, sarcomatoid|8074/3
C0349656|T191|PT|10288008|SNOMEDCT_US|Squamous cell carcinoma, spindle cell|8074/3
C0334250|T191|PT|355109|MEDCIN|Acantholytic squamous cell carcinoma|8075/3
C0334250|T191|PT|271417|MEDCIN|adenoid squamous cell carcinoma|8075/3
C0334250|T191|SY|355109|MEDCIN|malignant neoplasm carcinoma squamous cell acantholytic|8075/3
C0334250|T191|SY|C4106|NCI|Adenoid Squamous Carcinoma|8075/3
C0334250|T191|SY|C4106|NCI|Adenoid Squamous Cell Carcinoma|8075/3
C0334250|T191|SY|C4106|NCI|Pseudoglandular Epidermoid Carcinoma|8075/3
C0334250|T191|SY|C4106|NCI|Pseudoglandular Epidermoid Cell Carcinoma|8075/3
C0334250|T191|SY|C4106|NCI|Pseudoglandular Squamous Carcinoma|8075/3
C0334250|T191|PT|C4106|NCI|Pseudoglandular Squamous Cell Carcinoma|8075/3
C0334250|T191|AB|BB2G.|RCD|Adenoid squamous cell ca|8075/3
C0334250|T191|PT|BB2G.|RCD|Adenoid squamous cell carcinoma|8075/3
C0334250|T191|AB|BB2G.|RCD|Pseudoglandular SCC|8075/3
C0334250|T191|SY|BB2G.|RCD|Pseudoglandular squamous cell carcinoma|8075/3
C0334250|T191|PT|403901001|SNOMEDCT_US|Acantholytic squamous cell carcinoma|8075/3
C0334250|T191|SY|85956000|SNOMEDCT_US|Acantholytic squamous cell carcinoma|8075/3
C0334250|T191|PT|85956000|SNOMEDCT_US|Adenoid squamous cell carcinoma|8075/3
C0334250|T191|SY|85956000|SNOMEDCT_US|Pseudoglandular squamous cell carcinoma|8075/3
C4518234|T191|PT|733897002|SNOMEDCT_US|Pseudovascular squamous cell carcinoma|8075/3
C0334250|T191|SY|85956000|SNOMEDCT_US|Squamous cell carcinoma, acantholytic|8075/3
C0334251|T191|SY|271383|MEDCIN|carcinoma in situ squamous cell with questionable stromal invasion|8076/2
C0334251|T191|PT|271383|MEDCIN|squamous cell carcinoma in situ with questionable stromal invasion|8076/2
C0334251|T191|PT|C65176|NCI|Squamous Cell Carcinoma In Situ with Questionable Stromal Invasion|8076/2
C0334251|T191|AB|BB2H.|RCD|Epidermoid carcinoma in situ + questionable stromal invasion|8076/2
C0334251|T191|SY|BB2H.|RCD|Epidermoid carcinoma in situ with questionable stromal invasion|8076/2
C0334251|T191|AB|BB2H.|RCD|Epidermoid CIS+ ?stromal invas|8076/2
C0334251|T191|AB|BB2H.|RCD|SCC in situ+ ?stromal invasion|8076/2
C0334251|T191|AB|BB2H.|RCD|Squamous cell carcinoma in situ + ?stromal invasion|8076/2
C0334251|T191|PT|BB2H.|RCD|Squamous cell carcinoma in situ with questionable stromal invasion|8076/2
C0334251|T191|SY|5688000|SNOMEDCT_US|Epidermoid carcinoma in situ with questionable stromal invasion|8076/2
C0334251|T191|PT|5688000|SNOMEDCT_US|Squamous cell carcinoma in situ with questionable stromal invasion|8076/2
C0334252|T191|LLT|10073528|MDR|Microinvasive squamous cell carcinoma|8076/3
C0334252|T191|PT|271418|MEDCIN|microinvasive squamous cell carcinoma|8076/3
C0334252|T191|PT|C65178|NCI|Microinvasive Squamous Cell Carcinoma|8076/3
C0334252|T191|AB|BB2J.|RCD|Microinvasive squamous cell ca|8076/3
C0334252|T191|PT|BB2J.|RCD|Microinvasive squamous cell carcinoma|8076/3
C3164881|T191|SY|448406002|SNOMEDCT_US|CIN III with early stromal invasion|8076/3
C3164881|T191|PT|448406002|SNOMEDCT_US|Grade III squamous intraepithelial neoplasia with microinvasive squamous cell carcinoma|8076/3
C0334252|T191|SY|12478003|SNOMEDCT_US|Microinvasive squamous cell carcinoma|8076/3
C0334252|T191|PT|12478003|SNOMEDCT_US|Squamous cell carcinoma, microinvasive|8076/3
C0349458|T191|PT|BI00378|BI|cervical intra-epithelial neoplasm i|8077/0
C0349458|T191|AB|BI00378|BI|cin i|8077/0
C0349458|T191|PT|0059631|CCPSS|CERVICAL CANCER CIN I|8077/0
C0349458|T191|SY|0000031235|CHV|cin 1|8077/0
C0349458|T191|SY|0000031235|CHV|cin i|8077/0
C0349458|T191|SY|0000031235|CHV|mild cervical dysplasia|8077/0
C0349458|T191|PT|N87.0|ICD10|Mild cervical dysplasia|8077/0
C0349458|T191|PT|N87.0|ICD10CM|Mild cervical dysplasia|8077/0
C0349458|T191|AB|N87.0|ICD10CM|Mild cervical dysplasia|8077/0
C0349458|T191|AB|622.11|ICD9CM|Mild dysplasia of cervix|8077/0
C0349458|T191|PT|622.11|ICD9CM|Mild dysplasia of cervix|8077/0
C0349458|T191|PT|MTHU015897|ICPC2ICD10ENG|cervix; intraepithelial neoplasia, grade I|8077/0
C0349458|T191|PT|MTHU024459|ICPC2ICD10ENG|dysplasia; cervix, mild|8077/0
C0349458|T191|PT|MTHU052215|ICPC2ICD10ENG|neoplasia; intraepithelial, cervix, grade I|8077/0
C0349458|T191|PT|X86005|ICPC2P|CIN 1|8077/0
C0349458|T191|PTN|X86005|ICPC2P|CIN 1|8077/0
C0349458|T191|LLT|10049700|MDR|Cervical intraepithelial neoplasia I|8077/0
C1302773|T191|LLT|10064450|MDR|Low grade squamous intraepithelial lesion|8077/0
C1302773|T191|LLT|10064454|MDR|LSIL|8077/0
C0349458|T191|PT|275379|MEDCIN|mild cervical dysplasia|8077/0
C1302773|T191|PM|D000081483|MSH|Low Grade Squamous Intraepithelial Lesions|8077/0
C1302773|T191|PEP|D000081483|MSH|Low-Grade Squamous Intraepithelial Lesions|8077/0
C1302773|T191|PM|D000081483|MSH|LSIL, Low Grade Squamous Intraepithelial Lesions|8077/0
C1302773|T191|ET|D000081483|MSH|LSIL, Low-Grade Squamous Intraepithelial Lesions|8077/0
C0349458|T191|PN|NOCODE|MTH|Cervical intraepithelial neoplasia grade 1|8077/0
C1302773|T191|PN|NOCODE|MTH|Low Grade Squamous Intraepithelial Neoplasia|8077/0
C1334412|T191|AB|C27238|NCI|ASIN-L|8077/0
C1333458|T191|SY|C27427|NCI|Esophageal Low Grade Squamous Intraepithelial Neoplasia|8077/0
C1302773|T191|SY|C8335|NCI|Grade 1 Squamous Intraepithelial Neoplasia|8077/0
C1302798|T191|SY|C7351|NCI|Grade 2 Squamous Intraepithelial Lesion|8077/0
C1302798|T191|SY|C7351|NCI|Grade 2 Squamous Intraepithelial Neoplasia|8077/0
C1302773|T191|SY|C8335|NCI|Grade I Squamous Intraepithelial Neoplasia|8077/0
C1302798|T191|SY|C7351|NCI|Grade II Squamous Intraepithelial Lesion|8077/0
C1302798|T191|PT|C7351|NCI|Grade II Squamous Intraepithelial Neoplasia|8077/0
C1334412|T191|SY|C27238|NCI|Low Grade Anal Canal Intraepithelial Neoplasia|8077/0
C1334412|T191|SY|C27238|NCI|Low Grade Anal Canal Squamous Dysplasia|8077/0
C1334412|T191|PT|C27238|NCI|Low Grade Anal Canal Squamous Intraepithelial Neoplasia|8077/0
C1334412|T191|SY|C27238|NCI|Low Grade Anal Squamous Intraepithelial Neoplasia|8077/0
C0349458|T191|PT|C4630|NCI|Low Grade Cervical Intraepithelial Neoplasia|8077/0
C1333458|T191|SY|C27427|NCI|Low Grade Esophageal Squamous Dysplasia|8077/0
C1333458|T191|PT|C27427|NCI|Low Grade Esophageal Squamous Intraepithelial Neoplasia|8077/0
C1302773|T191|PT|C8335|NCI|Low Grade Squamous Intraepithelial Neoplasia|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Cervix Intraepithelial Neoplasia|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Cervix Uteri Intraepithelial Neoplasia|8077/0
C1334412|T191|SY|C27238|NCI|Low-Grade Intraepithelial Neoplasia of Anal Canal|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Intraepithelial Neoplasia of Cervix|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Intraepithelial Neoplasia of Cervix Uteri|8077/0
C1334412|T191|SY|C27238|NCI|Low-Grade Intraepithelial Neoplasia of the Anal Canal|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Intraepithelial Neoplasia of the Cervix|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Intraepithelial Neoplasia of the Cervix Uteri|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Intraepithelial Neoplasia of the Uterine Cervix|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Intraepithelial Neoplasia of Uterine Cervix|8077/0
C1302773|T191|SY|C8335|NCI|Low-Grade Squamous Intraepithelial Lesion|8077/0
C0349458|T191|SY|C4630|NCI|Low-Grade Uterine Cervix Intraepithelial Neoplasia|8077/0
C1302773|T191|AB|C8335|NCI|LSIL|8077/0
C1302773|T191|DN|C8335|NCI_CTRP|Low Grade Squamous Intraepithelial Neoplasia|8077/0
C1302773|T191|PT|CDR0000410514|NCI_NCI-GLOSS|low-grade squamous intraepithelial lesion|8077/0
C1302773|T191|PT|CDR0000410401|NCI_NCI-GLOSS|LSIL|8077/0
C0349458|T191|PT|CDR0000613645|PDQ|cervical intraepithelial neoplasia grade 1|8077/0
C0349458|T191|AB|CDR0000613645|PDQ|CIN1|8077/0
C1302773|T191|SY|CDR0000398204|PDQ|grade 1 squamous intraepithelial neoplasia|8077/0
C1302773|T191|SY|CDR0000398204|PDQ|grade I squamous intraepithelial neoplasia|8077/0
C1302773|T191|SY|CDR0000398204|PDQ|Low Grade Squamous Intraepithelial Neoplasia|8077/0
C1302773|T191|SY|CDR0000398204|PDQ|low-grade squamous intraepithelial lesion|8077/0
C1302773|T191|PT|CDR0000398204|PDQ|low-grade squamous intraepithelial neoplasia|8077/0
C1302773|T191|AB|CDR0000398204|PDQ|LSIL|8077/0
C0349458|T191|AB|Xa3HD|RCD|Cerv intraep neop grade I|8077/0
C0349458|T191|AB|Xa3HD|RCD|Cerv intraepith neoplasia 1|8077/0
C0349458|T191|PT|Xa3HD|RCD|Cervical intraepithelial neoplasia grade 1|8077/0
C0349458|T191|SY|Xa3HD|RCD|Cervical intraepithelial neoplasia grade I|8077/0
C0349458|T191|AB|Xa3HD|RCD|CIN I - Cerv intraep neopl 1|8077/0
C0349458|T191|SY|Xa3HD|RCD|CIN I - Cervical intraepithelial neoplasia 1|8077/0
C0349458|T191|SY|Xa3HD|RCD|Mild cervical dysplasia|8077/0
C0349458|T191|SY|Xa3HD|RCD|Mild dysplasia of cervix|8077/0
C0349458|T191|OAP|198342006|SNOMEDCT_US|Cervical intraepithelial neoplasia grade 1|8077/0
C0349458|T191|OF|198342006|SNOMEDCT_US|Cervical intraepithelial neoplasia grade 1|8077/0
C0349458|T191|PT|285836003|SNOMEDCT_US|Cervical intraepithelial neoplasia grade 1|8077/0
C0349458|T191|SY|285836003|SNOMEDCT_US|Cervical intraepithelial neoplasia grade I|8077/0
C0349458|T191|SY|285836003|SNOMEDCT_US|CIN I - Cervical intraepithelial neoplasia 1|8077/0
C1302773|T191|SY|112662005|SNOMEDCT_US|Low grade SIL|8077/0
C1302773|T191|PT|112662005|SNOMEDCT_US|Low-grade squamous intraepithelial lesion|8077/0
C1302773|T191|SY|112662005|SNOMEDCT_US|LSIL|8077/0
C0349458|T191|SY|285836003|SNOMEDCT_US|Mild cervical dysplasia|8077/0
C0349458|T191|SY|285836003|SNOMEDCT_US|Mild dysplasia of cervix|8077/0
C1302773|T191|PT|400002005|SNOMEDCT_US|Squamous intraepithelial neoplasia grade 1|8077/0
C1302798|T191|PT|400049009|SNOMEDCT_US|Squamous intraepithelial neoplasia grade 2|8077/0
C1302773|T191|SY|400002005|SNOMEDCT_US|Squamous intraepithelial neoplasia, grade I|8077/0
C1302798|T191|SY|400049009|SNOMEDCT_US|Squamous intraepithelial neoplasia, grade II|8077/0
C1302773|T191|PT|450595003|SNOMEDCT_US|Squamous intraepithelial neoplasia, low grade|8077/0
C0334245|T191|SY|0000029942|CHV|carcinoma squamous cell in situ|8077/2
C0333875|T191|SY|0000029841|CHV|high grade sil|8077/2
C0333875|T191|SY|0000029841|CHV|hsil|8077/2
C0334245|T191|SY|0000029942|CHV|in situ squamous cell carcinoma|8077/2
C0334245|T191|PT|0000029942|CHV|squamous cell carcinoma in situ|8077/2
C0333875|T191|LLT|10064451|MDR|High grade squamous intraepithelial lesion|8077/2
C0333875|T191|LLT|10064455|MDR|HSIL|8077/2
C0334245|T191|LLT|10022739|MDR|Intra-epidermal carcinoma|8077/2
C0334245|T191|LLT|10022782|MDR|Intraepidermal carcinoma|8077/2
C0334245|T191|PT|271382|MEDCIN|squamous cell carcinoma in situ|8077/2
C0333875|T191|PM|D000081483|MSH|High Grade Squamous Intraepithelial Lesions|8077/2
C0333875|T191|PEP|D000081483|MSH|High-Grade Squamous Intraepithelial Lesions|8077/2
C0333875|T191|PM|D000081483|MSH|HSIL, High Grade Squamous Intraepithelial Lesions|8077/2
C0333875|T191|ET|D000081483|MSH|HSIL, High-Grade Squamous Intraepithelial Lesions|8077/2
C0334245|T191|PN|NOCODE|MTH|Intraepithelial Squamous Cell Carcinoma|8077/2
C0334245|T191|SY|C27093|NCI|Epidermoid Carcinoma in situ|8077/2
C0334245|T191|SY|C27093|NCI|Epidermoid Cell Carcinoma in situ|8077/2
C1333451|T191|SY|C27426|NCI|Esophageal High-Grade Squamous Intraepithelial Neoplasia|8077/2
C0334245|T191|AB|C27093|NCI|Grade 3 SIN|8077/2
C0334245|T191|SY|C27093|NCI|Grade 3 Squamous Intraepithelial Neoplasia|8077/2
C0334245|T191|AB|C27093|NCI|Grade III SIN|8077/2
C0334245|T191|SY|C27093|NCI|Grade III Squamous Intraepithelial Neoplasia|8077/2
C1333451|T191|PT|C27426|NCI|High Grade Esophageal Squamous Intraepithelial Neoplasia|8077/2
C0333875|T191|PT|C8336|NCI|High Grade Squamous Intraepithelial Neoplasia|8077/2
C1333451|T191|SY|C27426|NCI|High-Grade Esophageal Squamous Dysplasia|8077/2
C1333451|T191|SY|C27426|NCI|High-Grade Esophageal Squamous Intraepithelial Neoplasia|8077/2
C0333875|T191|SY|C8336|NCI|High-Grade Squamous Intraepithelial Lesion|8077/2
C0333875|T191|AB|C8336|NCI|HSIL|8077/2
C0334245|T191|SY|C27093|NCI|Intraepithelial Squamous Cell Carcinoma|8077/2
C0334245|T191|SY|C27093|NCI|Squamous Carcinoma in situ|8077/2
C0334245|T191|SY|C27093|NCI|Squamous Cell Carcinoma in situ|8077/2
C0334245|T191|SY|C27093|NCI|Squamous Cell Carcinoma in-situ|8077/2
C0334245|T191|PT|C27093|NCI|Stage 0 Squamous Cell Carcinoma|8077/2
C0334245|T191|PT|C27093|NCI_CDISC|CARCINOMA, SQUAMOUS CELL, IN SITU, MALIGNANT|8077/2
C0334245|T191|SY|C27093|NCI_CDISC|Epidermoid Carcinoma In situ|8077/2
C0334245|T191|SY|C27093|NCI_CDISC|Epidermoid Cell Carcinoma In situ|8077/2
C0334245|T191|SY|C27093|NCI_CDISC|Grade 3 Squamous Intraepithelial Neoplasia|8077/2
C0334245|T191|SY|C27093|NCI_CDISC|Grade III Squamous Intraepithelial Neoplasia|8077/2
C0334245|T191|SY|C27093|NCI_CDISC|Intraepithelial Squamous Cell Carcinoma|8077/2
C0334245|T191|SY|C27093|NCI_CDISC|Squamous Carcinoma In situ|8077/2
C0334245|T191|SY|C27093|NCI_CDISC|Squamous Cell Carcinoma In situ|8077/2
C0333875|T191|DN|C8336|NCI_CTRP|High Grade Squamous Intraepithelial Neoplasia|8077/2
C0333875|T191|PT|CDR0000044762|NCI_NCI-GLOSS|high-grade squamous intraepithelial lesion|8077/2
C0333875|T191|PT|CDR0000409768|NCI_NCI-GLOSS|HSIL|8077/2
C0333875|T191|SY|CDR0000321379|PDQ|High Grade Squamous Intraepithelial Neoplasia|8077/2
C0333875|T191|PT|CDR0000321379|PDQ|high-grade squamous intraepithelial lesion|8077/2
C0333875|T191|SY|CDR0000321379|PDQ|high-grade squamous intraepithelial neoplasia|8077/2
C0333875|T191|SY|CDR0000321379|PDQ|HSIL|8077/2
C0334245|T191|SY|Xa98D|RCD|Epidermoid carcinoma in situ|8077/2
C0334245|T191|SY|Xa98D|RCD|IEC - Intraepidermal carcinoma|8077/2
C0334245|T191|SY|Xa98D|RCD|Intraepidermal carcinoma|8077/2
C0334245|T191|AB|Xa98D|RCD|Intraepithel squamous cell ca|8077/2
C0334245|T191|SY|Xa98D|RCD|Intraepithelial squamous cell carcinoma|8077/2
C0334245|T191|PT|X77n1|RCD|Squamous carcinoma in situ|8077/2
C0334245|T191|AB|Xa98D|RCD|Squamous cell ca in situ|8077/2
C0334245|T191|PT|Xa98D|RCD|Squamous cell carcinoma in situ|8077/2
C0334245|T191|AB|Xa98D|RCDSY|Squam cell ca-in-situ NOS|8077/2
C0334245|T191|SY|Xa98D|RCDSY|Squamous cell carcinoma in situ NOS|8077/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Epidermoid carcinoma in situ|8077/2
C0334245|T191|IS|59529006|SNOMEDCT_US|Epidermoid carcinoma in situ, NOS|8077/2
C0333875|T191|SY|22725004|SNOMEDCT_US|High grade SIL|8077/2
C0333875|T191|PT|22725004|SNOMEDCT_US|High-grade squamous intraepithelial lesion|8077/2
C0333875|T191|SY|22725004|SNOMEDCT_US|HSIL|8077/2
C0334245|T191|SY|59529006|SNOMEDCT_US|IEC - Intraepidermal carcinoma|8077/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Intraepidermal carcinoma|8077/2
C0334245|T191|IS|59529006|SNOMEDCT_US|Intraepidermal carcinoma, NOS|8077/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Intraepithelial squamous cell carcinoma|8077/2
C0334245|T191|PT|400066006|SNOMEDCT_US|Intraepithelial squamous cell carcinoma|8077/2
C0334245|T191|PT|252989001|SNOMEDCT_US|Squamous carcinoma in situ|8077/2
C0334245|T191|SY|252989001|SNOMEDCT_US|Squamous carcinoma in situ - category|8077/2
C0334245|T191|OF|189565007|SNOMEDCT_US|Squamous cell carcinoma in situ|8077/2
C0334245|T191|PT|189565007|SNOMEDCT_US|Squamous cell carcinoma in situ|8077/2
C0334245|T191|PT|59529006|SNOMEDCT_US|Squamous cell carcinoma in situ|8077/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Squamous cell carcinoma in situ, no ICD-O subtype|8077/2
C0334245|T191|SY|59529006|SNOMEDCT_US|Squamous cell carcinoma in situ, no International Classification of Diseases for Oncology subtype|8077/2
C0334245|T191|IS|59529006|SNOMEDCT_US|Squamous cell carcinoma in situ, NOS|8077/2
C0334245|T191|SY|20365006|SNOMEDCT_US|Squamous intraepithelial neoplasia, grade III|8077/2
C0334245|T191|PT|20365006|SNOMEDCT_US|Squamous intraepithelial neoplasia, high grade|8077/2
C1266004|T191|PT|271419|MEDCIN|squamous cell carcinoma with horn formation|8078/3
C1266004|T191|PT|C65179|NCI|Squamous Cell Carcinoma with Horn Formation|8078/3
C1266004|T191|PT|128633003|SNOMEDCT_US|Squamous cell carcinoma with horn formation|8078/3
C0154089|T191|PT|0000021388|CHV|erythroplasia of queyrat|8080/2
C0154089|T191|SY|0000021388|CHV|erythroplasia queyrat|8080/2
C0154089|T191|DI|U000595|DXP|ERYTHROPLASIA, QUEYRAT|8080/2
C0154089|T191|PX|D07.4|ICD10|Carcinoma in situ of penis|8080/2
C0154089|T191|PS|D07.4|ICD10|Penis|8080/2
C0154089|T191|PT|D07.4|ICD10CM|Carcinoma in situ of penis|8080/2
C0154089|T191|AB|D07.4|ICD10CM|Carcinoma in situ of penis|8080/2
C0154089|T191|ET|D07.4|ICD10CM|Erythroplasia of Queyrat NOS|8080/2
C0154089|T191|ET|D00-D09|ICD10CM|Queyrat's erythroplasia|8080/2
C0154089|T191|AB|233.5|ICD9CM|Ca in situ penis|8080/2
C0154089|T191|PT|233.5|ICD9CM|Carcinoma in situ of penis|8080/2
C0154089|T191|LLT|10007384|MDR|Carcinoma in situ of penis|8080/2
C0154089|T191|PT|10007384|MDR|Carcinoma in situ of penis|8080/2
C0154089|T191|LLT|10034328|MDR|Penis carcinoma in situ|8080/2
C0154089|T191|LLT|10037732|MDR|Queyrat erythroplasia|8080/2
C0154089|T191|PT|10037732|MDR|Queyrat erythroplasia|8080/2
C0154089|T191|PT|233440|MEDCIN|Bowen's disease of penis|8080/2
C0154089|T191|PT|97979|MEDCIN|carcinoma in situ of penis|8080/2
C0154089|T191|PT|355076|MEDCIN|Penile intraepithelial neoplasia grade III|8080/2
C0154089|T191|PT|233446|MEDCIN|Queyrat erythroplasia of glans penis|8080/2
C0154089|T191|PN|U000725|MTH|Carcinoma in situ of penis|8080/2
C0154089|T191|SY|C27790|NCI|Bowen Disease of the Penis|8080/2
C0154089|T191|SY|C27790|NCI|Bowen's Disease of Penis|8080/2
C0154089|T191|SY|C27790|NCI|Bowen's Disease of the Penis|8080/2
C0154089|T191|SY|C27790|NCI|Carcinoma in situ of Penis|8080/2
C0154089|T191|SY|C27790|NCI|Carcinoma in situ of the Penis|8080/2
C0154089|T191|SY|C27790|NCI|Erythroplasia of Queyrat|8080/2
C0154089|T191|SY|C27790|NCI|Grade III Penile Intraepithelial Neoplasia|8080/2
C0154089|T191|SY|C27790|NCI|Grade III Squamous Intraepithelial Lesion of Penis|8080/2
C0154089|T191|SY|C27790|NCI|Grade III Squamous Intraepithelial Lesion of the Penis|8080/2
C0154089|T191|PT|C27790|NCI|Penile Carcinoma In Situ|8080/2
C0154089|T191|SY|C27790|NCI|Penile Carcinoma In Situ AJCC v7|8080/2
C0154089|T191|SY|C27790|NCI|Queyrat Erythroplasia|8080/2
C0154089|T191|SY|C27790|NCI|Queyrat's Erythroplasia|8080/2
C0154089|T191|PT|CDR0000482355|NCI_NCI-GLOSS|stage 0 penile carcinoma in situ|8080/2
C0154089|T191|SY|X78il|RCD|Bowen's disease of glans penis|8080/2
C0154089|T191|SY|X78il|RCD|Bowen's disease of penis|8080/2
C0154089|T191|PT|B835.|RCD|Carcinoma in situ of penis|8080/2
C0154089|T191|AB|B835.|RCD|CIS - Carc in situ of penis|8080/2
C0154089|T191|SY|B835.|RCD|CIS - Carcinoma in situ of penis|8080/2
C0154089|T191|SY|X78il|RCD|Erythroplasia of Queyrat|8080/2
C0154089|T191|PT|X78il|RCD|Queyrat's erythroplasia|8080/2
C0154089|T191|OP|BB2K.|RCDSY|Queyrat's erythroplasia|8080/2
C0154089|T191|SY|398831006|SNOMEDCT_US|Bowen disease of penis|8080/2
C0154089|T191|OAS|255104003|SNOMEDCT_US|Bowen's disease of glans penis|8080/2
C0154089|T191|SY|398831006|SNOMEDCT_US|Bowen's disease of glans penis|8080/2
C0154089|T191|OAS|255104003|SNOMEDCT_US|Bowen's disease of penis|8080/2
C0154089|T191|PT|398831006|SNOMEDCT_US|Bowen's disease of penis|8080/2
C0154089|T191|SY|398831006|SNOMEDCT_US|Bowens disease of penis|8080/2
C0154089|T191|SY|92679008|SNOMEDCT_US|Cancer in situ of penis|8080/2
C0154089|T191|PT|92679008|SNOMEDCT_US|Carcinoma in situ of penis|8080/2
C0154089|T191|IS|92679008|SNOMEDCT_US|Carcinoma in situ of penis, NOS|8080/2
C0154089|T191|IS|92679008|SNOMEDCT_US|CIS - Carcinoma in situ of penis|8080/2
C0154089|T191|OAS|255104003|SNOMEDCT_US|Erythroplasia of Queyrat|8080/2
C0154089|T191|SY|398768004|SNOMEDCT_US|Erythroplasia of Queyrat|8080/2
C0154089|T191|PT|400092004|SNOMEDCT_US|Penile intraepithelial neoplasia grade III|8080/2
C0154089|T191|SY|398768004|SNOMEDCT_US|Queyrat erythroplasia|8080/2
C0154089|T191|SY|18348002|SNOMEDCT_US|Queyrat erythroplasia|8080/2
C0154089|T191|OF|255147003|SNOMEDCT_US|Queyrat's erythroplasia|8080/2
C0154089|T191|PT|398768004|SNOMEDCT_US|Queyrat's erythroplasia|8080/2
C0154089|T191|OAP|255104003|SNOMEDCT_US|Queyrat's erythroplasia|8080/2
C0154089|T191|PT|18348002|SNOMEDCT_US|Queyrat's erythroplasia|8080/2
C0154089|T191|OAP|255105002|SNOMEDCT_US|Queyrat's erythroplasia|8080/2
C0154089|T191|OAP|255147003|SNOMEDCT_US|Queyrat's erythroplasia|8080/2
C0154089|T191|OF|255105002|SNOMEDCT_US|Queyrat's erythroplasia|8080/2
C0154089|T191|OAS|189208007|SNOMEDCT_US|Queyrats's erythroplasia|8080/2
C0006079|T191|PT|0060852|CCPSS|BOWEN DISEASE|8081/2
C0006079|T191|SY|0000002117|CHV|bowen disease|8081/2
C0006079|T191|PT|0000002117|CHV|bowen's disease|8081/2
C0006079|T191|SY|0000002117|CHV|bowens disease|8081/2
C0006079|T191|SY|0000002117|CHV|disease bowen's|8081/2
C0006079|T191|PT|NOCODE|COSTAR|Bowen's Disease|8081/2
C0006079|T191|ET|D00-D09|ICD10CM|Bowen's disease|8081/2
C0006079|T191|PTN|S77001|ICPC2P|Bowens disease|8081/2
C0006079|T191|PT|S77001|ICPC2P|Disease;Bowens|8081/2
C0006079|T191|LLT|10006059|MDR|Bowen's disease|8081/2
C0006079|T191|PT|10006059|MDR|Bowen's disease|8081/2
C0006079|T191|PT|31503|MEDCIN|Bowen's disease|8081/2
C0006079|T191|DEV|D001913|MSH|BOWEN DIS|8081/2
C0006079|T191|ET|D001913|MSH|Bowen Disease|8081/2
C0006079|T191|MH|D001913|MSH|Bowen's Disease|8081/2
C0006079|T191|DEV|D001913|MSH|BOWENS DIS|8081/2
C0006079|T191|PM|D001913|MSH|Bowens Disease|8081/2
C0006079|T191|PM|D001913|MSH|Disease, Bowen|8081/2
C0006079|T191|PM|D001913|MSH|Disease, Bowen's|8081/2
C0006079|T191|PN|NOCODE|MTH|Bowen's Disease|8081/2
C0006079|T191|SY|C62571|NCI|Bowen Disease|8081/2
C0006079|T191|PT|C62571|NCI|Bowen Disease of the Skin|8081/2
C0006079|T191|SY|C62571|NCI|Bowen's Disease of the Skin|8081/2
C0006079|T191|SY|C62571|NCI|Intraepidermal Squamous Cell Carcinoma, Bowen Type|8081/2
C0006079|T191|DN|C62571|NCI_CTRP|Bowen Disease of the Skin|8081/2
C0006079|T191|PT|CDR0000044251|NCI_NCI-GLOSS|Bowen disease|8081/2
C0006079|T191|IS|X70Ld|RCD|BD - Bowen's disease|8081/2
C0006079|T191|IS|X70Ld|RCD|Bowen's disease|8081/2
C0006079|T191|OA|X70Ld|RCD|Intraepiderm SCC-Bowen's type|8081/2
C0006079|T191|OA|X70Ld|RCD|Intraepidermal SCC - Bowen's|8081/2
C0006079|T191|OP|X70Ld|RCD|Intraepidermal squamous cell carcinoma - Bowen's type|8081/2
C0006079|T191|IS|X70Ld|RCD|SCC - Intraepidermal squamous cell carcinoma - Bowen's type|8081/2
C0006079|T191|OP|BB2L.|RCDSY|Bowen's disease|8081/2
C0006079|T191|SY|84999002|SNOMEDCT_US|BD - Bowen's disease|8081/2
C0006079|T191|SY|84999002|SNOMEDCT_US|Bowen disease|8081/2
C0006079|T191|OAS|269582000|SNOMEDCT_US|Bowen's disease|8081/2
C0006079|T191|PT|84999002|SNOMEDCT_US|Bowen's disease|8081/2
C0006079|T191|OAS|154507009|SNOMEDCT_US|Bowen's disease|8081/2
C0006079|T191|OAS|189208007|SNOMEDCT_US|Bowen's disease|8081/2
C0006079|T191|SY|254656002|SNOMEDCT_US|Bowen's disease of skin|8081/2
C0006079|T191|OAP|240544007|SNOMEDCT_US|Intraepidermal squamous cell carcinoma - Bowen's type|8081/2
C0006079|T191|OF|240544007|SNOMEDCT_US|Intraepidermal squamous cell carcinoma - Bowen's type|8081/2
C0006079|T191|SY|84999002|SNOMEDCT_US|Intraepidermal squamous cell carcinoma, Bowen's type|8081/2
C0006079|T191|SY|84999002|SNOMEDCT_US|SCC - Intraepidermal squamous cell carcinoma - Bowen's type|8081/2
C0006079|T191|IT|1798|WHO|BOWEN'S DISEASE|8081/2
C0334254|T191|SY|0000029943|CHV|lymphoepithelial carcinoma|8082/3
C0334254|T191|PT|0000029943|CHV|lymphoepithelioma|8082/3
C0334254|T191|SY|0000029943|CHV|lymphoepithelioma-like carcinoma|8082/3
C0334254|T191|MTH_LLT|10082022|MDR|Lymphepithelioma|8082/3
C0334254|T191|LLT|10082023|MDR|Lymphoepithelial carcinoma|8082/3
C0334254|T191|LLT|10082022|MDR|Lymphoepithelioma|8082/3
C0334254|T191|PT|271420|MEDCIN|lymphoepithelial carcinoma|8082/3
C0334254|T191|PN|NOCODE|MTH|Lymphoepithelial carcinoma|8082/3
C0334254|T191|SY|C4107|NCI|Lymphoepithelial carcinoma|8082/3
C0334254|T191|SY|C4107|NCI|Lymphoepithelioma|8082/3
C0334254|T191|SY|C4107|NCI|Lymphoepithelioma-Like Carcinoma|8082/3
C0334254|T191|PT|C4107|NCI|Nasopharyngeal Type Undifferentiated Carcinoma|8082/3
C0334254|T191|SY|C4107|NCI|Schmincke Tumor|8082/3
C0334254|T191|PT|CDR0000044288|NCI_NCI-GLOSS|lymphoepithelioma|8082/3
C0334254|T191|PT|BB2M.|RCD|Lymphoepithelial carcinoma|8082/3
C0334254|T191|SY|BB2M.|RCD|Lymphoepithelioma|8082/3
C0334254|T191|SY|BB2M.|RCD|Schminke tumour|8082/3
C0334254|T191|SY|BB2M.|RCDAE|Lymphepithelioma|8082/3
C0334254|T191|SY|BB2M.|RCDAE|Schminke tumor|8082/3
C0334254|T191|PT|764938007|SNOMEDCT_US|Lymphoepithelial carcinoma|8082/3
C0334254|T191|PT|7300000|SNOMEDCT_US|Lymphoepithelial carcinoma|8082/3
C0334254|T191|SY|764938007|SNOMEDCT_US|Lymphoepithelial-like carcinoma|8082/3
C0334254|T191|SY|7300000|SNOMEDCT_US|Lymphoepithelioma|8082/3
C0334254|T191|SY|7300000|SNOMEDCT_US|Lymphoepithelioma-like carcinoma|8082/3
C0334254|T191|SY|7300000|SNOMEDCT_US|Schminke tumor|8082/3
C0334254|T191|SYGB|7300000|SNOMEDCT_US|Schminke tumour|8082/3
C1266005|T191|PT|271421|MEDCIN|basaloid squamous cell carcinoma|8083/3
C1266005|T191|SY|TCGA|NCI|Basaloid Squamous Cell Carcinoma|8083/3
C1266005|T191|PT|C54244|NCI|Basaloid Squamous Cell Carcinoma|8083/3
C1266005|T191|PT|128634009|SNOMEDCT_US|Basaloid squamous cell carcinoma|8083/3
C1266006|T191|PT|271422|MEDCIN|clear cell type squamous cell carcinoma|8084/3
C1266006|T191|SY|271422|MEDCIN|squamous cell carcinoma, clear cell type|8084/3
C1266006|T191|SY|TCGA|NCI|Squamous Cell Carcinoma, Clear Cell Type|8084/3
C1266006|T191|PT|C65180|NCI|Squamous Cell Carcinoma, Clear Cell Type|8084/3
C1266006|T191|PT|128635005|SNOMEDCT_US|Squamous cell carcinoma, clear cell type|8084/3
C0206710|T191|DEV|D018295|MSH|BASAL CELL NEOPL|8090/1
C0206710|T191|PM|D018295|MSH|Basal Cell Neoplasm|8090/1
C0206710|T191|ET|D018295|MSH|Basal Cell Neoplasms|8090/1
C0206710|T191|PM|D018295|MSH|Cell Neoplasm, Basal|8090/1
C0206710|T191|PM|D018295|MSH|Cell Neoplasms, Basal|8090/1
C0206710|T191|DEV|D018295|MSH|NEOPL BASAL CELL|8090/1
C0206710|T191|PM|D018295|MSH|Neoplasm, Basal Cell|8090/1
C0206710|T191|MH|D018295|MSH|Neoplasms, Basal Cell|8090/1
C0206710|T191|PN|NOCODE|MTH|Basal Cell Neoplasm|8090/1
C0206710|T191|PT|C3784|NCI|Basal Cell Neoplasm|8090/1
C0206710|T191|SY|C3784|NCI|Basal Cell Tumor|8090/1
C0206710|T191|PT|BB30.|RCD|Basal cell tumour|8090/1
C0206710|T191|PT|BB30.|RCDAE|Basal cell tumor|8090/1
C0206710|T191|OP|BB3z.|RCDSY|Basal cell neoplasm NOS|8090/1
C0206710|T191|OP|BB3..|RCDSY|Basal cell neoplasms|8090/1
C0206710|T191|SY|127570002|SNOMEDCT_US|Basal cell neoplasm|8090/1
C0206710|T191|PT|30649006|SNOMEDCT_US|Basal cell tumor|8090/1
C0206710|T191|SY|30649006|SNOMEDCT_US|Basal cell tumor, uncertain whether benign or malignant|8090/1
C0206710|T191|PTGB|30649006|SNOMEDCT_US|Basal cell tumour|8090/1
C4721806|T191|ET|0000004560|AOD|basal cell carcinoma|8090/3
C0007117|T191|PT|BI00572|BI|basal cell carcinoma|8090/3
C0007117|T191|AB|BI00572|BI|bcc|8090/3
C0007117|T191|PT|0033261|CCPSS|BASAL CELL CARCINOMA|8090/3
C4721806|T191|SD|NEO026|CCSR_10|Skin cancers - basal cell carcinoma|8090/3
C4721806|T191|PT|0000002425|CHV|basal cell carcinoma|8090/3
C4721806|T191|SY|0000002425|CHV|basal cell carcinoma of skin|8090/3
C4721806|T191|SY|0000002425|CHV|basal cell carcinoma of the skin|8090/3
C4721806|T191|SY|0000002425|CHV|basal cell carcinomas|8090/3
C4721806|T191|SY|0000002425|CHV|basal cell epithelioma|8090/3
C4721806|T191|SY|0000002425|CHV|basal cell skin cancer|8090/3
C4721806|T191|SY|0000002425|CHV|basalioma|8090/3
C4721806|T191|SY|0000002425|CHV|rodent ulcer|8090/3
C4721806|T191|PT|0000057894|CHV|rodent ulcer|8090/3
C4721806|T191|SY|0000002425|CHV|rodent ulcers|8090/3
C4721806|T191|PT|099|COSTAR|BASAL CELL CARCINOMA OF SKIN|8090/3
C4721806|T191|PT|100|COSTAR|BASAL CELL EPITHELIOMA|8090/3
C4721806|T191|PT|2000-2719|CSP|basal cell carcinoma|8090/3
C4721806|T191|GT|CARCINOMA SKIN|CST|BASAL CELL CARCINOMA|8090/3
C0007117|T191|DI|U000197|DXP|BASAL CELL CARCINOMA|8090/3
C4721806|T191|SY|NOCODE|DXP|EPITHELIOMA, BASAL CELL|8090/3
C4721806|T191|SY|NOCODE|DXP|SKIN CANCER, BASAL CELL CARCINOMA|8090/3
C4721806|T191|PT|HP:0002671|HPO|Basal cell carcinoma|8090/3
C4721806|T191|SY|HP:0002671|HPO|Basal cell carcinomas|8090/3
C4721806|T191|SY|HP:0002671|HPO|Basal cell epithelioma|8090/3
C4721806|T191|SY|HP:0002671|HPO|Basalioma|8090/3
C0007117|T191|PT|S77008|ICPC2P|Basal cell carcinoma|8090/3
C0007117|T191|PTN|S77008|ICPC2P|basal cell carcinoma|8090/3
C0007117|T191|PTN|S77007|ICPC2P|rodent ulcer|8090/3
C0007117|T191|PT|S77007|ICPC2P|Ulcer;rodent|8090/3
C0007117|T191|PT|U006152|LCH|Rodent ulcer|8090/3
C0007117|T191|PT|sh85114800|LCH_NW|Basal cell carcinoma|8090/3
C4721806|T191|LLT|10004146|MDR|Basal cell carcinoma|8090/3
C4721806|T191|PT|10004146|MDR|Basal cell carcinoma|8090/3
C4721806|T191|LLT|10004150|MDR|Basal cell epithelioma|8090/3
C4721806|T191|LLT|10077422|MDR|Basalioma|8090/3
C4721806|T191|LLT|10007286|MDR|Carcinoma basal cell|8090/3
C1304299|T191|LLT|10073090|MDR|Keratotic basal cell carcinoma|8090/3
C1368275|T191|LLT|10035029|MDR|Pigmented basal cell carcinoma|8090/3
C4721806|T191|LLT|10039208|MDR|Rodent ulcer|8090/3
C1304299|T191|PT|352406|MEDCIN|Basal cell carcinoma - keratotic|8090/3
C4721806|T191|PT|31723|MEDCIN|basal cell carcinoma of skin|8090/3
C0346016|T191|PT|355699|MEDCIN|Basal cell carcinoma with eccrine differentiation|8090/3
C1302747|T191|PT|352408|MEDCIN|Basal cell carcinoma with matrical differentiation|8090/3
C0334683|T191|PT|352411|MEDCIN|Basal cell carcinoma with sebaceous differentiation|8090/3
C4721806|T191|PT|356404|MEDCIN|Basal cell epithelioma|8090/3
C1304299|T191|SY|352406|MEDCIN|malignant neoplasm carcinoma basal cell keratotic|8090/3
C1302747|T191|SY|352408|MEDCIN|malignant neoplasm carcinoma basal cell with matrical differentiation|8090/3
C0334683|T191|SY|352411|MEDCIN|malignant neoplasm carcinoma basal cell with sebaceous differentiation|8090/3
C4721806|T191|SY|356404|MEDCIN|malignant neoplasm carcinoma epithelioma basal cell|8090/3
C1368275|T191|PT|355694|MEDCIN|Pigmented basal cell carcinoma|8090/3
C1368275|T191|SY|355694|MEDCIN|skin neoplasm malignant carcinoma basal cell pigmented|8090/3
C0346016|T191|SY|355699|MEDCIN|skin neoplasm malignant carcinoma basal cell with eccrine differentiation|8090/3
C0007117|T191|ET|405|MEDLINEPLUS|Basal Cell Carcinoma|8090/3
C4721806|T191|PM|D002280|MSH|Basal Cell Carcinoma|8090/3
C1304297|T191|CE|C537655|MSH|Basal cell carcinoma with follicular differentiation|8090/3
C1304297|T191|NM|C537655|MSH|Basal cell carcinoma, infundibulocystic|8090/3
C4721806|T191|PM|D002280|MSH|Basal Cell Carcinomas|8090/3
C4721806|T191|PM|D002280|MSH|Basal Cell Epithelioma|8090/3
C4721806|T191|PM|D002280|MSH|Basal Cell Epitheliomas|8090/3
C4721806|T191|MH|D002280|MSH|Carcinoma, Basal Cell|8090/3
C1368275|T191|PEP|D002280|MSH|Carcinoma, Basal Cell, Pigmented|8090/3
C4721806|T191|PM|D002280|MSH|Carcinomas, Basal Cell|8090/3
C4721806|T191|ET|D002280|MSH|Epithelioma, Basal Cell|8090/3
C4721806|T191|PM|D002280|MSH|Epitheliomas, Basal Cell|8090/3
C1304297|T191|CE|C537655|MSH|Infundibulocystic basal cell carcinoma|8090/3
C4721806|T191|ET|D002280|MSH|Rodent Ulcer|8090/3
C4721806|T191|PM|D002280|MSH|Rodent Ulcers|8090/3
C4721806|T191|ET|D002280|MSH|Ulcer, Rodent|8090/3
C4721806|T191|PM|D002280|MSH|Ulcers, Rodent|8090/3
C0007117|T191|PN|NOCODE|MTH|Basal cell carcinoma|8090/3
C4721806|T191|PT|100|MTH|BASAL CELL CARCINOMA OF SKIN|8090/3
C1368275|T191|PN|NOCODE|MTH|Pigmented Basal Cell Carcinoma|8090/3
C4721806|T191|PN|NOCODE|MTH|Skin Basal Cell Carcinoma|8090/3
C0334683|T191|PN|NOCODE|MTH|Skin Basal Cell Carcinoma with Sebaceous Differentiation|8090/3
C4721806|T191|SY|C2921|NCI|Basal Cell Cancer|8090/3
C4721806|T191|SY|C2921|NCI|Basal Cell Carcinoma|8090/3
C0007117|T191|PT|C156767|NCI|Basal Cell Carcinoma|8090/3
C4721806|T191|SY|C2921|NCI|Basal Cell Carcinoma of Skin|8090/3
C4721806|T191|SY|C2921|NCI|Basal Cell Carcinoma of the Skin|8090/3
C0334683|T191|SY|C4346|NCI|Basal Cell Carcinoma with Sebaceous Differentiation|8090/3
C4721806|T191|SY|C2921|NCI|Basal Cell Epithelioma|8090/3
C0334683|T191|SY|C4346|NCI|Basal Cell Epithelioma with Sebaceous Differentiation|8090/3
C4721806|T191|SY|C2921|NCI|Basal Cell Skin Carcinoma|8090/3
C0334683|T191|SY|C4346|NCI|Basosebaceous Epithelioma|8090/3
C4721806|T191|AB|C2921|NCI|BCC|8090/3
C1304297|T191|SY|C27540|NCI|Infundibulocystic Basal Cell Carcinoma|8090/3
C1304299|T191|SY|C54665|NCI|Keratotic Basal Cell Carcinoma|8090/3
C1368275|T191|SY|C9359|NCI|Pigmented Basal Cell Carcinoma|8090/3
C1304299|T191|SY|C54665|NCI|Pilar Basal Cell Carcinoma|8090/3
C0334683|T191|SY|C4346|NCI|Sebaceous Epithelioma|8090/3
C4721806|T191|PT|C2921|NCI|Skin Basal Cell Carcinoma|8090/3
C0334683|T191|PT|C4346|NCI|Skin Basal Cell Carcinoma with Sebaceous Differentiation|8090/3
C1304297|T191|PT|C27540|NCI|Skin Infundibulocystic Basal Cell Carcinoma|8090/3
C1304299|T191|PT|C54665|NCI|Skin Keratotic Basal Cell Carcinoma|8090/3
C1368275|T191|PT|C9359|NCI|Skin Pigmented Basal Cell Carcinoma|8090/3
C0007117|T191|PT|C156767|NCI_CPTAC|Basal Cell Carcinoma|8090/3
C4721806|T191|PT|C2921|NCI_CPTAC|Skin Basal Cell Carcinoma|8090/3
C4721806|T191|PT|10004146|NCI_CTEP-SDC|Basal cell carcinoma|8090/3
C0007117|T191|DN|C156767|NCI_CTRP|Basal Cell Carcinoma|8090/3
C4721806|T191|DN|C2921|NCI_CTRP|Skin Basal Cell Cancer|8090/3
C4721806|T191|PT|CDR0000667109|NCI_NCI-GLOSS|basal cell cancer|8090/3
C4721806|T191|PT|CDR0000046515|NCI_NCI-GLOSS|basal cell carcinoma|8090/3
C4721806|T191|ET|CDR0000039109|PDQ|basal cell carcinoma of the skin|8090/3
C4721806|T191|PSC|CDR0000039109|PDQ|basal cell carcinoma of the skin|8090/3
C4721806|T191|SY|CDR0000039109|PDQ|carcinoma of the skin, basal cell|8090/3
C4721806|T191|SY|CDR0000039109|PDQ|carcinoma, basal cell, skin|8090/3
C0007117|T191|PT|Xa98G|RCD|Basal cell carcinoma|8090/3
C4721806|T191|PT|X78SS|RCD|Basal cell carcinoma of skin|8090/3
C0346016|T191|PT|X78Sg|RCD|Basal cell carcinoma with eccrine differentiation|8090/3
C4721806|T191|SY|X78SS|RCD|Basalioma|8090/3
C4721806|T191|AB|X78SS|RCD|BCC - Basal cell carc of skin|8090/3
C0007117|T191|SY|Xa98G|RCD|BCC - Basal cell carcinoma|8090/3
C4721806|T191|SY|X78SS|RCD|BCC - Basal cell carcinoma of skin|8090/3
C0346016|T191|AB|X78Sg|RCD|BCC with eccrine differentn|8090/3
C4721806|T191|OP|XM1ML|RCD|Epithelioma basal cell|8090/3
C1368275|T191|SY|Xa98G|RCD|Pigmented basal cell carcinoma|8090/3
C4721806|T191|SY|X78SS|RCD|Rodent ulcer|8090/3
C4721806|T191|SY|X78SS|RCD|RU - Rodent ulcer|8090/3
C0007117|T191|OP|BB31.|RCDSY|Basal cell carcinoma NOS|8090/3
C0007117|T191|PT|1338007|SNOMEDCT_US|Basal cell carcinoma|8090/3
C0007117|T191|OAS|154507009|SNOMEDCT_US|Basal cell carcinoma|8090/3
C0007117|T191|OAS|188083002|SNOMEDCT_US|Basal cell carcinoma|8090/3
C4721806|T191|OAS|269582000|SNOMEDCT_US|Basal cell carcinoma|8090/3
C1304299|T191|PT|402528005|SNOMEDCT_US|Basal cell carcinoma - keratotic|8090/3
C4721806|T191|PT|254701007|SNOMEDCT_US|Basal cell carcinoma of skin|8090/3
C1302446|T191|PT|399487002|SNOMEDCT_US|Basal cell carcinoma with adnexal differentiation|8090/3
C0346016|T191|PT|399470004|SNOMEDCT_US|Basal cell carcinoma with eccrine differentiation|8090/3
C0346016|T191|PT|254710004|SNOMEDCT_US|Basal cell carcinoma with eccrine differentiation|8090/3
C1304297|T191|PT|399746002|SNOMEDCT_US|Basal cell carcinoma with follicular differentiation|8090/3
C1302747|T191|PT|402530007|SNOMEDCT_US|Basal cell carcinoma with matrical differentiation|8090/3
C1302747|T191|PT|399958006|SNOMEDCT_US|Basal cell carcinoma with matrical differentiation|8090/3
C0334683|T191|PT|402533009|SNOMEDCT_US|Basal cell carcinoma with sebaceous differentiation|8090/3
C0334683|T191|PT|400087001|SNOMEDCT_US|Basal cell carcinoma with sebaceous differentiation|8090/3
C0007117|T191|IS|1338007|SNOMEDCT_US|Basal cell carcinoma, NOS|8090/3
C4721806|T191|SY|1338007|SNOMEDCT_US|Basal cell epithelioma|8090/3
C4721806|T191|SY|254701007|SNOMEDCT_US|Basalioma|8090/3
C0007117|T191|SY|1338007|SNOMEDCT_US|Basiloma|8090/3
C0007117|T191|SY|1338007|SNOMEDCT_US|BCC - Basal cell carcinoma|8090/3
C4721806|T191|SY|254701007|SNOMEDCT_US|BCC - Basal cell carcinoma of skin|8090/3
C4721806|T191|SY|254701007|SNOMEDCT_US|Cancer of skin, basal cell|8090/3
C0346016|T191|SY|399470004|SNOMEDCT_US|Eccrine basal cell carcinoma|8090/3
C4721806|T191|OAS|188083002|SNOMEDCT_US|Epithelioma basal cell|8090/3
C4721806|T191|PT|275265005|SNOMEDCT_US|Epithelioma basal cell|8090/3
C1304297|T191|SY|399746002|SNOMEDCT_US|Infundibulocystic basal cell carcinoma|8090/3
C1304299|T191|PT|399547009|SNOMEDCT_US|Keratotic basal cell carcinoma|8090/3
C1368275|T191|SY|1338007|SNOMEDCT_US|Pigmented basal cell carcinoma|8090/3
C1368275|T191|PT|403909004|SNOMEDCT_US|Pigmented basal cell carcinoma|8090/3
C1368275|T191|PT|399585007|SNOMEDCT_US|Pigmented basal cell carcinoma|8090/3
C4721806|T191|SY|254701007|SNOMEDCT_US|Rodent ulcer|8090/3
C4721806|T191|OAS|269582000|SNOMEDCT_US|Rodent ulcer|8090/3
C0007117|T191|IS|399049001|SNOMEDCT_US|Rodent ulcer|8090/3
C0007117|T191|OAS|188083002|SNOMEDCT_US|Rodent ulcer|8090/3
C0007117|T191|OAS|154507009|SNOMEDCT_US|Rodent ulcer|8090/3
C0007117|T191|SY|1338007|SNOMEDCT_US|Rodent ulcer|8090/3
C4721806|T191|SY|254701007|SNOMEDCT_US|RU - Rodent ulcer|8090/3
C4721806|T191|PT|1240|WHO|BASAL CELL CARCINOMA|8090/3
C4721806|T191|IT|1240|WHO|CARCINOMA BASAL CELL|8090/3
C0334256|T191|SY|C4108|NCI|Multicentric Basal Cell Carcinoma|8091/3
C0334256|T191|PT|C4108|NCI|Superficial Multifocal Basal Cell Carcinoma|8091/3
C0334256|T191|AB|BB32.|RCD|Multicentric basal cell ca|8091/3
C0334256|T191|PT|BB32.|RCD|Multicentric basal cell carcinoma|8091/3
C0334256|T191|SY|61098004|SNOMEDCT_US|Multicentric basal cell carcinoma|8091/3
C0334256|T191|PT|61098004|SNOMEDCT_US|Multifocal superficial basal cell carcinoma|8091/3
C0555191|T191|LLT|10027981|MDR|Morpheaform basal cell carcinoma|8092/3
C0555191|T191|LLT|10062787|MDR|Morphoeaform basal cell carcinoma|8092/3
C0555191|T191|SY|355700|MEDCIN|malignant neoplasm carcinoma basal cell morpheic|8092/3
C0555191|T191|PT|355700|MEDCIN|Morpheic basal cell carcinoma|8092/3
C0334257|T191|PN|NOCODE|MTH|Infiltrating basal cell carcinoma|8092/3
C0555191|T191|PN|NOCODE|MTH|Morpheic basal cell carcinoma|8092/3
C0555191|T191|SY|C27182|NCI|Basal Cell Carcinoma Sclerosing Type|8092/3
C0334257|T191|SY|C27539|NCI|Infiltrating Basal Cell Carcinoma|8092/3
C0555191|T191|SY|C27182|NCI|Morphea-Type Basal Cell Carcinoma|8092/3
C0555191|T191|SY|C27182|NCI|Morpheaform Basal Cell Carcinoma|8092/3
C0555191|T191|SY|C27182|NCI|Sclerosing Type Basal Cell Carcinoma|8092/3
C0334257|T191|PT|C27539|NCI|Skin Infiltrating Basal Cell Carcinoma|8092/3
C0555191|T191|AB|Xa98H|RCD|Basal cell ca, sclerosing type|8092/3
C0555191|T191|OA|BB33.|RCD|Basal cell carcinoma - morphoe|8092/3
C0555191|T191|OP|BB33.|RCD|Basal cell carcinoma - morphoeic|8092/3
C0555191|T191|PT|Xa98H|RCD|Basal cell carcinoma - sclerosing type|8092/3
C0555191|T191|PT|134152008|SNOMEDCT_US|Basal cell carcinoma - morpheic|8092/3
C0555191|T191|PTGB|134152008|SNOMEDCT_US|Basal cell carcinoma - morphoeic|8092/3
C0555191|T191|PT|302821007|SNOMEDCT_US|Basal cell carcinoma - sclerosing type|8092/3
C5230950|T191|PT|816972004|SNOMEDCT_US|Basal cell carcinoma with sarcomatoid differentiation|8092/3
C0334257|T191|SY|56665009|SNOMEDCT_US|Basal cell carcinoma, desmoplastic type|8092/3
C0555191|T191|IS|56665009|SNOMEDCT_US|Basal cell carcinoma, morphea|8092/3
C0555191|T191|SY|56665009|SNOMEDCT_US|Basal cell carcinoma, morpheic|8092/3
C0555191|T191|SY|302821007|SNOMEDCT_US|Basal cell carcinoma, sclerosing type|8092/3
C0555191|T191|SY|403913006|SNOMEDCT_US|Cicatrising basal cell carcinoma|8092/3
C0334257|T191|PT|56665009|SNOMEDCT_US|Infiltrating basal cell carcinoma|8092/3
C0334257|T191|SY|56665009|SNOMEDCT_US|Infiltrating basal cell carcinoma, non-sclerosing|8092/3
C0334257|T191|SY|56665009|SNOMEDCT_US|Infiltrating basal cell carcinoma, sclerosing|8092/3
C0555191|T191|SY|134152008|SNOMEDCT_US|Morpheaform basal cell carcinoma|8092/3
C0555191|T191|PT|403913006|SNOMEDCT_US|Morpheic basal cell carcinoma|8092/3
C0346013|T191|PT|0000031041|CHV|fibroepithelioma|8093/3
C0346013|T191|SY|0000031041|CHV|fibroepithelioma of pinkus|8093/3
C0346013|T191|SY|0000031041|CHV|fibroepithelioma pinkus|8093/3
C0346013|T191|SY|0000031041|CHV|pinkus tumor|8093/3
C0346013|T191|SY|0000031041|CHV|pinkus tumour|8093/3
C0346013|T191|LLT|10073089|MDR|Fibroepithelial basal cell carcinoma|8093/3
C0346013|T191|LLT|10016625|MDR|Fibroepithelioma of pinkus|8093/3
C0346013|T191|PT|356501|MEDCIN|Fibroepithelioma of Pinkus|8093/3
C0346013|T191|SY|356501|MEDCIN|skin neoplasm malignant carcinoma basal cell fibroepithelioma of pinkus|8093/3
C0346013|T191|SY|C4109|NCI|Fibroepithelial Basal Cell Carcinoma|8093/3
C0346013|T191|SY|C4109|NCI|Fibroepithelioma of Pinkus|8093/3
C0346013|T191|SY|C4109|NCI|Pinkus Tumor|8093/3
C0346013|T191|PT|C4109|NCI|Skin Fibroepithelial Basal Cell Carcinoma|8093/3
C0346013|T191|AB|BB34.|RCD|Fibroepithelial basal cell ca|8093/3
C0346013|T191|PT|BB34.|RCD|Fibroepithelial basal cell carcinoma|8093/3
C0346013|T191|PT|X78SU|RCD|Fibroepithelioma of Pinkus|8093/3
C0346013|T191|SY|X78SU|RCD|Pinkus tumour|8093/3
C0346013|T191|SY|X78SU|RCDAE|Pinkus tumor|8093/3
C0346013|T191|PT|43369006|SNOMEDCT_US|Basal cell carcinoma, fibroepithelial|8093/3
C0346013|T191|SY|43369006|SNOMEDCT_US|Fibroepithelial basal cell carcinoma|8093/3
C0346013|T191|SY|43369006|SNOMEDCT_US|Fibroepithelial basal cell carcinoma, Pinkus type|8093/3
C0346013|T191|SY|43369006|SNOMEDCT_US|Fibroepithelioma|8093/3
C0346013|T191|PT|254703005|SNOMEDCT_US|Fibroepithelioma of Pinkus|8093/3
C0346013|T191|SY|43369006|SNOMEDCT_US|Fibroepithelioma of Pinkus type|8093/3
C0346013|T191|SY|43369006|SNOMEDCT_US|Pinkus tumor|8093/3
C0346013|T191|SY|254703005|SNOMEDCT_US|Pinkus tumor|8093/3
C0346013|T191|SYGB|254703005|SNOMEDCT_US|Pinkus tumour|8093/3
C0346013|T191|SYGB|43369006|SNOMEDCT_US|Pinkus tumour|8093/3
C0007118|T191|SY|0000002426|CHV|basosquamous carcinoma|8094/3
C0007118|T191|PT|0000002426|CHV|basosquamous cell carcinoma|8094/3
C0007118|T191|PT|2000-2932|CSP|basosquamous cell carcinoma|8094/3
C0007118|T191|GT|CARCINOMA SKIN|CST|CARCINOMA BASOSQUAMOUS|8094/3
C0007118|T191|LLT|10004154|MDR|Basal squamous cell carcinoma|8094/3
C0007118|T191|LLT|10004162|MDR|Basi squamous cell carcinoma|8094/3
C0007118|T191|LLT|10004178|MDR|Basosquamous carcinoma|8094/3
C0007118|T191|PT|10004178|MDR|Basosquamous carcinoma|8094/3
C0007118|T191|LLT|10004179|MDR|Basosquamous carcinoma of skin|8094/3
C0007118|T191|PT|10004179|MDR|Basosquamous carcinoma of skin|8094/3
C0007118|T191|LLT|10007287|MDR|Carcinoma basosquamous|8094/3
C0007118|T191|LLT|10007288|MDR|Carcinoma basosquamous of skin|8094/3
C0007118|T191|LLT|10027492|MDR|Metatypical basal cell carcinoma|8094/3
C0007118|T191|PT|313918|MEDCIN|basosquamous carcinoma of skin|8094/3
C0007118|T191|SY|313918|MEDCIN|skin neoplasm malignant carcinoma basosquamous|8094/3
C0007118|T191|PM|D002281|MSH|Basosquamous Carcinoma|8094/3
C0007118|T191|PM|D002281|MSH|Basosquamous Carcinomas|8094/3
C0007118|T191|MH|D002281|MSH|Carcinoma, Basosquamous|8094/3
C0007118|T191|PM|D002281|MSH|Carcinomas, Basosquamous|8094/3
C0007118|T191|SY|C2922|NCI|Basosquamous Carcinoma|8094/3
C0007118|T191|SY|C2922|NCI|Basosquamous Cell Carcinoma|8094/3
C0007118|T191|PT|C2922|NCI|Skin Basosquamous Cell Carcinoma|8094/3
C0007118|T191|SY|C2922|NCI|Skin Mixed Basal and Squamous Cell Carcinoma|8094/3
C0007118|T191|SY|C2922|NCI_CDISC|Basosquamous Carcinoma|8094/3
C0007118|T191|SY|C2922|NCI_CDISC|Basosquamous Cell Carcinoma|8094/3
C0007118|T191|PT|C2922|NCI_CDISC|BASOSQUAMOUS TUMOR, MALIGNANT|8094/3
C0007118|T191|SY|C2922|NCI_CDISC|Skin Mixed Basal and Squamous Cell Carcinoma|8094/3
C0007118|T191|PT|BB35.|RCD|Basosquamous carcinoma|8094/3
C0007118|T191|PT|X78ST|RCD|Basosquamous carcinoma of skin|8094/3
C0007118|T191|SY|X78ST|RCD|BCC - Metatypical basal cell carcinoma of skin|8094/3
C0007118|T191|SY|X78ST|RCD|Metatypical basal cell carcinoma of skin|8094/3
C0007118|T191|AB|X78ST|RCD|Metatypical BCC of skin|8094/3
C0007118|T191|PT|BB36.|RCD|Metatypical carcinoma|8094/3
C0007118|T191|AB|BB35.|RCD|Mixed basal - squamous cell ca|8094/3
C0007118|T191|SY|BB35.|RCD|Mixed basal - squamous cell carcinoma|8094/3
C0007118|T191|SY|37304002|SNOMEDCT_US|Basisquamous cell carcinoma|8094/3
C0007118|T191|PT|37304002|SNOMEDCT_US|Basosquamous carcinoma|8094/3
C0007118|T191|PT|254702000|SNOMEDCT_US|Basosquamous carcinoma of skin|8094/3
C0007118|T191|SY|254702000|SNOMEDCT_US|BCC - Metatypical basal cell carcinoma of skin|8094/3
C0007118|T191|SY|254702000|SNOMEDCT_US|Metatypical basal cell carcinoma of skin|8094/3
C0007118|T191|PT|6641007|SNOMEDCT_US|Metatypical carcinoma|8094/3
C0007118|T191|SY|37304002|SNOMEDCT_US|Mixed basal - squamous cell carcinoma|8094/3
C0007118|T191|SY|37304002|SNOMEDCT_US|Mixed basal-squamous cell carcinoma|8094/3
C0007118|T191|SY|0000002426|CHV|basosquamous carcinoma|8095/3
C0007118|T191|PT|0000002426|CHV|basosquamous cell carcinoma|8095/3
C0007118|T191|PT|2000-2932|CSP|basosquamous cell carcinoma|8095/3
C0007118|T191|GT|CARCINOMA SKIN|CST|CARCINOMA BASOSQUAMOUS|8095/3
C0007118|T191|LLT|10004154|MDR|Basal squamous cell carcinoma|8095/3
C0007118|T191|LLT|10004162|MDR|Basi squamous cell carcinoma|8095/3
C0007118|T191|LLT|10004178|MDR|Basosquamous carcinoma|8095/3
C0007118|T191|PT|10004178|MDR|Basosquamous carcinoma|8095/3
C0007118|T191|LLT|10004179|MDR|Basosquamous carcinoma of skin|8095/3
C0007118|T191|PT|10004179|MDR|Basosquamous carcinoma of skin|8095/3
C0007118|T191|LLT|10007287|MDR|Carcinoma basosquamous|8095/3
C0007118|T191|LLT|10007288|MDR|Carcinoma basosquamous of skin|8095/3
C0007118|T191|LLT|10027492|MDR|Metatypical basal cell carcinoma|8095/3
C0007118|T191|PT|313918|MEDCIN|basosquamous carcinoma of skin|8095/3
C0007118|T191|SY|313918|MEDCIN|skin neoplasm malignant carcinoma basosquamous|8095/3
C0007118|T191|PM|D002281|MSH|Basosquamous Carcinoma|8095/3
C0007118|T191|PM|D002281|MSH|Basosquamous Carcinomas|8095/3
C0007118|T191|MH|D002281|MSH|Carcinoma, Basosquamous|8095/3
C0007118|T191|PM|D002281|MSH|Carcinomas, Basosquamous|8095/3
C0007118|T191|SY|C2922|NCI|Basosquamous Carcinoma|8095/3
C0007118|T191|SY|C2922|NCI|Basosquamous Cell Carcinoma|8095/3
C0007118|T191|PT|C2922|NCI|Skin Basosquamous Cell Carcinoma|8095/3
C1883040|T191|SY|C66903|NCI|Skin Metatypical Basal Cell Carcinoma|8095/3
C1883040|T191|PT|C66903|NCI|Skin Metatypical Carcinoma|8095/3
C0007118|T191|SY|C2922|NCI|Skin Mixed Basal and Squamous Cell Carcinoma|8095/3
C0007118|T191|SY|C2922|NCI_CDISC|Basosquamous Carcinoma|8095/3
C0007118|T191|SY|C2922|NCI_CDISC|Basosquamous Cell Carcinoma|8095/3
C0007118|T191|PT|C2922|NCI_CDISC|BASOSQUAMOUS TUMOR, MALIGNANT|8095/3
C0007118|T191|SY|C2922|NCI_CDISC|Skin Mixed Basal and Squamous Cell Carcinoma|8095/3
C0007118|T191|PT|BB35.|RCD|Basosquamous carcinoma|8095/3
C0007118|T191|PT|X78ST|RCD|Basosquamous carcinoma of skin|8095/3
C0007118|T191|SY|X78ST|RCD|BCC - Metatypical basal cell carcinoma of skin|8095/3
C0007118|T191|SY|X78ST|RCD|Metatypical basal cell carcinoma of skin|8095/3
C0007118|T191|AB|X78ST|RCD|Metatypical BCC of skin|8095/3
C0007118|T191|PT|BB36.|RCD|Metatypical carcinoma|8095/3
C0007118|T191|AB|BB35.|RCD|Mixed basal - squamous cell ca|8095/3
C0007118|T191|SY|BB35.|RCD|Mixed basal - squamous cell carcinoma|8095/3
C0007118|T191|SY|37304002|SNOMEDCT_US|Basisquamous cell carcinoma|8095/3
C0007118|T191|PT|37304002|SNOMEDCT_US|Basosquamous carcinoma|8095/3
C0007118|T191|PT|254702000|SNOMEDCT_US|Basosquamous carcinoma of skin|8095/3
C0007118|T191|SY|254702000|SNOMEDCT_US|BCC - Metatypical basal cell carcinoma of skin|8095/3
C0007118|T191|SY|254702000|SNOMEDCT_US|Metatypical basal cell carcinoma of skin|8095/3
C0007118|T191|PT|6641007|SNOMEDCT_US|Metatypical carcinoma|8095/3
C0007118|T191|SY|37304002|SNOMEDCT_US|Mixed basal - squamous cell carcinoma|8095/3
C0007118|T191|SY|37304002|SNOMEDCT_US|Mixed basal-squamous cell carcinoma|8095/3
C2937231|T191|PN|NOCODE|MTH|Intraepidermal epithelioma of Jadassohn|8096/0
C2937231|T191|OP|C4110|NCI|Borst-Jadassohn Intraepidermal Carcinoma|8096/0
C2937231|T191|PT|C4110|NCI|Intraepidermal Epithelioma of Jadassohn|8096/0
C2937231|T191|OP|C4110|NCI|Intraepidermal Epithelioma of Jadassohn|8096/0
C2937231|T191|AB|XM1F8|RCD|Borst-Jadassohn intraepid ca|8096/0
C2937231|T191|SY|XM1F8|RCD|Borst-Jadassohn intraepidermal carcinoma|8096/0
C2937231|T191|SY|XM1F8|RCD|Borst-Jadassohn phenomenon|8096/0
C2937231|T191|AB|XM1F8|RCD|Clonal intraepidermal carcinom|8096/0
C2937231|T191|SY|XM1F8|RCD|Clonal intraepidermal carcinoma|8096/0
C2937231|T191|AB|XM1F8|RCD|Intraep epithelio of Jadassohn|8096/0
C2937231|T191|AB|XM1F8|RCD|Intraepi epithelioma Borsst-J|8096/0
C2937231|T191|SY|XM1F8|RCD|Intraepidermal epithelioma of Borsst-Jadassohn|8096/0
C2937231|T191|PT|XM1F8|RCD|Intraepidermal epithelioma of Jadassohn|8096/0
C2937231|T191|OA|BB37.|RCDSY|Intraepid.epith.- Jadassohn|8096/0
C2937231|T191|OP|BB37.|RCDSY|Intraepidermal epithelioma of Jadassohn|8096/0
C2937231|T191|SY|274897005|SNOMEDCT_US|Borst-Jadassohn intraepidermal carcinoma|8096/0
C2937231|T191|SY|274897005|SNOMEDCT_US|Borst-Jadassohn phenomenon|8096/0
C2937231|T191|SY|274897005|SNOMEDCT_US|Clonal intraepidermal carcinoma|8096/0
C2937231|T191|IS|274897005|SNOMEDCT_US|Intraepidermal epithelioma of Borsst-Jadassohn|8096/0
C2937231|T191|SY|274897005|SNOMEDCT_US|Intraepidermal epithelioma of Borst-Jadassohn|8096/0
C2937231|T191|PT|274897005|SNOMEDCT_US|Intraepidermal epithelioma of Jadassohn|8096/0
C2937231|T191|PT|39332000|SNOMEDCT_US|Intraepidermal epithelioma of Jadassohn|8096/0
C4083056|T191|SY|0000057721|CHV|basal cell carcinoma nodular|8097/3
C4083056|T191|PT|0000057721|CHV|nodular basal cell carcinoma|8097/3
C1367861|T191|LLT|10073092|MDR|Micronodular basal cell carcinoma|8097/3
C4083056|T191|LLT|10073093|MDR|Nodular basal cell carcinoma|8097/3
C1367861|T191|PT|352407|MEDCIN|Basal cell carcinoma - micronodular|8097/3
C1879347|T191|PT|355695|MEDCIN|Circumscribed solid basal cell carcinoma|8097/3
C1367861|T191|SY|352407|MEDCIN|malignant neoplasm carcinoma basal cell micronodular|8097/3
C1879347|T191|SY|355695|MEDCIN|skin neoplasm malignant carcinoma basal cell circumscribed solid|8097/3
C4083056|T191|PN|NOCODE|MTH|Basal cell carcinoma, nodular|8097/3
C1879347|T191|PN|NOCODE|MTH|Skin Nodular Solid Basal Cell Carcinoma|8097/3
C1367861|T191|SY|C27541|NCI|Micronodular Basal Cell Carcinoma|8097/3
C1367861|T191|PT|C27541|NCI|Skin Micronodular Basal Cell Carcinoma|8097/3
C1879347|T191|PT|C5616|NCI|Skin Nodular Solid Basal Cell Carcinoma|8097/3
C1367861|T191|PT|402529002|SNOMEDCT_US|Basal cell carcinoma - micronodular|8097/3
C1367861|T191|IS|128636006|SNOMEDCT_US|Basal cell carcinoma, micronodular|8097/3
C1367861|T191|PT|400071004|SNOMEDCT_US|Basal cell carcinoma, micronodular|8097/3
C4083056|T191|PT|128636006|SNOMEDCT_US|Basal cell carcinoma, nodular|8097/3
C1879347|T191|PT|403910009|SNOMEDCT_US|Circumscribed solid basal cell carcinoma|8097/3
C4083056|T191|IS|403910009|SNOMEDCT_US|Nodular basal cell carcinoma|8097/3
C1304296|T191|PT|352403|MEDCIN|Basal cell carcinoma - adenoid|8098/3
C1304296|T191|SY|352403|MEDCIN|malignant neoplasm carcinoma basal cell adenoid|8098/3
C1304296|T191|SY|C27535|NCI|Adenoid Basal Cell Carcinoma|8098/3
C1304296|T191|PT|C27535|NCI|Skin Adenoid Basal Cell Carcinoma|8098/3
C1266007|T191|PT|128637002|SNOMEDCT_US|Adenoid basal carcinoma|8098/3
C1304296|T191|PT|402525008|SNOMEDCT_US|Basal cell carcinoma - adenoid|8098/3
C0349658|T191|SY|0000029944|CHV|epithelioma adenoides cysticum|8100/0
C0349658|T191|PT|0000029944|CHV|trichoepithelioma|8100/0
C0349658|T191|SY|0000029944|CHV|trichoepitheliomas|8100/0
C0349658|T191|PT|HP:0025367|HPO|Trichoepithelioma|8100/0
C0349658|T191|PT|10015106|MDR|Epithelioma adenoides cysticum|8100/0
C0349658|T191|LLT|10015106|MDR|Epithelioma adenoides cysticum|8100/0
C0349658|T191|LLT|10063951|MDR|Trichoblastoma|8100/0
C0349658|T191|LLT|10044610|MDR|Trichoepithelioma|8100/0
C0349658|T191|PT|312994|MEDCIN|trichoepithelioma|8100/0
C0349658|T191|PN|NOCODE|MTH|Trichoepithelioma|8100/0
C0349658|T191|SY|C27132|NCI|Brooke's Tumor|8100/0
C0349658|T191|PT|C27132|NCI|Trichoblastoma|8100/0
C0349658|T191|SY|C27132|NCI|Trichoepithelioma|8100/0
C0349658|T191|SY|C27132|NCI|Trichogenic Adnexal Tumor|8100/0
C0349658|T191|SY|C27132|NCI|Trichogenic Trichoblastoma|8100/0
C0349658|T191|SY|C27132|NCI_CDISC|Brooke's Tumor|8100/0
C0349658|T191|SY|C27132|NCI_CDISC|Trichoepithelioma|8100/0
C0349658|T191|PT|C27132|NCI_CDISC|TRICHOEPITHELIOMA, BENIGN|8100/0
C0349658|T191|SY|C27132|NCI_CDISC|Trichogenic Adnexal Tumor|8100/0
C0349658|T191|SY|C27132|NCI_CDISC|Trichogenic Trichoblastoma|8100/0
C0349658|T191|SY|XM1F9|RCD|Brooke's tumour|8100/0
C0349658|T191|SY|XM1F9|RCD|Epithelioma adenoides cysticum|8100/0
C0349658|T191|PT|Xa0ZO|RCD|Trichoblastoma|8100/0
C0349658|T191|PT|XM1F9|RCD|Trichoepithelioma|8100/0
C0349658|T191|SY|XM1F9|RCDAE|Brooke's tumor|8100/0
C0349658|T191|OP|BB38.|RCDSY|Trichoepithelioma|8100/0
C0349658|T191|SY|59186007|SNOMEDCT_US|Brooke's tumor|8100/0
C0349658|T191|SY|274898000|SNOMEDCT_US|Brooke's tumor|8100/0
C0349658|T191|SYGB|59186007|SNOMEDCT_US|Brooke's tumour|8100/0
C0349658|T191|SYGB|274898000|SNOMEDCT_US|Brooke's tumour|8100/0
C0349658|T191|SY|59186007|SNOMEDCT_US|Epithelioma adenoides cysticum|8100/0
C0349658|T191|SY|274898000|SNOMEDCT_US|Epithelioma adenoides cysticum|8100/0
C0349658|T191|PT|277942005|SNOMEDCT_US|Trichoblastoma|8100/0
C0349658|T191|PT|59186007|SNOMEDCT_US|Trichoepithelioma|8100/0
C0349658|T191|PT|274898000|SNOMEDCT_US|Trichoepithelioma|8100/0
C0334262|T191|PT|0000029945|CHV|trichofolliculoma|8101/0
C0334262|T191|LLT|10044611|MDR|Trichofolliculoma|8101/0
C0334262|T191|CE|C536553|MSH|Recurrent trichofolliculoma|8101/0
C0334262|T191|NM|C536553|MSH|Trichofolliculoma|8101/0
C0334262|T191|PN|NOCODE|MTH|Trichofolliculoma|8101/0
C0334262|T191|PT|C4112|NCI|Trichofolliculoma|8101/0
C0334262|T191|PT|XM1FA|RCD|Trichofolliculoma|8101/0
C0334262|T191|OP|BB39.|RCDSY|Trichofolliculoma|8101/0
C0334262|T191|PT|33059009|SNOMEDCT_US|Trichofolliculoma|8101/0
C0334262|T191|PT|274899008|SNOMEDCT_US|Trichofolliculoma|8101/0
C0334263|T191|PT|0000029946|CHV|trichilemmoma|8102/0
C0334263|T191|SY|0000029946|CHV|trichilemmomas|8102/0
C0334263|T191|SY|0000029946|CHV|tricholemmoma|8102/0
C0334263|T191|SY|0000029946|CHV|tricholemmomas|8102/0
C0334263|T191|PT|HP:0012844|HPO|Trichilemmoma|8102/0
C0334263|T191|SY|HP:0012844|HPO|Tricholemmoma|8102/0
C0334263|T191|LLT|10057991|MDR|Trichilemmoma|8102/0
C0334263|T191|LLT|10044612|MDR|Tricholemmoma|8102/0
C0334263|T191|PT|C4113|NCI|Trichilemmoma|8102/0
C0334263|T191|SY|C4113|NCI|Tricholemmoma|8102/0
C0334263|T191|PT|C4113|NCI_CDISC|TRICHOLEMMOMA, BENIGN|8102/0
C0334263|T191|PT|XM1FB|RCD|Tricholemmoma|8102/0
C0334263|T191|OP|BB3A.|RCDSY|Tricholemmoma|8102/0
C0334263|T191|PT|46199002|SNOMEDCT_US|Trichilemmoma|8102/0
C0334263|T191|PT|274900003|SNOMEDCT_US|Trichilemmoma|8102/0
C0334263|T191|SY|46199002|SNOMEDCT_US|Tricholemmoma|8102/0
C0334263|T191|SY|274900003|SNOMEDCT_US|Tricholemmoma|8102/0
C0334263|T191|PT|0000029946|CHV|trichilemmoma|8102/2
C0334263|T191|SY|0000029946|CHV|trichilemmomas|8102/2
C0334263|T191|SY|0000029946|CHV|tricholemmoma|8102/2
C0334263|T191|SY|0000029946|CHV|tricholemmomas|8102/2
C0334263|T191|PT|HP:0012844|HPO|Trichilemmoma|8102/2
C0334263|T191|SY|HP:0012844|HPO|Tricholemmoma|8102/2
C0334263|T191|LLT|10057991|MDR|Trichilemmoma|8102/2
C0334263|T191|LLT|10044612|MDR|Tricholemmoma|8102/2
C0334263|T191|PT|C4113|NCI|Trichilemmoma|8102/2
C0334263|T191|SY|C4113|NCI|Tricholemmoma|8102/2
C0334263|T191|PT|C4113|NCI_CDISC|TRICHOLEMMOMA, BENIGN|8102/2
C0334263|T191|PT|XM1FB|RCD|Tricholemmoma|8102/2
C0334263|T191|OP|BB3A.|RCDSY|Tricholemmoma|8102/2
C0334263|T191|PT|274900003|SNOMEDCT_US|Trichilemmoma|8102/2
C0334263|T191|PT|46199002|SNOMEDCT_US|Trichilemmoma|8102/2
C0334263|T191|SY|46199002|SNOMEDCT_US|Tricholemmoma|8102/2
C0334263|T191|SY|274900003|SNOMEDCT_US|Tricholemmoma|8102/2
C1266009|T191|SY|355112|MEDCIN|skin neoplasm malignant trichilemmal carcinoma|8102/3
C1266009|T191|PT|355112|MEDCIN|Trichilemmal carcinoma|8102/3
C1266009|T191|SY|C43326|NCI|Trichilemmal Carcinoma|8102/3
C1266009|T191|PT|C43326|NCI|Trichilemmocarcinoma|8102/3
C1266009|T191|SY|128624000|SNOMEDCT_US|Trichilemmal carcinoma|8102/3
C1266009|T191|PT|403929003|SNOMEDCT_US|Trichilemmal carcinoma|8102/3
C1266009|T191|PT|128624000|SNOMEDCT_US|Trichilemmocarcinoma|8102/3
C0345992|T191|PT|0000031036|CHV|pilar tumor|8103/0
C0345992|T191|SY|0000031036|CHV|pilar tumors|8103/0
C0345992|T191|SY|0000031036|CHV|proliferating trichilemmal cyst|8103/0
C0345992|T191|PN|NOCODE|MTH|Pilar tumor|8103/0
C0345992|T191|ET|704.42|MTHICD9|Trichilemmal proliferating cyst|8103/0
C0345992|T191|SY|C27125|NCI|Pilar Cyst|8103/0
C0345992|T191|SY|C27125|NCI|Pilar Tumor|8103/0
C0345992|T191|PT|C27125|NCI|Proliferating Pilar Tumor|8103/0
C0345992|T191|SY|C27125|NCI|Proliferating Trichilemmal Cyst|8103/0
C0345992|T191|SY|C27125|NCI|Proliferating Trichilemmal Tumor|8103/0
C0345992|T191|SY|C27125|NCI|Proliferating Tricholemmal Tumor|8103/0
C0345992|T191|AB|X78Ru|RCD|Proliferat trichilemmal cyst|8103/0
C0345992|T191|PT|X78Ru|RCD|Proliferating pilar cyst|8103/0
C0345992|T191|SY|X78Ru|RCD|Proliferating trichilemmal cyst|8103/0
C0345992|T191|SY|419093005|SNOMEDCT_US|Pilar cyst|8103/0
C0345992|T191|PT|128638007|SNOMEDCT_US|Pilar tumor|8103/0
C0345992|T191|PTGB|128638007|SNOMEDCT_US|Pilar tumour|8103/0
C0345992|T191|PT|254678009|SNOMEDCT_US|Proliferating pilar cyst|8103/0
C0345992|T191|SY|128638007|SNOMEDCT_US|Proliferating trichilemmal cyst|8103/0
C0345992|T191|SY|254678009|SNOMEDCT_US|Proliferating trichilemmal cyst|8103/0
C0345992|T191|SY|128638007|SNOMEDCT_US|Proliferating trichilemmal tumor|8103/0
C0345992|T191|SYGB|128638007|SNOMEDCT_US|Proliferating trichilemmal tumour|8103/0
C0345992|T191|SY|128638007|SNOMEDCT_US|Proliferating tricholemmal cyst|8103/0
C0345992|T191|PT|0000031036|CHV|pilar tumor|8103/1
C0345992|T191|SY|0000031036|CHV|pilar tumors|8103/1
C0345992|T191|SY|0000031036|CHV|proliferating trichilemmal cyst|8103/1
C0345992|T191|PN|NOCODE|MTH|Pilar tumor|8103/1
C2959585|T191|PN|NOCODE|MTH|Proliferating trichilemmal tumor|8103/1
C0345992|T191|ET|704.42|MTHICD9|Trichilemmal proliferating cyst|8103/1
C0345992|T191|SY|C27125|NCI|Pilar Cyst|8103/1
C0345992|T191|SY|C27125|NCI|Pilar Tumor|8103/1
C0345992|T191|PT|C27125|NCI|Proliferating Pilar Tumor|8103/1
C0345992|T191|SY|C27125|NCI|Proliferating Trichilemmal Cyst|8103/1
C0345992|T191|SY|C27125|NCI|Proliferating Trichilemmal Tumor|8103/1
C0345992|T191|SY|C27125|NCI|Proliferating Tricholemmal Tumor|8103/1
C0345992|T191|AB|X78Ru|RCD|Proliferat trichilemmal cyst|8103/1
C0345992|T191|PT|X78Ru|RCD|Proliferating pilar cyst|8103/1
C0345992|T191|SY|X78Ru|RCD|Proliferating trichilemmal cyst|8103/1
C0345992|T191|SY|419093005|SNOMEDCT_US|Pilar cyst|8103/1
C0345992|T191|PT|128638007|SNOMEDCT_US|Pilar tumor|8103/1
C0345992|T191|PTGB|128638007|SNOMEDCT_US|Pilar tumour|8103/1
C0345992|T191|PT|254678009|SNOMEDCT_US|Proliferating pilar cyst|8103/1
C0345992|T191|SY|254678009|SNOMEDCT_US|Proliferating trichilemmal cyst|8103/1
C0345992|T191|SY|128638007|SNOMEDCT_US|Proliferating trichilemmal cyst|8103/1
C0345992|T191|SY|128638007|SNOMEDCT_US|Proliferating trichilemmal tumor|8103/1
C2959585|T191|PT|446023005|SNOMEDCT_US|Proliferating trichilemmal tumor|8103/1
C2959585|T191|PTGB|446023005|SNOMEDCT_US|Proliferating trichilemmal tumour|8103/1
C0345992|T191|SYGB|128638007|SNOMEDCT_US|Proliferating trichilemmal tumour|8103/1
C0345992|T191|SY|128638007|SNOMEDCT_US|Proliferating tricholemmal cyst|8103/1
C0206711|T191|SY|0000021039|CHV|calcifying epithelioma malherbe|8110/0
C0206711|T191|SY|0000021039|CHV|pilomatricoma|8110/0
C0206711|T191|SY|0000021039|CHV|pilomatricomas|8110/0
C0206711|T191|PT|0000021039|CHV|pilomatrixoma|8110/0
C0206711|T191|PT|HP:0030434|HPO|Pilomatrixoma|8110/0
C0206711|T191|LLT|10035040|MDR|Pilomatricoma|8110/0
C0206711|T191|ET|D018296|MSH|Benign Pilomatricoma|8110/0
C0206711|T191|ET|D018296|MSH|Benign Pilomatrixoma|8110/0
C0206711|T191|ET|D018296|MSH|Calcifying Epithelioma of Malherbe|8110/0
C0206711|T191|ET|D018296|MSH|Epithelioma Calcificans Of Malherbe|8110/0
C0206711|T191|ET|D018296|MSH|Malherbe Calcifying Epithelioma|8110/0
C0206711|T191|ET|D018296|MSH|Pilomatricoma|8110/0
C0206711|T191|PM|D018296|MSH|Pilomatricoma, Benign|8110/0
C0206711|T191|MH|D018296|MSH|Pilomatrixoma|8110/0
C0206711|T191|PM|D018296|MSH|Pilomatrixoma, Benign|8110/0
C0206711|T191|PN|NOCODE|MTH|Pilomatrixoma|8110/0
C0206711|T191|SY|C7368|NCI|Benign Pilomatricoma|8110/0
C0206711|T191|SY|C7368|NCI|Benign Pilomatrixoma|8110/0
C0206711|T191|SY|C7368|NCI|Calcifying Epithelioma of Malherbe|8110/0
C0206711|T191|PT|C7368|NCI|Pilomatricoma|8110/0
C0206711|T191|SY|C7368|NCI|Pilomatrixoma|8110/0
C0206711|T191|SY|C7368|NCI_CDISC|Benign Hair Follicle Neoplasm|8110/0
C0206711|T191|SY|C7368|NCI_CDISC|Benign Pilomatricoma|8110/0
C0206711|T191|SY|C7368|NCI_CDISC|Benign Pilomatrixoma|8110/0
C0206711|T191|SY|C7368|NCI_CDISC|Calcifying Epitherlioma of Malherbe|8110/0
C0206711|T191|SY|C7368|NCI_CDISC|Pilomatrixoma|8110/0
C0206711|T191|PT|C7368|NCI_CDISC|PILOMATRIXOMA, BENIGN|8110/0
C0206711|T191|AB|XM1FC|RCD|Ben calci epithelioma-Malherbe|8110/0
C0206711|T191|SY|XM1FC|RCD|Benign calcifying epithelioma of Malherbe|8110/0
C0206711|T191|AB|XM1FC|RCD|Calcif epithelioma of Malherbe|8110/0
C0206711|T191|SY|XM1FC|RCD|Calcifying epithelioma of Malherbe|8110/0
C0206711|T191|SY|XM1FC|RCD|Pilomatricoma|8110/0
C0206711|T191|PT|XM1FC|RCD|Pilomatrixoma|8110/0
C0206711|T191|OP|BB3B.|RCDSY|Pilomatrixoma|8110/0
C0206711|T191|SY|44155009|SNOMEDCT_US|Benign calcifying epithelioma|8110/0
C0206711|T191|SY|274901004|SNOMEDCT_US|Benign calcifying epithelioma of Malherbe|8110/0
C0206711|T191|SY|274901004|SNOMEDCT_US|Calcifying epithelioma of Malherbe|8110/0
C0206711|T191|SY|44155009|SNOMEDCT_US|Calcifying epithelioma of Malherbe|8110/0
C5230949|T191|PT|816971006|SNOMEDCT_US|Melanocytic matricoma|8110/0
C0206711|T191|SY|44155009|SNOMEDCT_US|Pilomatricoma|8110/0
C0206711|T191|SY|274901004|SNOMEDCT_US|Pilomatricoma|8110/0
C0206711|T191|PT|274901004|SNOMEDCT_US|Pilomatrixoma|8110/0
C0206711|T191|PT|44155009|SNOMEDCT_US|Pilomatrixoma|8110/0
C0206711|T191|IS|44155009|SNOMEDCT_US|Pilomatrixoma, NOS|8110/0
C0585475|T191|LLT|10075614|MDR|Pilomatrix carcinoma|8110/3
C0585475|T191|PT|10075614|MDR|Pilomatrix carcinoma|8110/3
C0585475|T191|PT|231610|MEDCIN|pilomatrix carcinoma of skin|8110/3
C0585475|T191|SY|C4114|NCI|Invasive Pilomatrixoma|8110/3
C0585475|T191|SY|C4114|NCI|Matrical Carcinoma|8110/3
C0585475|T191|PT|C4114|NCI|Pilomatrical Carcinoma|8110/3
C0585475|T191|SY|C4114|NCI|Pilomatrix Carcinoma|8110/3
C0585475|T191|SY|C4114|NCI|Pilomatrix Carcinoma of Skin|8110/3
C0585475|T191|SY|C4114|NCI|Pilomatrix Carcinoma of the Skin|8110/3
C0585475|T191|SY|C4114|NCI|Pilomatrix Skin Carcinoma|8110/3
C0585475|T191|SY|X77nB|RCD|Malignant pilomatrixoma|8110/3
C0585475|T191|PT|X77nB|RCD|Pilomatrix carcinoma|8110/3
C0585475|T191|PT|XaBB4|RCD|Pilomatrix carcinoma of skin|8110/3
C0585475|T191|SY|24762001|SNOMEDCT_US|Malignant pilomatrixoma|8110/3
C0585475|T191|SY|24762001|SNOMEDCT_US|Matrical carcinoma|8110/3
C0585475|T191|SY|24762001|SNOMEDCT_US|Pilomatricoma, malignant|8110/3
C0585475|T191|PT|24762001|SNOMEDCT_US|Pilomatrix carcinoma|8110/3
C0585475|T191|PT|307610008|SNOMEDCT_US|Pilomatrix carcinoma of skin|8110/3
C0585475|T191|SY|24762001|SNOMEDCT_US|Pilomatrixoma, malignant|8110/3
C0334266|T191|PT|C4115|NCI|Transitional Cell Papilloma|8120/0
C0334266|T191|SY|C4115|NCI|Transitional Papilloma|8120/0
C0334266|T191|PT|C4115|NCI_CDISC|PAPILLOMA, TRANSITIONAL CELL, BENIGN|8120/0
C0334266|T191|SY|C4115|NCI_CDISC|Transitional Papilloma|8120/0
C0334266|T191|PT|Xa98I|RCD|Transitional cell papilloma|8120/0
C0334266|T191|SY|Xa98I|RCD|Transitional papilloma|8120/0
C0334266|T191|OA|BB40.|RCDSY|Transit.cell papilloma NOS|8120/0
C0334266|T191|OP|BB40.|RCDSY|Transitional cell papilloma NOS|8120/0
C0334266|T191|SY|45083001|SNOMEDCT_US|Transitional cell papilloma|8120/0
C0334266|T191|PT|44342003|SNOMEDCT_US|Transitional cell papilloma, benign|8120/0
C0334266|T191|IS|44342003|SNOMEDCT_US|Transitional cell papilloma, NOS|8120/0
C0334266|T191|SY|44342003|SNOMEDCT_US|Transitional papilloma|8120/0
C0235754|T191|PT|0000023601|CHV|bladder papilloma|8120/1
C0235754|T191|SY|0000023601|CHV|bladder wart|8120/1
C0235754|T191|SY|0000023601|CHV|bladder warts|8120/1
C0235754|T191|SY|0000023601|CHV|papilloma bladder|8120/1
C0235754|T191|SY|0000023601|CHV|papilloma of bladder|8120/1
C0235754|T191|SY|0000023601|CHV|papilloma urinary bladder|8120/1
C0235754|T191|GT|NEOPL BLADDER|CST|BLADDER PAPILLOMA|8120/1
C0235754|T191|DI|U000221|DXP|BLADDER, PAPILLOMA|8120/1
C0235754|T191|PT|MTHU011081|ICPC2ICD10ENG|bladder; papilloma|8120/1
C0235754|T191|PT|MTHU057335|ICPC2ICD10ENG|papilloma; bladder|8120/1
C0235754|T191|PTN|U78006|ICPC2P|bladder papillomata|8120/1
C0235754|T191|PT|U78006|ICPC2P|Papillomata;bladder|8120/1
C0235754|T191|LLT|10005064|MDR|Bladder papilloma|8120/1
C0235754|T191|PT|10005064|MDR|Bladder papilloma|8120/1
C0235754|T191|LLT|10005086|MDR|Bladder wart|8120/1
C0235754|T191|LLT|10033717|MDR|Papilloma of bladder|8120/1
C0235754|T191|PN|NOCODE|MTH|Bladder papilloma|8120/1
C0235754|T191|PT|C3842|NCI|Urothelial Papilloma|8120/1
C0235754|T191|SY|BB41.|RCD|Papilloma of bladder|8120/1
C0235754|T191|SY|BB41.|RCD|Urinary bladder papilloma|8120/1
C0235754|T191|PT|BB41.|RCD|Urothelial papilloma|8120/1
C0235754|T191|OAS|269642004|SNOMEDCT_US|Bladder papilloma NOS|8120/1
C0235754|T191|OAS|154620001|SNOMEDCT_US|Bladder papilloma NOS|8120/1
C0235754|T191|OAP|313414002|SNOMEDCT_US|Bladder papilloma NOS|8120/1
C0235754|T191|OAS|154620001|SNOMEDCT_US|Papilloma bladder NOS|8120/1
C0235754|T191|OAS|269642004|SNOMEDCT_US|Papilloma bladder NOS|8120/1
C0235754|T191|SY|45083001|SNOMEDCT_US|Papilloma of bladder|8120/1
C0235754|T191|SY|45083001|SNOMEDCT_US|Papilloma of urinary bladder|8120/1
C0235754|T191|SY|45083001|SNOMEDCT_US|Urinary bladder papilloma|8120/1
C0235754|T191|PT|45083001|SNOMEDCT_US|Urothelial papilloma|8120/1
C0235754|T191|PT|0765|WHO|BLADDER PAPILLOMA|8120/1
C0334267|T191|PT|271384|MEDCIN|transitional cell carcinoma in situ|8120/2
C0334267|T191|PN|NOCODE|MTH|Transitional cell carcinoma in situ|8120/2
C0334267|T191|PT|C4116|NCI|Stage 0 Transitional Cell Carcinoma|8120/2
C0334267|T191|SY|C4116|NCI|Transitional Carcinoma in situ|8120/2
C0334267|T191|SY|C4116|NCI|Transitional Cell Carcinoma in situ|8120/2
C0334267|T191|AB|BB42.|RCD|Transit cell carcinoma in situ|8120/2
C0334267|T191|PT|BB42.|RCD|Transitional cell carcinoma in situ|8120/2
C0334267|T191|PT|53530009|SNOMEDCT_US|Transitional cell carcinoma in situ|8120/2
C0334267|T191|IS|53530009|SNOMEDCT_US|Urothelial carcinoma in situ|8120/2
C0334267|T191|SY|53530009|SNOMEDCT_US|Urothelial carcinoma in situ|8120/2
C0007138|T191|PT|0012180|CCPSS|TRANSITIONAL CELL CARCINOMA|8120/3
C0007138|T191|SY|0000002438|CHV|carcinoma cell transitional|8120/3
C0007138|T191|SY|0000002438|CHV|carcinomas urothelial|8120/3
C0007138|T191|SY|0000002438|CHV|transitional carcinoma|8120/3
C0007138|T191|PT|0000002438|CHV|transitional cell carcinoma|8120/3
C0007138|T191|SY|0000002438|CHV|transitional cell carcinomas|8120/3
C0007138|T191|SY|0000002438|CHV|urothelial carcinoma|8120/3
C0007138|T191|PT|2000-9838|CSP|transitional cell carcinoma|8120/3
C0007138|T191|GT|CARCINOMA|CST|CARCINOMA TRANSITIONAL CELL|8120/3
C0007138|T191|PT|A79011|ICPC2P|Transitional cell carcinoma|8120/3
C0007138|T191|PTN|A79011|ICPC2P|transitional cell carcinoma|8120/3
C0007138|T191|LLT|10007477|MDR|Carcinoma transitional cell|8120/3
C0007138|T191|LLT|10044412|MDR|Transitional cell carcinoma|8120/3
C0007138|T191|PT|10044412|MDR|Transitional cell carcinoma|8120/3
C0007138|T191|LLT|10064467|MDR|Urothelial carcinoma|8120/3
C0007138|T191|PT|271430|MEDCIN|transitional cell carcinoma|8120/3
C0007138|T191|MH|D002295|MSH|Carcinoma, Transitional Cell|8120/3
C0007138|T191|PM|D002295|MSH|Carcinomas, Transitional Cell|8120/3
C0007138|T191|PM|D002295|MSH|Cell Carcinoma, Transitional|8120/3
C0007138|T191|PM|D002295|MSH|Cell Carcinomas, Transitional|8120/3
C0007138|T191|PM|D002295|MSH|Transitional Cell Carcinoma|8120/3
C0007138|T191|PM|D002295|MSH|Transitional Cell Carcinomas|8120/3
C0007138|T191|PN|NOCODE|MTH|Carcinoma, Transitional Cell|8120/3
C0007138|T191|SY|C2930|NCI|Transitional Carcinoma|8120/3
C0007138|T191|PT|C2930|NCI|Transitional Cell Carcinoma|8120/3
C0007138|T191|PT|C2930|NCI_CDISC|CARCINOMA, UROTHELIAL, MALIGNANT|8120/3
C0007138|T191|SY|C2930|NCI_CDISC|Transitional Cell Carcinoma|8120/3
C0007138|T191|PT|C2930|NCI_CPTAC|Transitional Cell Carcinoma|8120/3
C0007138|T191|PT|CDR0000046629|NCI_NCI-GLOSS|transitional cell carcinoma|8120/3
C0007138|T191|PT|C2930|NCI_NICHD|Transitional Cell Carcinoma|8120/3
C0007138|T191|SY|Xa98J|RCD|TCC - Transitional cell carcinoma|8120/3
C0007138|T191|AB|Xa98J|RCD|TCC-Transitionl cell carcinoma|8120/3
C0007138|T191|SY|Xa98J|RCD|Transitional carcinoma|8120/3
C0007138|T191|PT|Xa98J|RCD|Transitional cell carcinoma|8120/3
C0007138|T191|SY|Xa98J|RCD|Urothelial carcinoma|8120/3
C0007138|T191|OA|BB43.|RCDSY|Transitional cell ca. NOS|8120/3
C0007138|T191|OP|BB43.|RCDSY|Transitional cell carcinoma NOS|8120/3
C3164997|T191|PT|449330007|SNOMEDCT_US|Papillary and solid transitional cell carcinoma|8120/3
C0007138|T191|SY|27090000|SNOMEDCT_US|TCC - Transitional cell carcinoma|8120/3
C0007138|T191|SY|27090000|SNOMEDCT_US|Transitional carcinoma|8120/3
C3164997|T191|SY|449330007|SNOMEDCT_US|Transitional carcinoma with mixed papillary and solid growth pattern|8120/3
C0007138|T191|PT|27090000|SNOMEDCT_US|Transitional cell carcinoma|8120/3
C1302510|T191|PT|399564007|SNOMEDCT_US|Transitional cell carcinoma with glandular differentiation|8120/3
C1302431|T191|PT|399464005|SNOMEDCT_US|Transitional cell carcinoma with squamous differentiation|8120/3
C0007138|T191|IS|27090000|SNOMEDCT_US|Transitional cell carcinoma, NOS|8120/3
C0007138|T191|SY|27090000|SNOMEDCT_US|Urothelial carcinoma|8120/3
C0334268|T191|PT|0000029947|CHV|schneiderian papilloma|8121/0
C0334268|T191|SY|0000029947|CHV|sinonasal papilloma|8121/0
C0334268|T191|LLT|10082317|MDR|Schneiderian papilloma|8121/0
C0334268|T191|LLT|10071665|MDR|Sinonasal papilloma|8121/0
C0334268|T191|PT|10071665|MDR|Sinonasal papilloma|8121/0
C1334282|T191|SY|C6192|NCI|Inverted Papilloma of Urinary Tract|8121/0
C1334282|T191|PT|C6192|NCI|Inverted Urothelial Papilloma|8121/0
C0334268|T191|PT|C4117|NCI|Schneiderian Papilloma|8121/0
C1334282|T191|SY|C6192|NCI|Urinary Tract Inverted Papilloma|8121/0
C0334268|T191|PT|BB44.|RCD|Schneiderian papilloma|8121/0
C5231008|T191|PT|818961002|SNOMEDCT_US|Benign columnar cell papilloma|8121/0
C5231007|T191|PT|818960001|SNOMEDCT_US|Benign cylindrical cell papilloma|8121/0
C5231003|T191|SY|818956004|SNOMEDCT_US|Benign exophytic sinonasal papilloma|8121/0
C5231003|T191|SY|818956004|SNOMEDCT_US|Benign fungiform sinonasal papilloma|8121/0
C0334268|T191|PT|818954001|SNOMEDCT_US|Benign inverted transitional cell papilloma|8121/0
C0334268|T191|SY|818954001|SNOMEDCT_US|Benign inverted transitional papilloma|8121/0
C5231003|T191|SY|818956004|SNOMEDCT_US|Benign Schneiderian papilloma|8121/0
C5231003|T191|PT|818956004|SNOMEDCT_US|Benign sinonasal papilloma|8121/0
C5231003|T191|SY|818956004|SNOMEDCT_US|Benign sinonasal papilloma, exophytic|8121/0
C5231003|T191|SY|818956004|SNOMEDCT_US|Benign sinonasal papilloma, fungiform|8121/0
C0334268|T191|SY|818954001|SNOMEDCT_US|Benign transitional cell papilloma, inverted|8121/0
C0334268|T191|SY|818954001|SNOMEDCT_US|Benign transitional papilloma, inverted|8121/0
C1334282|T191|PT|733845009|SNOMEDCT_US|Inverted urothelial papilloma|8121/0
C0334268|T191|OAP|50894008|SNOMEDCT_US|Schneiderian papilloma|8121/0
C0334268|T191|OAS|50894008|SNOMEDCT_US|Sinonasal papilloma|8121/0
C0334268|T191|OAS|50894008|SNOMEDCT_US|Sinonasal papilloma, exophytic|8121/0
C0334268|T191|OAS|50894008|SNOMEDCT_US|Sinonasal papilloma, fungiform|8121/0
C0334268|T191|OAS|50894008|SNOMEDCT_US|Transitional cell papilloma, inverted, benign|8121/0
C0334268|T191|OAS|50894008|SNOMEDCT_US|Transitional papilloma, inverted, benign|8121/0
C0334269|T191|SY|0000029948|CHV|columnar cell papilloma|8121/1
C0334269|T191|PT|0000029948|CHV|cylindrical cell papilloma|8121/1
C0334269|T191|PT|C4118|NCI|Inverted Transitional Cell Papilloma|8121/1
C0334269|T191|SY|C4118|NCI|Inverted Transitional Papilloma|8121/1
C0334269|T191|AB|BB45.|RCD|Invert transit cell papilloma|8121/1
C0334269|T191|PT|BB45.|RCD|Inverted transitional cell papilloma|8121/1
C0334269|T191|IS|46580000|SNOMEDCT_US|Columnar cell papilloma|8121/1
C5231004|T191|PT|818957008|SNOMEDCT_US|Columnar cell papilloma uncertain whether benign or malignant|8121/1
C0334269|T191|IS|46580000|SNOMEDCT_US|Cylindrical cell papilloma|8121/1
C5231005|T191|PT|818958003|SNOMEDCT_US|Cylindrical cell papilloma uncertain whether benign or malignant|8121/1
C5231002|T191|PT|818955000|SNOMEDCT_US|Inverted sinonasal papilloma uncertain whether benign or malignant|8121/1
C0334269|T191|IS|46580000|SNOMEDCT_US|Inverted transitional cell papilloma|8121/1
C0334269|T191|PT|46580000|SNOMEDCT_US|Inverted transitional cell papilloma uncertain whether benign or malignant|8121/1
C0334269|T191|SY|46580000|SNOMEDCT_US|Inverted transitional papilloma uncertain whether benign or malignant|8121/1
C5231002|T191|SY|818955000|SNOMEDCT_US|Oncocytic Schneiderian papilloma uncertain whether benign or malignant|8121/1
C5231002|T191|SY|818955000|SNOMEDCT_US|Schneiderian papilloma, oncocytic, uncertain whether benign or malignant|8121/1
C5231002|T191|SY|818955000|SNOMEDCT_US|Sinonasal papilloma, inverted, uncertain whether benign or malignant|8121/1
C0334269|T191|IS|46580000|SNOMEDCT_US|Transitional cell papilloma, inverted|8121/1
C0334269|T191|SY|46580000|SNOMEDCT_US|Transitional cell papilloma, inverted, uncertain whether benign or malignant|8121/1
C0334269|T191|IS|46580000|SNOMEDCT_US|Transitional papilloma, inverted|8121/1
C0334269|T191|SY|46580000|SNOMEDCT_US|Transitional papilloma, inverted, uncertain whether benign or malignant|8121/1
C0334270|T191|SY|271434|MEDCIN|malignant neoplasm carcinoma Schneiderian|8121/3
C0334270|T191|PT|271434|MEDCIN|Schneiderian carcinoma|8121/3
C0334270|T191|PT|C54287|NCI|Non-Keratinizing Sinonasal Squamous Cell Carcinoma|8121/3
C0334270|T191|SY|C54287|NCI|Ringertz Carcinoma|8121/3
C0334270|T191|SY|C54287|NCI|Schneiderian Carcinoma|8121/3
C0334270|T191|SY|C54287|NCI|Sinonasal Cylindrical Cell Carcinoma|8121/3
C0334270|T191|SY|C54287|NCI|Sinonasal Schneiderian Carcinoma|8121/3
C0334270|T191|SY|C54287|NCI|Sinonasal Transitional Cell Carcinoma|8121/3
C0334270|T191|PT|BB46.|RCD|Schneiderian carcinoma|8121/3
C0334270|T191|SY|5600009|SNOMEDCT_US|Cylindrical cell carcinoma|8121/3
C0334270|T191|PT|5600009|SNOMEDCT_US|Schneiderian carcinoma|8121/3
C0334271|T191|PT|271431|MEDCIN|spindle cell transitional cell carcinoma|8122/3
C0334271|T191|SY|271431|MEDCIN|transitional cell carcinoma, spindle cell|8122/3
C0334271|T191|PT|C4120|NCI|Sarcomatoid Transitional Cell Carcinoma|8122/3
C0334271|T191|SY|C4120|NCI|Transitional Cell Spindle Cell Carcinoma|8122/3
C0334271|T191|SY|C4120|NCI|Transitional Spindle Cell Carcinoma|8122/3
C0334271|T191|AB|BB47.|RCD|Transit cell ca-spindle cell|8122/3
C0334271|T191|PT|BB47.|RCD|Transitional cell carcinoma - spindle cell|8122/3
C0334271|T191|SY|112676006|SNOMEDCT_US|Transitional cell carcinoma - spindle cell|8122/3
C0334271|T191|SY|112676006|SNOMEDCT_US|Transitional cell carcinoma, sarcomatoid|8122/3
C0334271|T191|PT|112676006|SNOMEDCT_US|Transitional cell carcinoma, spindle cell|8122/3
C1704216|T191|PT|0000029949|CHV|basaloid carcinoma|8123/3
C1704216|T191|SY|0000029949|CHV|carcinoma basaloid|8123/3
C1704216|T191|PT|271435|MEDCIN|basaloid carcinoma|8123/3
C1704216|T191|SY|TCGA|NCI|Basaloid Carcinoma|8123/3
C1704216|T191|PT|C4121|NCI|Basaloid Carcinoma|8123/3
C1704216|T191|PT|C4121|NCI_CPTAC|Basaloid Carcinoma|8123/3
C1704216|T191|PT|BB48.|RCD|Basaloid carcinoma|8123/3
C1704216|T191|PT|5843004|SNOMEDCT_US|Basaloid carcinoma|8123/3
C0334273|T191|PT|271436|MEDCIN|cloacogenic carcinoma|8124/3
C0334273|T191|PT|217583|MEDCIN|cloacogenic carcinoma of anal canal|8124/3
C0334273|T191|PT|217712|MEDCIN|cloacogenic carcinoma of anus|8124/3
C0334273|T191|PCE|C563020|MSH|Cloacogenic Carcinoma|8124/3
C0334273|T191|PT|C8255|NCI|Anal Canal Cloacogenic Carcinoma|8124/3
C0334273|T191|SY|C8255|NCI|Anal Canal Transitional Zone Carcinoma|8124/3
C0334273|T191|SY|C8255|NCI|Anal Cloacogenic Carcinoma|8124/3
C0334273|T191|SY|C8255|NCI|Cloacogenic Anal Carcinoma|8124/3
C0334273|T191|SY|C8255|NCI|Cloacogenic Carcinoma|8124/3
C0334273|T191|SY|C8255|NCI|Cloacogenic Carcinoma of Anus|8124/3
C0334273|T191|SY|C8255|NCI|Cloacogenic Carcinoma of the Anus|8124/3
C0334273|T191|DN|C8255|NCI_CTRP|Anal Canal Cloacogenic Cancer|8124/3
C0334273|T191|SY|CDR0000040845|PDQ|Anal Canal Cloacogenic Carcinoma|8124/3
C0334273|T191|SY|CDR0000040845|PDQ|anal cancer, cloacogenic carcinoma|8124/3
C0334273|T191|SY|CDR0000040845|PDQ|Anal Cloacogenic Carcinoma|8124/3
C0334273|T191|SY|CDR0000040845|PDQ|anus cancer, cloacogenic carcinoma|8124/3
C0334273|T191|SY|CDR0000040845|PDQ|Cloacogenic Anal Carcinoma|8124/3
C0334273|T191|SY|CDR0000040845|PDQ|Cloacogenic Carcinoma|8124/3
C0334273|T191|SY|CDR0000040845|PDQ|Cloacogenic Carcinoma of Anus|8124/3
C0334273|T191|PT|CDR0000040845|PDQ|cloacogenic carcinoma of the anus|8124/3
C0334273|T191|PT|BB49.|RCD|Cloacogenic carcinoma|8124/3
C0334273|T191|PT|84570003|SNOMEDCT_US|Cloacogenic carcinoma|8124/3
C1266010|T191|SY|C27884|NCI|Bladder Papillary Neoplasm of Low Malignant Potential|8130/1
C1266010|T191|SY|C27884|NCI|Bladder Papillary Transitional Cell Neoplasm of Low Malignant Potential|8130/1
C1266010|T191|PT|C27884|NCI|Bladder Papillary Urothelial Neoplasm of Low Malignant Potential|8130/1
C1266010|T191|SY|C27884|NCI|Bladder PUNLMP|8130/1
C1266010|T191|PT|128625004|SNOMEDCT_US|Papillary transitional cell neoplasm of low malignant potential|8130/1
C1266010|T191|SY|128625004|SNOMEDCT_US|Papillary urothelial neoplasm of low malignant potential|8130/1
C1266011|T191|PT|C65181|NCI|Non-Invasive Papillary Transitional Cell Carcinoma|8130/2
C1266011|T191|PT|128877008|SNOMEDCT_US|Papillary transitional cell carcinoma, non-invasive|8130/2
C1266011|T191|SY|128877008|SNOMEDCT_US|Papillary urothelial carcinoma, non-invasive|8130/2
C0334274|T191|PT|271432|MEDCIN|papillary transitional cell carcinoma|8130/3
C0334274|T191|SY|C4122|NCI|Papillary Transitional Carcinoma|8130/3
C0334274|T191|PT|C4122|NCI|Papillary Transitional Cell Carcinoma|8130/3
C0334274|T191|AB|BB4A.|RCD|Papillary transitional cell ca|8130/3
C0334274|T191|PT|BB4A.|RCD|Papillary transitional cell carcinoma|8130/3
C0334274|T191|PT|12400006|SNOMEDCT_US|Papillary transitional cell carcinoma|8130/3
C1266012|T191|SY|271433|MEDCIN|malignant neoplasm carcinoma transitional cell micropapillary|8131/3
C1266012|T191|PT|271433|MEDCIN|micropapillary transitional cell carcinoma|8131/3
C1266012|T191|PT|C65182|NCI|Micropapillary Transitional Cell Carcinoma|8131/3
C1266012|T191|PT|128639004|SNOMEDCT_US|Transitional cell carcinoma, micropapillary|8131/3
C0001430|T191|DE|0000004524|AOD|adenoma|8140/0
C0001430|T191|PT|0011787|CCPSS|ADENOMA NOS|8140/0
C0001430|T191|SY|0000000716|CHV|adenoma|8140/0
C0334684|T191|SY|0000030022|CHV|adenoma renal|8140/0
C0001430|T191|SY|0000000716|CHV|adenomas|8140/0
C0334684|T191|SY|0000053236|CHV|adenomas kidney|8140/0
C0334684|T191|SY|0000030022|CHV|adenomas renal|8140/0
C0001430|T191|SY|0000000716|CHV|benign adenoma|8140/0
C0334684|T191|PT|0000053236|CHV|kidney adenoma|8140/0
C0334684|T191|PT|0000030022|CHV|renal adenoma|8140/0
C0334684|T191|SY|0000030022|CHV|renal cell adenoma|8140/0
C0001430|T191|PT|0000000716|CHV|tumor of the gland|8140/0
C0001430|T191|PT|027|COSTAR|ADENOMA|8140/0
C0001430|T191|PT|2000-1015|CSP|adenoma|8140/0
C0001430|T191|PT|ADENOMA|CST|ADENOMA|8140/0
C0001430|T191|PT|U000067|LCH|Adenoma|8140/0
C0001430|T191|PT|sh85000843|LCH_NW|Adenoma|8140/0
C0001430|T191|LA|LA15390-0|LNC|Adenoma, NOS|8140/0
C0001430|T191|LLT|10001231|MDR|Adenoma|8140/0
C0001430|T191|LLT|10001233|MDR|Adenoma benign|8140/0
C0001430|T191|PT|10001233|MDR|Adenoma benign|8140/0
C0001430|T191|LLT|10001234|MDR|Adenoma benign NOS|8140/0
C0001430|T191|LLT|10001236|MDR|Adenoma NOS|8140/0
C0334684|T191|LLT|10051926|MDR|Kidney adenoma|8140/0
C0334684|T191|LLT|10051948|MDR|Renal adenoma|8140/0
C0334684|T191|PT|10051948|MDR|Renal adenoma|8140/0
C0334684|T191|PT|31537|MEDCIN|adenoma of kidney|8140/0
C0334684|T191|SY|31537|MEDCIN|renal adenoma|8140/0
C0001430|T191|ET|3585|MEDLINEPLUS|Adenoma|8140/0
C0001430|T191|MH|D000236|MSH|Adenoma|8140/0
C0001430|T191|PM|D000236|MSH|Adenomas|8140/0
C0001430|T191|PN|NOCODE|MTH|Adenoma|8140/0
C0334688|T191|PN|NOCODE|MTH|Medullary adenoma|8140/0
C0334684|T191|PN|NOCODE|MTH|Renal Adenoma|8140/0
C0001430|T191|PT|C2855|NCI|Adenoma|8140/0
C0334684|T191|PT|C8383|NCI|Kidney Adenoma|8140/0
C0334684|T191|SY|C8383|NCI|Renal Adenoma|8140/0
C0001430|T191|PT|C2855|NCI_CDISC|ADENOMA, BENIGN|8140/0
C0334684|T191|PT|C8383|NCI_CDISC|ADENOMA, RENAL CELL, BENIGN|8140/0
C0334684|T191|SY|C8383|NCI_CDISC|Renal Tubule Adenoma|8140/0
C0001430|T191|PT|CDR0000046217|NCI_NCI-GLOSS|adenoma|8140/0
C0001430|T191|PT|Xa98K|RCD|Adenoma|8140/0
C0001430|T191|OP|BB50.|RCDSY|Adenoma NOS|8140/0
C0001430|T191|SY|443416007|SNOMEDCT_US|Adenoma|8140/0
C0001430|T191|PT|32048006|SNOMEDCT_US|Adenoma|8140/0
C0001430|T191|SY|32048006|SNOMEDCT_US|Adenoma, no subtype|8140/0
C0001430|T191|IS|32048006|SNOMEDCT_US|Adenoma, NOS|8140/0
C0001430|T191|SY|443416007|SNOMEDCT_US|Benign adenoma|8140/0
C0001430|T191|PT|443416007|SNOMEDCT_US|Benign adenomatous neoplasm|8140/0
C0334688|T191|SY|9098000|SNOMEDCT_US|C cell adenoma|8140/0
C4511908|T191|PT|726545001|SNOMEDCT_US|Intestinal-type adenoma|8140/0
C0334690|T191|PT|12583009|SNOMEDCT_US|Lobular adenoma|8140/0
C0334688|T191|PT|9098000|SNOMEDCT_US|Medullary adenoma|8140/0
C0334686|T191|PT|24017008|SNOMEDCT_US|Meibomian adenoma|8140/0
C0334688|T191|SY|9098000|SNOMEDCT_US|Parafollicular cell adenoma|8140/0
C0334684|T191|SY|41627005|SNOMEDCT_US|Renal adenoma|8140/0
C0334684|T191|PT|41627005|SNOMEDCT_US|Renal cell adenoma|8140/0
C1305409|T191|PN|NOCODE|MTH|Atypical adenoma|8140/1
C1305409|T191|PT|C7559|NCI|Atypical Adenoma|8140/1
C1302701|T191|PT|399890002|SNOMEDCT_US|Adenomatous neoplasm of borderline malignancy|8140/1
C1305409|T191|PT|24482001|SNOMEDCT_US|Atypical adenoma|8140/1
C0334276|T191|PT|0000029950|CHV|adenocarcinoma in situ|8140/2
C0334276|T191|SY|0000029950|CHV|adenocarcinoma in-situ|8140/2
C0334276|T191|SY|0000029950|CHV|adenocarcinoma situ|8140/2
C0334276|T191|SY|0000029950|CHV|in situ adenocarcinoma|8140/2
C0334276|T191|PT|271386|MEDCIN|adenocarcinoma in situ|8140/2
C0334276|T191|MH|D065311|MSH|Adenocarcinoma in Situ|8140/2
C0334276|T191|PM|D065311|MSH|Adenocarcinoma in Situs|8140/2
C0334276|T191|ET|D065311|MSH|Adenocarcinoma, Intraepithelial|8140/2
C0334276|T191|ET|D065311|MSH|Adenocarcinoma, Preinvasive|8140/2
C0334276|T191|PM|D065311|MSH|Adenocarcinomas, Intraepithelial|8140/2
C0334276|T191|PM|D065311|MSH|Adenocarcinomas, Preinvasive|8140/2
C0334276|T191|PM|D065311|MSH|in Situ, Adenocarcinoma|8140/2
C0334276|T191|PM|D065311|MSH|Intraepithelial Adenocarcinoma|8140/2
C0334276|T191|PM|D065311|MSH|Intraepithelial Adenocarcinomas|8140/2
C0334276|T191|PM|D065311|MSH|Preinvasive Adenocarcinoma|8140/2
C0334276|T191|PM|D065311|MSH|Preinvasive Adenocarcinomas|8140/2
C0334276|T191|PM|D065311|MSH|Situ, Adenocarcinoma in|8140/2
C0334276|T191|PN|NOCODE|MTH|Adenocarcinoma in Situ|8140/2
C0334276|T191|PT|C4123|NCI|Adenocarcinoma In Situ|8140/2
C0334276|T191|SY|C4123|NCI|Adenocarcinoma in situ|8140/2
C0334276|T191|SY|C4123|NCI|AIS|8140/2
C0334276|T191|PT|BB51.|RCD|Adenocarcinoma in situ|8140/2
C0334276|T191|SY|BB51.|RCD|AIS - Adenocarcinoma in situ|8140/2
C0334276|T191|PT|51642000|SNOMEDCT_US|Adenocarcinoma in situ|8140/2
C0334276|T191|IS|51642000|SNOMEDCT_US|Adenocarcinoma in situ, NOS|8140/2
C0334276|T191|SY|51642000|SNOMEDCT_US|AIS - Adenocarcinoma in situ|8140/2
C0001418|T191|DE|0000004528|AOD|adenocarcinoma|8140/3
C0001418|T191|PT|0062849|CCPSS|ADENOCARCINOMA|8140/3
C0001418|T191|PT|0000000709|CHV|adenocarcinoma|8140/3
C0001418|T191|SY|0000000709|CHV|adenocarcinomas|8140/3
C0001418|T191|PT|026|COSTAR|ADENOCARCINOMA NOS|8140/3
C0001418|T191|PT|2000-0386|CSP|adenocarcinoma|8140/3
C0001418|T191|GT|CARCINOMA|CST|ADENOCARCINOMA|8140/3
C0001418|T191|GT|CARCINOMA|CST|ADENOCARCINOMA NOS|8140/3
C0001418|T191|PT|U000063|LCH|Adenocarcinoma|8140/3
C0001418|T191|PT|sh85000835|LCH_NW|Adenocarcinoma|8140/3
C0001418|T191|LA|LA11900-0|LNC|Adenocarcinoma|8140/3
C0001418|T191|LA|LA26493-9|LNC|Adenocarcinoma, NOS|8140/3
C0001418|T191|LLT|10001141|MDR|Adenocarcinoma|8140/3
C0001418|T191|PT|10001141|MDR|Adenocarcinoma|8140/3
C0001418|T191|LLT|10001166|MDR|Adenocarcinoma NOS|8140/3
C0001418|T191|LLT|10076630|MDR|Carcinoma in adenoma|8140/3
C0001418|T191|PT|271455|MEDCIN|adenocarcinoma|8140/3
C0431095|T191|PT|271466|MEDCIN|adenocarcinoma with metaplasia|8140/3
C0001418|T191|PT|351909|MEDCIN|Malignant adenomatous neoplasm|8140/3
C0001418|T191|MH|D000230|MSH|Adenocarcinoma|8140/3
C0001418|T191|PM|D000230|MSH|Adenocarcinomas|8140/3
C0001418|T191|ET|D000230|MSH|Adenoma, Malignant|8140/3
C0001418|T191|PM|D000230|MSH|Adenomas, Malignant|8140/3
C0001418|T191|PM|D000230|MSH|Malignant Adenoma|8140/3
C0001418|T191|PM|D000230|MSH|Malignant Adenomas|8140/3
C0001418|T191|PN|NOCODE|MTH|Adenocarcinoma|8140/3
C0001418|T191|PT|C2852|NCI|Adenocarcinoma|8140/3
C0001418|T191|SY|TCGA|NCI|Adenocarcinoma|8140/3
C0431095|T191|PT|C4712|NCI|Adenocarcinoma with Metaplasia|8140/3
C0001418|T191|PT|C2852|NCI_CDISC|ADENOCARCINOMA, MALIGNANT|8140/3
C0001418|T191|PT|C2852|NCI_CPTAC|Adenocarcinoma|8140/3
C0001418|T191|SY|C2852|NCI_CPTAC|Adenocarcinoma, NOS|8140/3
C0001418|T191|PT|10001166|NCI_CTEP-SDC|Adenocarcinoma, NOS|8140/3
C0001418|T191|PT|CDR0000046216|NCI_NCI-GLOSS|adenocarcinoma|8140/3
C0001418|T191|PT|X77nE|RCD|Adenocarcinoma|8140/3
C0431095|T191|PT|X77o2|RCD|Adenocarcinoma with metaplasia|8140/3
C0001418|T191|OP|BB52.|RCDSY|Adenocarcinoma NOS|8140/3
C0001418|T191|PT|35917007|SNOMEDCT_US|Adenocarcinoma|8140/3
C0001418|T191|SY|443961001|SNOMEDCT_US|Adenocarcinoma|8140/3
C0431095|T191|PT|253026002|SNOMEDCT_US|Adenocarcinoma with metaplasia|8140/3
C0001418|T191|SY|35917007|SNOMEDCT_US|Adenocarcinoma, no subtype|8140/3
C1531704|T191|PT|413447005|SNOMEDCT_US|Adenocarcinoma, no subtype, high grade|8140/3
C1531705|T191|PT|413448000|SNOMEDCT_US|Adenocarcinoma, no subtype, intermediate grade|8140/3
C1531706|T191|PT|413449008|SNOMEDCT_US|Adenocarcinoma, no subtype, low grade|8140/3
C0001418|T191|IS|35917007|SNOMEDCT_US|Adenocarcinoma, NOS|8140/3
C0334685|T191|PT|10146008|SNOMEDCT_US|Chief cell adenocarcinoma|8140/3
C0334685|T191|SY|10146008|SNOMEDCT_US|Chief cell carcinoma|8140/3
C0001418|T191|PT|443961001|SNOMEDCT_US|Malignant adenomatous neoplasm|8140/3
C0522636|T191|PT|103692002|SNOMEDCT_US|Meibomian adenocarcinoma|8140/3
C4518548|T191|PT|732977002|SNOMEDCT_US|Non-intestinal type adenocarcinoma|8140/3
C4518548|T191|SY|732977002|SNOMEDCT_US|Nonintestinal type adenocarcinoma|8140/3
C1270225|T191|PT|388676006|SNOMEDCT_US|Well differentiated adenocarcinoma, gastric foveolar type|8140/3
C0001418|T191|PT|1289|WHO|ADENOCARCINOMA NOS|8140/3
C0334277|T191|PT|0062844|CCPSS|ADENOCARCINOMA METASTATIC|8140/6
C0334277|T191|SY|0000029951|CHV|adenocarcinoma metastatic|8140/6
C0334277|T191|PT|0000029951|CHV|metastatic adenocarcinoma|8140/6
C0334277|T191|PT|C4124|NCI|Metastatic Adenocarcinoma|8140/6
C0334277|T191|DN|C4124|NCI_CTRP|Metastatic Adenocarcinoma|8140/6
C0334277|T191|PT|Xa98L|RCD|Metastatic adenocarcinoma|8140/6
C0334277|T191|OA|BB53.|RCDSY|Adenocarc., metastatic NOS|8140/6
C0334277|T191|OP|BB53.|RCDSY|Adenocarcinoma, metastatic, NOS|8140/6
C0334277|T191|PT|4590003|SNOMEDCT_US|Adenocarcinoma, metastatic|8140/6
C0334277|T191|IS|4590003|SNOMEDCT_US|Adenocarcinoma, metastatic, NOS|8140/6
C0334277|T191|SY|4590003|SNOMEDCT_US|Metastatic adenocarcinoma|8140/6
C0007135|T191|SY|0000002436|CHV|adenocarcinoma scirrhous|8141/3
C0007135|T191|SY|0000002436|CHV|scirrhous adenocarcinoma|8141/3
C0007135|T191|PT|0000002436|CHV|scirrhous carcinoma|8141/3
C0007135|T191|SY|271456|MEDCIN|malignant neoplasm adenocarcinoma scirrhous|8141/3
C0007135|T191|PT|271456|MEDCIN|scirrhous adenocarcinoma|8141/3
C0007135|T191|MH|D002293|MSH|Adenocarcinoma, Scirrhous|8141/3
C0007135|T191|PM|D002293|MSH|Adenocarcinomas, Scirrhous|8141/3
C0007135|T191|ET|D002293|MSH|Carcinoma, Scirrhous|8141/3
C0007135|T191|PM|D002293|MSH|Carcinomas, Scirrhous|8141/3
C0007135|T191|PM|D002293|MSH|Scirrhous Adenocarcinoma|8141/3
C0007135|T191|PM|D002293|MSH|Scirrhous Adenocarcinomas|8141/3
C0007135|T191|PM|D002293|MSH|Scirrhous Carcinoma|8141/3
C0007135|T191|PM|D002293|MSH|Scirrhous Carcinomas|8141/3
C0007135|T191|SY|C2928|NCI|Adenocarcinoma with Productive Fibrosis|8141/3
C0007135|T191|PT|C2928|NCI|Scirrhous Adenocarcinoma|8141/3
C0007135|T191|SY|C2928|NCI_CDISC|Adenocarcinoma With Productive Fibrosis|8141/3
C0007135|T191|PT|C2928|NCI_CDISC|FIBROADENOCARCINOMA, MALIGNANT|8141/3
C0007135|T191|SY|C2928|NCI_CDISC|Fibrocarcinoma|8141/3
C0007135|T191|SY|C2928|NCI_CDISC|Scirrhous Carcinoma|8141/3
C0007135|T191|AB|BB54.|RCD|Carcinoma +productive fibrosis|8141/3
C0007135|T191|SY|BB54.|RCD|Carcinoma with productive fibrosis|8141/3
C0007135|T191|PT|BB54.|RCD|Scirrhous adenocarcinoma|8141/3
C0007135|T191|SY|BB54.|RCD|Scirrhous carcinoma|8141/3
C0007135|T191|SY|4584002|SNOMEDCT_US|Carcinoma with productive fibrosis|8141/3
C0007135|T191|PT|4584002|SNOMEDCT_US|Scirrhous adenocarcinoma|8141/3
C0007135|T191|SY|4584002|SNOMEDCT_US|Scirrhous carcinoma|8141/3
C0023743|T191|SY|0000007438|CHV|leather bottle stomach|8142/3
C0023743|T191|SY|0000007438|CHV|leather-bottle stomach|8142/3
C0023743|T191|PT|0000007438|CHV|linitis plastica|8142/3
C0023743|T191|PT|MTHU090277|ICPC2ICD10ENG|leather bottle stomach|8142/3
C0023743|T191|PT|MTHU045489|ICPC2ICD10ENG|linitis plastica|8142/3
C0023743|T191|PT|10024520|MDR|Linitis plastica|8142/3
C0023743|T191|LLT|10024520|MDR|Linitis plastica|8142/3
C0023743|T191|SY|31765|MEDCIN|gastric adenocarcinoma linitis plastica|8142/3
C0023743|T191|PT|31765|MEDCIN|linitis plastica|8142/3
C0023743|T191|MH|D008039|MSH|Linitis Plastica|8142/3
C0023743|T191|PT|C3190|NCI|Linitis Plastica|8142/3
C0023743|T191|SY|XaBAo|RCD|Leather-bottle stomach|8142/3
C0023743|T191|PT|XaBAo|RCD|Linitis plastica|8142/3
C0023743|T191|PT|BB55.|RCDSY|Linitis plastica|8142/3
C0023743|T191|OAS|307594007|SNOMEDCT_US|Leather-bottle stomach|8142/3
C0023743|T191|PT|37995004|SNOMEDCT_US|Linitis plastica|8142/3
C0023743|T191|OAP|307594007|SNOMEDCT_US|Linitis plastica|8142/3
C0023743|T191|OF|307594007|SNOMEDCT_US|Linitis plastica|8142/3
C0334278|T191|SY|271457|MEDCIN|malignant neoplasm adenocarcinoma superficial spreading|8143/3
C0334278|T191|PT|271457|MEDCIN|superficial spreading adenocarcinoma|8143/3
C0334278|T191|OP|C4125|NCI|Superficial Spreading Adenocarcinoma|8143/3
C0334278|T191|PT|C4125|NCI|Superficial Spreading Adenocarcinoma|8143/3
C0334278|T191|AB|BB56.|RCD|Superficial spreading adenoca|8143/3
C0334278|T191|PT|BB56.|RCD|Superficial spreading adenocarcinoma|8143/3
C0334278|T191|PT|81446001|SNOMEDCT_US|Superficial spreading adenocarcinoma|8143/3
C0334279|T191|SY|C4126|NCI|Intestinal Type Carcinoma|8144/3
C0334279|T191|PT|C4126|NCI|Intestinal-Type Adenocarcinoma|8144/3
C0334279|T191|PT|BB57.|RCD|Adenocarcinoma - intestinal type|8144/3
C0334279|T191|AB|BB57.|RCD|Adenocarcinoma-intestinal type|8144/3
C0334279|T191|SY|BB57.|RCD|Carcinoma - intestinal type|8144/3
C0334279|T191|SY|25190001|SNOMEDCT_US|Adenocarcinoma - intestinal type|8144/3
C0334279|T191|PT|25190001|SNOMEDCT_US|Adenocarcinoma, intestinal type|8144/3
C0334279|T191|SY|25190001|SNOMEDCT_US|Carcinoma - intestinal type|8144/3
C0334279|T191|SY|25190001|SNOMEDCT_US|Carcinoma, intestinal type|8144/3
C0334280|T191|PT|MTHU014739|ICPC2ICD10ENG|carcinoma; diffuse type, unspecified site|8145/3
C0334280|T191|PT|C4127|NCI|Diffuse Type Adenocarcinoma|8145/3
C0334280|T191|SY|C4127|NCI|Diffuse Type Carcinoma|8145/3
C0334280|T191|SY|BB58.|RCD|Adenocarcinoma - diffuse type|8145/3
C0334280|T191|PT|BB58.|RCD|Carcinoma - diffuse type|8145/3
C0334280|T191|SY|24505004|SNOMEDCT_US|Adenocarcinoma - diffuse type|8145/3
C0334280|T191|SY|24505004|SNOMEDCT_US|Adenocarcinoma, diffuse type|8145/3
C0334280|T191|SY|24505004|SNOMEDCT_US|Carcinoma - diffuse type|8145/3
C0334280|T191|PT|24505004|SNOMEDCT_US|Carcinoma, diffuse type|8145/3
C0205649|T191|PT|0000020667|CHV|monomorphic adenoma|8146/0
C0205649|T191|PEP|D000236|MSH|Adenoma, Monomorphic|8146/0
C0205649|T191|PM|D000236|MSH|Adenomas, Monomorphic|8146/0
C0205649|T191|PM|D000236|MSH|Monomorphic Adenoma|8146/0
C0205649|T191|PM|D000236|MSH|Monomorphic Adenomas|8146/0
C0205649|T191|PT|C3686|NCI|Salivary Gland Monomorphic Adenoma|8146/0
C0205649|T191|PT|BB59.|RCD|Monomorphic adenoma|8146/0
C0205649|T191|PT|77653004|SNOMEDCT_US|Monomorphic adenoma|8146/0
C0205646|T191|PT|MTHU003473|ICPC2ICD10ENG|adenoma; basal cell|8147/0
C0205646|T191|PT|MTHU009781|ICPC2ICD10ENG|basal cell; adenoma|8147/0
C0205646|T191|PT|39558|MEDCIN|basal cell adenoma of salivary gland|8147/0
C0205646|T191|PEP|D000236|MSH|Adenoma, Basal Cell|8147/0
C0205646|T191|PM|D000236|MSH|Adenomas, Basal Cell|8147/0
C0205646|T191|PM|D000236|MSH|Basal Cell Adenoma|8147/0
C0205646|T191|PM|D000236|MSH|Basal Cell Adenomas|8147/0
C0205646|T191|PN|NOCODE|MTH|Adenoma, Basal Cell|8147/0
C0205646|T191|SY|C5950|NCI|Basal Cell Adenoma|8147/0
C0205646|T191|SY|C5950|NCI|Basal Cell Adenoma of Salivary Gland|8147/0
C0205646|T191|SY|C5950|NCI|Basal Cell Adenoma of the Salivary Gland|8147/0
C0205646|T191|PT|C5950|NCI|Salivary Gland Basal Cell Adenoma|8147/0
C0205646|T191|PT|BB5A.|RCD|Basal cell adenoma|8147/0
C0205646|T191|PT|27230006|SNOMEDCT_US|Basal cell adenoma|8147/0
C3697865|T191|PT|698198009|SNOMEDCT_US|Membranous basal cell adenoma|8147/0
C0205641|T191|PT|0000020662|CHV|basal cell adenocarcinoma|8147/3
C2243086|T191|LLT|10079199|MDR|Basal cell adenocarcinoma of salivary gland|8147/3
C0205641|T191|PT|271458|MEDCIN|basal cell adenocarcinoma|8147/3
C2243086|T191|PT|39576|MEDCIN|basal cell adenocarcinoma of salivary gland|8147/3
C0205641|T191|PEP|D000230|MSH|Adenocarcinoma, Basal Cell|8147/3
C0205641|T191|PM|D000230|MSH|Adenocarcinomas, Basal Cell|8147/3
C0205641|T191|PM|D000230|MSH|Basal Cell Adenocarcinoma|8147/3
C0205641|T191|PM|D000230|MSH|Basal Cell Adenocarcinomas|8147/3
C0205641|T191|PN|NOCODE|MTH|Adenocarcinoma, Basal Cell|8147/3
C2243086|T191|PN|NOCODE|MTH|basal cell adenocarcinoma of salivary gland|8147/3
C2243086|T191|SY|C3678|NCI|Basal Cell Adenocarcinoma|8147/3
C2243086|T191|SY|C3678|NCI|Basal Cell Adenocarcinoma of Salivary Gland|8147/3
C2243086|T191|SY|C3678|NCI|Basal Cell Adenocarcinoma of the Salivary Gland|8147/3
C2243086|T191|PT|C3678|NCI|Salivary Gland Basal Cell Adenocarcinoma|8147/3
C0205641|T191|PT|X77nF|RCD|Basal cell adenocarcinoma|8147/3
C0205641|T191|PT|34603009|SNOMEDCT_US|Basal cell adenocarcinoma|8147/3
C0205641|T191|OAP|189654005|SNOMEDCT_US|Basal cell adenocarcinoma|8147/3
C0205641|T191|OF|189654005|SNOMEDCT_US|Basal cell adenocarcinoma|8147/3
C1334423|T191|LA|LA26488-9|LNC|Glandular intraepithelial neoplasia, low grade|8148/0
C2348873|T191|PT|C67491|NCI|Biliary Intraepithelial Neoplasia-1|8148/0
C2348873|T191|AB|C67491|NCI|BilIN-1|8148/0
C1333457|T191|SY|C27428|NCI|Esophageal Low Grade Glandular Intraepithelial Neoplasia|8148/0
C2348873|T191|SY|C67491|NCI|Grade 1 Biliary Intraepithelial Neoplasia|8148/0
C1334423|T191|SY|C7661|NCI|Grade 1 Glandular Intraepithelial Neoplasia|8148/0
C1333861|T191|SY|C7660|NCI|Grade 2 Glandular Intraepithelial Neoplasia|8148/0
C1334423|T191|SY|C7661|NCI|Grade I Glandular Intraepithelial Neoplasia|8148/0
C1333861|T191|PT|C7660|NCI|Grade II Glandular Intraepithelial Neoplasia|8148/0
C1333457|T191|SY|C27428|NCI|Low Grade Esophageal Glandular Dysplasia|8148/0
C1333457|T191|PT|C27428|NCI|Low Grade Esophageal Glandular Intraepithelial Neoplasia|8148/0
C1334423|T191|PT|C7661|NCI|Low Grade Glandular Intraepithelial Neoplasia|8148/0
C2348873|T191|SY|C67491|NCI|Mild Biliary System Dysplasia|8148/0
C1333861|T191|SY|C7660|NCI|Moderate Glandular Dysplasia|8148/0
C1334423|T191|PT|450890000|SNOMEDCT_US|Glandular intraepithelial neoplasia, low grade|8148/0
C1334014|T191|LA|LA26489-7|LNC|Glandular intraepithelial neoplasia, high grade|8148/2
C3272438|T191|PT|C95918|NCI|Ampullary Flat Intraepithelial Neoplasia, High Grade|8148/2
C2348875|T191|PT|C67493|NCI|Biliary Intraepithelial Neoplasia-3|8148/2
C2348875|T191|AB|C67493|NCI|BilIN-3|8148/2
C1333450|T191|PT|C27425|NCI|Esophageal High Grade Intraepithelial Neoplasia|8148/2
C1333450|T191|SY|C27425|NCI|Esophageal High-Grade Dysplasia|8148/2
C1333449|T191|SY|C27429|NCI|Esophageal High-Grade Glandular Intraepithelial Neoplasia|8148/2
C1333450|T191|SY|C27425|NCI|Esophageal High-Grade Intraepithelial Neoplasia|8148/2
C2348875|T191|SY|C67493|NCI|Grade 3 Biliary Intraepithelial Neoplasia|8148/2
C1266013|T191|PT|C6877|NCI|Grade III Glandular Intraepithelial Neoplasia|8148/2
C1333449|T191|PT|C27429|NCI|High Grade Esophageal Glandular Intraepithelial Neoplasia|8148/2
C1334014|T191|PT|C7662|NCI|High Grade Glandular Intraepithelial Neoplasia|8148/2
C1333449|T191|SY|C27429|NCI|High-Grade Esophageal Glandular Dysplasia|8148/2
C1333449|T191|SY|C27429|NCI|High-Grade Esophageal Glandular Intraepithelial Neoplasia|8148/2
C1334014|T191|SY|818948002|SNOMEDCT_US|Glandular intraepithelial neoplasia grade III|8148/2
C1266013|T191|OAP|128640002|SNOMEDCT_US|Glandular intraepithelial neoplasia, grade III|8148/2
C1334014|T191|SY|818948002|SNOMEDCT_US|High grade flat intraepithelial neoplasia|8148/2
C1334014|T191|PT|818948002|SNOMEDCT_US|High grade glandular intraepithelial neoplasia|8148/2
C1335896|T191|PT|39562|MEDCIN|canalicular adenoma of salivary gland|8149/0
C1335896|T191|SY|C5979|NCI|Canalicular Adenoma of Salivary Gland|8149/0
C1335896|T191|SY|C5979|NCI|Canalicular Adenoma of the Salivary Gland|8149/0
C1335896|T191|PT|C5979|NCI|Salivary Gland Canalicular Adenoma|8149/0
C1266014|T191|PT|128641003|SNOMEDCT_US|Canalicular adenoma|8149/0
C0022134|T191|SY|0000006942|CHV|islet cell adenoma|8150/0
C0022134|T191|PT|0000006942|CHV|nesidioblastoma|8150/0
C0022134|T191|MH|D007516|MSH|Adenoma, Islet Cell|8150/0
C0022134|T191|PM|D007516|MSH|Adenomas, Islet Cell|8150/0
C0022134|T191|PM|D007516|MSH|Islet Cell Adenoma|8150/0
C0022134|T191|PM|D007516|MSH|Islet Cell Adenomas|8150/0
C0022134|T191|PN|NOCODE|MTH|Islet Cell Adenoma|8150/0
C0022134|T191|OP|C65184|NCI|Islet Cell Adenoma|8150/0
C0022134|T191|PT|C65184|NCI|Islet Cell Adenoma|8150/0
C1709454|T191|SY|C45834|NCI|Pancreatic Endocrine Microadenoma|8150/0
C1709454|T191|PT|C45834|NCI|Pancreatic Neuroendocrine Microadenoma|8150/0
C0022134|T191|PT|BB5B0|RCD|Islet cell adenoma|8150/0
C0022134|T191|OAP|189586007|SNOMEDCT_US|Islet cell adenoma|8150/0
C0022134|T191|SY|76345009|SNOMEDCT_US|Islet cell adenoma|8150/0
C0022134|T191|SY|76345009|SNOMEDCT_US|Islet cell tumor, benign|8150/0
C0022134|T191|SYGB|76345009|SNOMEDCT_US|Islet cell tumour, benign|8150/0
C0022134|T191|PT|76345009|SNOMEDCT_US|Pancreatic endocrine tumor, benign|8150/0
C0022134|T191|PTGB|76345009|SNOMEDCT_US|Pancreatic endocrine tumour, benign|8150/0
C3838828|T191|PT|703815005|SNOMEDCT_US|Pancreatic microadenoma|8150/0
C0242363|T191|SY|0000030747|CHV|endocrine pancreas tumor|8150/1
C0242363|T191|SY|0000030747|CHV|endocrine pancreas tumors|8150/1
C0242363|T191|SY|0000030747|CHV|endocrine pancreatic tumors|8150/1
C0242363|T191|SY|0000024792|CHV|islet cell adenoma|8150/1
C0242363|T191|PT|0000024792|CHV|islet cell tumor|8150/1
C0242363|T191|SY|0000024792|CHV|islet cell tumors|8150/1
C0242363|T191|SY|0000024792|CHV|islet cell tumour|8150/1
C0242363|T191|SY|0000024792|CHV|nesidioblastoma|8150/1
C0242363|T191|PT|0000030747|CHV|pancreatic endocrine tumor|8150/1
C0242363|T191|SY|NOCODE|DXP|NESIDIOBLASTOMA|8150/1
C0242363|T191|PT|HP:0030405|HPO|Pancreatic endocrine tumor|8150/1
C0242363|T191|ET|D13.7|ICD10CM|Islet cell tumor|8150/1
C0242363|T191|PT|MTHU025135|ICPC2ICD10ENG|islet cell tumor; pancreas|8150/1
C0242363|T191|PT|MTHU025134|ICPC2ICD10ENG|islet cell; tumor, pancreas|8150/1
C0242363|T191|PT|MTHU052294|ICPC2ICD10ENG|nesidioblastoma; pancreas|8150/1
C0242363|T191|PT|MTHU052293|ICPC2ICD10ENG|nesidioblastoma; unspecified site|8150/1
C0242363|T191|PT|MTHU057116|ICPC2ICD10ENG|pancreas; islet cell tumor|8150/1
C0242363|T191|PT|MTHU057144|ICPC2ICD10ENG|pancreas; nesidioblastoma|8150/1
C0242363|T191|PT|MTHU057162|ICPC2ICD10ENG|pancreas; tumor, islet cell|8150/1
C0242363|T191|PT|MTHU077050|ICPC2ICD10ENG|tumor; islet cell, pancreas|8150/1
C0242363|T191|LLT|10067518|MDR|Pancreatic neuroendocrine tumor|8150/1
C0242363|T191|MTH_PT|10067517|MDR|Pancreatic neuroendocrine tumor|8150/1
C0242363|T191|LLT|10067517|MDR|Pancreatic neuroendocrine tumour|8150/1
C0242363|T191|PT|10067517|MDR|Pancreatic neuroendocrine tumour|8150/1
C0242363|T191|PT|38714|MEDCIN|neoplasm of islets of Langerhans|8150/1
C0242363|T191|ET|D007516|MSH|Island Cell Tumor|8150/1
C0242363|T191|PM|D007516|MSH|Island Cell Tumors|8150/1
C0242363|T191|PEP|D007516|MSH|Islet Cell Tumor|8150/1
C0242363|T191|PM|D007516|MSH|Islet Cell Tumors|8150/1
C0242363|T191|ET|D007516|MSH|Nesidioblastoma|8150/1
C0242363|T191|PM|D007516|MSH|Tumor, Island Cell|8150/1
C0242363|T191|PM|D007516|MSH|Tumor, Islet Cell|8150/1
C0242363|T191|PM|D007516|MSH|Tumors, Island Cell|8150/1
C0242363|T191|PM|D007516|MSH|Tumors, Islet Cell|8150/1
C0242363|T191|PN|NOCODE|MTH|Islet Cell Tumor|8150/1
C1337011|T191|PN|NOCODE|MTH|Well Differentiated Pancreatic Endocrine Tumor|8150/1
C0242363|T191|ET|211.7|MTHICD9|Islet cell tumor|8150/1
C1337011|T191|SY|C27720|NCI|Islet Cell Tumor|8150/1
C0242363|T191|SY|C27031|NCI|Pancreatic Endocrine Neoplasm|8150/1
C1337011|T191|SY|C27720|NCI|Pancreatic NET|8150/1
C0242363|T191|PT|C27031|NCI|Pancreatic Neuroendocrine Neoplasm|8150/1
C1337011|T191|PT|C27720|NCI|Pancreatic Neuroendocrine Tumor|8150/1
C1337011|T191|AB|C27720|NCI|PanNET|8150/1
C1337011|T191|SY|C27720|NCI|Well Differentiated Pancreatic Endocrine Neoplasm|8150/1
C1337011|T191|SY|C27720|NCI|Well Differentiated Pancreatic Endocrine Tumor|8150/1
C1337011|T191|PT|C27720|NCI_CPTAC|Pancreatic Neuroendocrine Tumor|8150/1
C1337011|T191|SY|10033630|NCI_CTEP-SDC|Islet cell tumors - pancreas|8150/1
C1337011|T191|PT|10033630|NCI_CTEP-SDC|Islet cell tumors of the pancreas|8150/1
C1337011|T191|DN|C27720|NCI_CTRP|Pancreatic Neuroendocrine Tumor|8150/1
C1337011|T191|PT|CDR0000573196|NCI_NCI-GLOSS|islet cell tumor|8150/1
C0242363|T191|SY|CDR0000550688|PDQ|islet cell tumor|8150/1
C0242363|T191|SY|CDR0000550688|PDQ|pancreatic neuroendocrine neoplasm|8150/1
C0242363|T191|ET|CDR0000550688|PDQ|pancreatic neuroendocrine tumor|8150/1
C0242363|T191|PT|CDR0000550688|PDQ|pancreatic neuroendocrine tumor|8150/1
C0242363|T191|SY|BB5B0|RCD|Islet cell tumour|8150/1
C0242363|T191|SY|BB5B0|RCD|Nesidioblastoma|8150/1
C0242363|T191|SY|X40J0|RCD|Pancreatic endocrine tumour|8150/1
C0242363|T191|PT|X40J0|RCD|Tumour of endocrine pancreas|8150/1
C0242363|T191|SY|BB5B0|RCDAE|Islet cell tumor|8150/1
C0242363|T191|SY|X40J0|RCDAE|Pancreatic endocrine tumor|8150/1
C0242363|T191|PT|X40J0|RCDAE|Tumor of endocrine pancreas|8150/1
C0242363|T191|OAS|188855000|SNOMEDCT_US|Endocrine tumor of pancreas|8150/1
C0242363|T191|OAS|188855000|SNOMEDCT_US|Endocrine tumour of pancreas|8150/1
C0242363|T191|PT|399528006|SNOMEDCT_US|Islet cell neoplasm|8150/1
C0242363|T191|IS|261713004|SNOMEDCT_US|Islet cell tumor|8150/1
C0242363|T191|SY|128878003|SNOMEDCT_US|Islet cell tumor|8150/1
C0242363|T191|IS|76345009|SNOMEDCT_US|Islet cell tumor|8150/1
C0242363|T191|OAS|154609001|SNOMEDCT_US|Islet cell tumor|8150/1
C0242363|T191|OAS|269636003|SNOMEDCT_US|Islet cell tumor|8150/1
C0242363|T191|IS|261713004|SNOMEDCT_US|Islet cell tumour|8150/1
C0242363|T191|OAS|269636003|SNOMEDCT_US|Islet cell tumour|8150/1
C0242363|T191|OAS|154609001|SNOMEDCT_US|Islet cell tumour|8150/1
C0242363|T191|SYGB|128878003|SNOMEDCT_US|Islet cell tumour|8150/1
C0242363|T191|PT|126864006|SNOMEDCT_US|Neoplasm of endocrine pancreas|8150/1
C0242363|T191|SY|126864006|SNOMEDCT_US|Neoplasm of islets of Langerhans|8150/1
C0242363|T191|SY|76345009|SNOMEDCT_US|Nesidioblastoma|8150/1
C0242363|T191|SY|126864006|SNOMEDCT_US|Pancreatic endocrine tumor|8150/1
C0242363|T191|OAS|188855000|SNOMEDCT_US|Pancreatic endocrine tumor|8150/1
C0242363|T191|OAS|237596009|SNOMEDCT_US|Pancreatic endocrine tumor|8150/1
C0242363|T191|PT|128878003|SNOMEDCT_US|Pancreatic endocrine tumor|8150/1
C0242363|T191|OAS|188855000|SNOMEDCT_US|Pancreatic endocrine tumour|8150/1
C0242363|T191|OAS|237596009|SNOMEDCT_US|Pancreatic endocrine tumour|8150/1
C0242363|T191|PTGB|128878003|SNOMEDCT_US|Pancreatic endocrine tumour|8150/1
C0242363|T191|SYGB|126864006|SNOMEDCT_US|Pancreatic endocrine tumour|8150/1
C0242363|T191|SY|126864006|SNOMEDCT_US|Tumor of endocrine pancreas|8150/1
C0242363|T191|OAP|237596009|SNOMEDCT_US|Tumor of endocrine pancreas|8150/1
C0242363|T191|SYGB|126864006|SNOMEDCT_US|Tumour of endocrine pancreas|8150/1
C0242363|T191|OAP|237596009|SNOMEDCT_US|Tumour of endocrine pancreas|8150/1
C1328479|T191|PT|0000021022|CHV|islet cell carcinoma|8150/3
C1328479|T191|ET|C25.4|ICD10CM|Malignant neoplasm of islets of Langerhans|8150/3
C1328479|T191|AB|157.4|ICD9CM|Mal neo islet langerhans|8150/3
C1328479|T191|PT|157.4|ICD9CM|Malignant neoplasm of islets of langerhans|8150/3
C1328479|T191|PT|MTHU014747|ICPC2ICD10ENG|carcinoma; islet cell, pancreas|8150/3
C1328479|T191|PT|MTHU014746|ICPC2ICD10ENG|carcinoma; islet cell, unspecified site|8150/3
C1328479|T191|PT|MTHU025130|ICPC2ICD10ENG|islet cell; carcinoma, pancreas|8150/3
C1328479|T191|PT|MTHU025129|ICPC2ICD10ENG|islet cell; carcinoma, unspecified site|8150/3
C1328479|T191|PT|MTHU057103|ICPC2ICD10ENG|pancreas; carcinoma, islet cell|8150/3
C1328479|T191|PT|MTHU057115|ICPC2ICD10ENG|pancreas; islet cell carcinoma|8150/3
C1328479|T191|LLT|10025997|MDR|Malignant neoplasm of islets of Langerhans|8150/3
C1328479|T191|PT|10025997|MDR|Malignant neoplasm of islets of Langerhans|8150/3
C1328479|T191|LLT|10026664|MDR|Malignant pancreatic islet neoplasm|8150/3
C1328479|T191|LLT|10062715|MDR|Pancreatic islet cell carcinoma|8150/3
C1328479|T191|LLT|10033630|MDR|Pancreatic islet cell neoplasm malignant NOS|8150/3
C1328479|T191|PT|350413|MEDCIN|Carcinoma of endocrine pancreas|8150/3
C1328479|T191|PT|271423|MEDCIN|islet cell carcinoma|8150/3
C1328479|T191|PT|218345|MEDCIN|islet cell carcinoma of pancreas|8150/3
C1328479|T191|SY|351055|MEDCIN|malignant neoplasm endocrine glands islets of langerhans|8150/3
C1328479|T191|PT|351055|MEDCIN|malignant neoplasm of Islets of Langerhans|8150/3
C1328479|T191|SY|350413|MEDCIN|pancreatic neoplasm malignant carcinoma endocrine pancreas|8150/3
C1328479|T191|ET|469|MEDLINEPLUS|Islet Cell Carcinoma|8150/3
C1328479|T191|MH|D018273|MSH|Carcinoma, Islet Cell|8150/3
C1328479|T191|PM|D018273|MSH|Carcinomas, Islet Cell|8150/3
C1328479|T191|PM|D018273|MSH|Islet Cell Carcinoma|8150/3
C1328479|T191|PM|D018273|MSH|Islet Cell Carcinomas|8150/3
C1328479|T191|ET|D018273|MSH|Islet Cell Tumor, Malignant|8150/3
C1334977|T191|NM|C536126|MSH|Non functioning pancreatic endocrine tumor|8150/3
C1334977|T191|CE|C536126|MSH|Non-functioning endocrine pancreatic tumors|8150/3
C1328479|T191|PN|NOCODE|MTH|Pancreatic Endocrine Carcinoma|8150/3
C1328479|T191|ET|157.4|MTHICD9|Malignant neoplasm of Islets of Langerhans, any part of pancreas|8150/3
C1328479|T191|SY|C3770|NCI|High Grade Pancreatic Neuroendocrine Carcinoma|8150/3
C1328479|T191|SY|C3770|NCI|High-Grade Pancreatic Neuroendocrine Carcinoma|8150/3
C1334977|T191|SY|C45837|NCI|Inactive Pancreatic Endocrine Tumor|8150/3
C1328479|T191|SY|C3770|NCI|Islet Cell Carcinoma|8150/3
C1334977|T191|SY|C45837|NCI|Non-Functional Pancreatic Neuroendocrine Tumor|8150/3
C1334977|T191|SY|C45837|NCI|Non-Functioning Pancreatic Endocrine Tumor|8150/3
C1334977|T191|SY|C45837|NCI|Non-Functioning Pancreatic NET|8150/3
C1334977|T191|PT|C45837|NCI|Non-Functioning Pancreatic Neuroendocrine Tumor|8150/3
C1334977|T191|SY|C45837|NCI|Non-Functioning Well Differentiated Pancreatic Endocrine Tumor|8150/3
C1334977|T191|SY|C45837|NCI|Non-Syndromic Pancreatic NET|8150/3
C1334977|T191|SY|C45837|NCI|Non-Syndromic Pancreatic Neuroendocrine Tumor|8150/3
C1334977|T191|SY|C45837|NCI|Nonfunctional Pancreatic NET|8150/3
C1334977|T191|SY|C45837|NCI|Nonfunctional Pancreatic Neuroendocrine Tumor|8150/3
C1334977|T191|SY|C45837|NCI|Nonfunctioning Pancreatic Neuroendocrine Tumor|8150/3
C1334977|T191|SY|C45837|NCI|Nonsyndromic Pancreatic Endocrine Tumor|8150/3
C1334977|T191|SY|C45837|NCI|Nonsyndromic Pancreatic Neuroendocrine Tumor|8150/3
C1328479|T191|SY|C3770|NCI|Pancreatic Endocrine Carcinoma|8150/3
C1328479|T191|SY|C3770|NCI|Pancreatic NEC|8150/3
C1328479|T191|SY|C3770|NCI|Pancreatic NEC G3|8150/3
C1328479|T191|PT|C3770|NCI|Pancreatic Neuroendocrine Carcinoma|8150/3
C1328479|T191|AB|C3770|NCI|PanNEC|8150/3
C1328479|T191|SY|C3770|NCI|Poorly Differentiated Neuroendocrine Neoplasm|8150/3
C1328479|T191|SY|C3770|NCI|Poorly Differentiated Pancreatic Endocrine Carcinoma|8150/3
C1328479|T191|PT|C3770|NCI_CDISC|CARCINOMA, ISLET CELL, MALIGNANT|8150/3
C1328479|T191|SY|C3770|NCI_CDISC|Islet Cell Cancer|8150/3
C1328479|T191|SY|C3770|NCI_CDISC|Islet Cell Carcinoma|8150/3
C1328479|T191|SY|C3770|NCI_CDISC|Malignant Islet Cell Tumor|8150/3
C1328479|T191|SY|C3770|NCI_CDISC|Malignant Pancreatic Endocrine Tumor|8150/3
C1328479|T191|SY|C3770|NCI_CDISC|Pancreatic Neuroendocrine Carcinoma|8150/3
C1328479|T191|PT|C3770|NCI_CPTAC|Pancreatic Neuroendocrine Carcinoma|8150/3
C1334977|T191|DN|C45837|NCI_CTRP|Non-Functioning Pancreatic Neuroendocrine Tumor|8150/3
C1328479|T191|DN|C3770|NCI_CTRP|Pancreatic Neuroendocrine Cancer|8150/3
C1328479|T191|PT|CDR0000046343|NCI_NCI-GLOSS|islet cell cancer|8150/3
C1328479|T191|PT|CDR0000530385|NCI_NCI-GLOSS|pancreatic endocrine cancer|8150/3
C1328479|T191|SY|CDR0000043353|PDQ|cancer of the endocrine pancreas|8150/3
C1328479|T191|SY|CDR0000043353|PDQ|carcinoma of the endocrine pancreas|8150/3
C1328479|T191|SY|CDR0000043353|PDQ|endocrine pancreatic cancer|8150/3
C1328479|T191|PSC|CDR0000043353|PDQ|islet cell carcinoma|8150/3
C1328479|T191|SY|CDR0000043353|PDQ|pancreatic endocrine cancer|8150/3
C1328479|T191|SY|CDR0000043353|PDQ|pancreatic endocrine carcinoma|8150/3
C1328479|T191|OA|X78Pg|RCD|Carcinoma endocrine pancreas|8150/3
C1328479|T191|OP|X78Pg|RCD|Carcinoma of endocrine pancreas|8150/3
C1328479|T191|IS|X78Pg|RCD|Endocrine pancreatic carcinoma|8150/3
C1328479|T191|SY|BB5B1|RCD|Islet cell adenocarcinoma|8150/3
C1328479|T191|PT|BB5B1|RCD|Islet cell carcinoma|8150/3
C1328479|T191|OA|B174.|RCD|Malig neop Islets Langerhans|8150/3
C1328479|T191|OA|B174.|RCD|Malign tumour Islet Langerhans|8150/3
C1328479|T191|IS|B174.|RCD|Malignant Islet cell tumour|8150/3
C1328479|T191|IS|B174.|RCD|Malignant neoplasm of Islets of Langerhans|8150/3
C1328479|T191|OP|B174.|RCD|Malignant tumour of Islets of Langerhans|8150/3
C1328479|T191|OA|B174.|RCDAE|Malign tumor Islet Langerhans|8150/3
C1328479|T191|IS|B174.|RCDAE|Malignant Islet cell tumor|8150/3
C1328479|T191|OP|B174.|RCDAE|Malignant tumor of Islets of Langerhans|8150/3
C1328479|T191|PT|254612002|SNOMEDCT_US|Carcinoma of endocrine pancreas|8150/3
C1328479|T191|SY|254612002|SNOMEDCT_US|Endocrine pancreatic carcinoma|8150/3
C1328479|T191|SY|60346004|SNOMEDCT_US|Islet cell adenocarcinoma|8150/3
C1328479|T191|SY|60346004|SNOMEDCT_US|Islet cell carcinoma|8150/3
C1328479|T191|SY|187794005|SNOMEDCT_US|Malignant Islet cell tumor|8150/3
C1328479|T191|SYGB|187794005|SNOMEDCT_US|Malignant Islet cell tumour|8150/3
C1328479|T191|IS|93843007|SNOMEDCT_US|Malignant neoplasm of islets of Langerhans|8150/3
C1328479|T191|SY|187794005|SNOMEDCT_US|Malignant neoplasm of Islets of Langerhans|8150/3
C1328479|T191|PT|187794005|SNOMEDCT_US|Malignant tumor of Islets of Langerhans|8150/3
C1328479|T191|PTGB|187794005|SNOMEDCT_US|Malignant tumour of Islets of Langerhans|8150/3
C1328479|T191|PT|60346004|SNOMEDCT_US|Pancreatic endocrine tumor, malignant|8150/3
C3839703|T191|PT|703816006|SNOMEDCT_US|Pancreatic endocrine tumor, nonfunctioning|8150/3
C1328479|T191|PTGB|60346004|SNOMEDCT_US|Pancreatic endocrine tumour, malignant|8150/3
C3839703|T191|PTGB|703816006|SNOMEDCT_US|Pancreatic endocrine tumour, nonfunctioning|8150/3
C1276147|T191|PT|261713004|SNOMEDCT_US|Metastatic islet cell carcinoma|8150/6
C0021670|T191|PT|0048177|CCPSS|INSULINOMA|8151/0
C0021670|T191|PT|0000006789|CHV|insulinoma|8151/0
C0021670|T191|SY|0000006789|CHV|insulinomas|8151/0
C0021670|T191|SY|0000006789|CHV|insuloma|8151/0
C0021670|T191|SY|0000006789|CHV|pancreatic insulinoma|8151/0
C0021670|T191|ET|2014-4965|CSP|insulinoma|8151/0
C0021670|T191|SY|NOCODE|DXP|INSULINOMA|8151/0
C0021670|T191|SY|NOCODE|DXP|INSULOMA|8151/0
C0021670|T191|DI|U001399|DXP|PANCREAS, ISLET-CELL TUMOR, INSULIN-PRODUCING|8151/0
C0021670|T191|PT|HP:0012197|HPO|Insulinoma|8151/0
C0021670|T191|SY|HP:0012197|HPO|Pancreatic insulinoma|8151/0
C0021670|T191|PT|MTHU003478|ICPC2ICD10ENG|adenoma; beta-cell, pancreas|8151/0
C0021670|T191|PT|MTHU010446|ICPC2ICD10ENG|beta-cell; adenoma, pancreas|8151/0
C0021670|T191|PT|MTHU010450|ICPC2ICD10ENG|beta-cell; tumor, pancreas|8151/0
C0021670|T191|PT|MTHU010449|ICPC2ICD10ENG|beta-cell; tumor, unspecified site|8151/0
C0021670|T191|PT|MTHU039746|ICPC2ICD10ENG|insulinoma; pancreas|8151/0
C0021670|T191|PT|MTHU039745|ICPC2ICD10ENG|insulinoma; unspecified site|8151/0
C0021670|T191|PT|MTHU057085|ICPC2ICD10ENG|pancreas; adenoma, beta-cell|8151/0
C0021670|T191|PT|MTHU057099|ICPC2ICD10ENG|pancreas; beta-cell tumor|8151/0
C0021670|T191|PT|MTHU057132|ICPC2ICD10ENG|pancreas; insulinoma|8151/0
C0021670|T191|PT|MTHU057160|ICPC2ICD10ENG|pancreas; tumor, beta-cell|8151/0
C0021670|T191|PT|MTHU077025|ICPC2ICD10ENG|tumor; beta-cell, pancreas|8151/0
C0021670|T191|PT|MTHU077024|ICPC2ICD10ENG|tumor; beta-cell, unspecified site|8151/0
C0021670|T191|PTN|T73009|ICPC2P|insulinoma|8151/0
C0021670|T191|PT|T73009|ICPC2P|Insulinoma|8151/0
C0021670|T191|LLT|10022498|MDR|Insulinoma|8151/0
C0021670|T191|PT|10022498|MDR|Insulinoma|8151/0
C0021670|T191|PM|D007340|MSH|Adenoma, beta Cell|8151/0
C0021670|T191|ET|D007340|MSH|Adenoma, beta-Cell|8151/0
C0021670|T191|PM|D007340|MSH|Adenomas, beta-Cell|8151/0
C0021670|T191|PM|D007340|MSH|beta Cell Tumor|8151/0
C0021670|T191|PM|D007340|MSH|beta-Cell Adenoma|8151/0
C0021670|T191|PM|D007340|MSH|beta-Cell Adenomas|8151/0
C0021670|T191|ET|D007340|MSH|beta-Cell Tumor|8151/0
C0021670|T191|PM|D007340|MSH|beta-Cell Tumors|8151/0
C0021670|T191|MH|D007340|MSH|Insulinoma|8151/0
C0021670|T191|PM|D007340|MSH|Insulinomas|8151/0
C0021670|T191|ET|D007340|MSH|Insuloma|8151/0
C0021670|T191|PM|D007340|MSH|Insulomas|8151/0
C0021670|T191|PM|D007340|MSH|Tumor, beta-Cell|8151/0
C0021670|T191|PM|D007340|MSH|Tumors, beta-Cell|8151/0
C0021670|T191|PN|NOCODE|MTH|insulinoma|8151/0
C0021670|T191|SY|C3140|NCI|Beta Cell Tumor|8151/0
C0021670|T191|SY|C3140|NCI|Beta Cell Tumor of Pancreas|8151/0
C0021670|T191|SY|C3140|NCI|Beta Cell Tumor of the Pancreas|8151/0
C0021670|T191|SY|C3140|NCI|Insulin-Producing Islet Cell Tumor|8151/0
C0021670|T191|SY|C3140|NCI|Insulin-Producing Tumor of Islet Cells|8151/0
C0021670|T191|SY|C3140|NCI|Insulin-Producing Tumor of the Islet Cells|8151/0
C0021670|T191|SY|C95598|NCI|Insulinoma|8151/0
C0021670|T191|SY|C3140|NCI|Pancreatic Beta Cell Tumor|8151/0
C0021670|T191|SY|C3140|NCI|Pancreatic Insulin Producing Neoplasm|8151/0
C0021670|T191|SY|C3140|NCI|Pancreatic Insulin Producing NET|8151/0
C0021670|T191|SY|C3140|NCI|Pancreatic Insulin Producing Tumor|8151/0
C0021670|T191|PT|C3140|NCI|Pancreatic Insulin-Producing Neuroendocrine Tumor|8151/0
C0021670|T191|PT|C95598|NCI|Pancreatic Insulinoma|8151/0
C0021670|T191|DN|C3140|NCI_CTRP|Pancreatic Insulin-Producing Neuroendocrine Tumor|8151/0
C0021670|T191|DN|C95598|NCI_CTRP|Pancreatic Insulinoma|8151/0
C0021670|T191|PT|CDR0000657854|NCI_NCI-GLOSS|beta cell neoplasm|8151/0
C0021670|T191|PT|CDR0000657855|NCI_NCI-GLOSS|beta cell tumor of the pancreas|8151/0
C0021670|T191|PT|CDR0000657853|NCI_NCI-GLOSS|insulinoma|8151/0
C0021670|T191|PT|CDR0000657856|NCI_NCI-GLOSS|pancreatic insulin-producing tumor|8151/0
C0021670|T191|PT|C95598|NCI_NICHD|Insulinoma|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Neoplasm|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Neoplasm of Pancreas|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Neoplasm of the Pancreas|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Tumor|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Tumor of Pancreas|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Tumor of the Pancreas|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Islet Cell Neoplasm|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Islet Cell Tumor|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Neoplasm of Islet Cells|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Neoplasm of the Islet Cells|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Tumor of Islet Cells|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Tumor of the Islet Cells|8151/0
C0021670|T191|PSC|CDR0000038792|PDQ|insulinoma|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Insulinoma|8151/0
C0021670|T191|SY|CDR0000038792|PDQ|islet cell insulinoma|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Pancreatic Beta Cell Tumor|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Pancreatic Insulin Producing Neoplasm|8151/0
C0021670|T191|SY|CDR0000040018|PDQ|Pancreatic Insulin Producing Tumor|8151/0
C0021670|T191|SY|CDR0000038792|PDQ|pancreatic insulinoma|8151/0
C0021670|T191|PT|R0121652|QMR|INSULINOMA|8151/0
C0021670|T191|SY|Xa98M|RCD|Beta cell adenoma|8151/0
C0021670|T191|PT|Xa98M|RCD|Insulinoma|8151/0
C0021670|T191|PT|BB5B2|RCDSY|Insulinoma NOS|8151/0
C5229670|T191|SY|788388009|SNOMEDCT_US|Benign beta cell adenoma|8151/0
C5229670|T191|PT|788388009|SNOMEDCT_US|Benign insulinoma|8151/0
C5229670|T191|PT|788390005|SNOMEDCT_US|Benign insulinoma|8151/0
C0021670|T191|OAS|25324008|SNOMEDCT_US|Beta cell adenoma|8151/0
C0021670|T191|OAS|302822000|SNOMEDCT_US|Beta cell adenoma|8151/0
C0021670|T191|OAP|25324008|SNOMEDCT_US|Insulinoma|8151/0
C0021670|T191|OAP|302822000|SNOMEDCT_US|Insulinoma|8151/0
C0021670|T191|IS|25324008|SNOMEDCT_US|Insulinoma, NOS|8151/0
C0021670|T191|PT|0048177|CCPSS|INSULINOMA|8151/1
C0021670|T191|PT|0000006789|CHV|insulinoma|8151/1
C0021670|T191|SY|0000006789|CHV|insulinomas|8151/1
C0021670|T191|SY|0000006789|CHV|insuloma|8151/1
C0021670|T191|SY|0000006789|CHV|pancreatic insulinoma|8151/1
C0021670|T191|ET|2014-4965|CSP|insulinoma|8151/1
C0021670|T191|SY|NOCODE|DXP|INSULINOMA|8151/1
C0021670|T191|SY|NOCODE|DXP|INSULOMA|8151/1
C0021670|T191|DI|U001399|DXP|PANCREAS, ISLET-CELL TUMOR, INSULIN-PRODUCING|8151/1
C0021670|T191|PT|HP:0012197|HPO|Insulinoma|8151/1
C0021670|T191|SY|HP:0012197|HPO|Pancreatic insulinoma|8151/1
C0021670|T191|PT|MTHU003478|ICPC2ICD10ENG|adenoma; beta-cell, pancreas|8151/1
C0021670|T191|PT|MTHU010446|ICPC2ICD10ENG|beta-cell; adenoma, pancreas|8151/1
C0021670|T191|PT|MTHU010450|ICPC2ICD10ENG|beta-cell; tumor, pancreas|8151/1
C0021670|T191|PT|MTHU010449|ICPC2ICD10ENG|beta-cell; tumor, unspecified site|8151/1
C0021670|T191|PT|MTHU039746|ICPC2ICD10ENG|insulinoma; pancreas|8151/1
C0021670|T191|PT|MTHU039745|ICPC2ICD10ENG|insulinoma; unspecified site|8151/1
C0021670|T191|PT|MTHU057085|ICPC2ICD10ENG|pancreas; adenoma, beta-cell|8151/1
C0021670|T191|PT|MTHU057099|ICPC2ICD10ENG|pancreas; beta-cell tumor|8151/1
C0021670|T191|PT|MTHU057132|ICPC2ICD10ENG|pancreas; insulinoma|8151/1
C0021670|T191|PT|MTHU057160|ICPC2ICD10ENG|pancreas; tumor, beta-cell|8151/1
C0021670|T191|PT|MTHU077025|ICPC2ICD10ENG|tumor; beta-cell, pancreas|8151/1
C0021670|T191|PT|MTHU077024|ICPC2ICD10ENG|tumor; beta-cell, unspecified site|8151/1
C0021670|T191|PTN|T73009|ICPC2P|insulinoma|8151/1
C0021670|T191|PT|T73009|ICPC2P|Insulinoma|8151/1
C0021670|T191|LLT|10022498|MDR|Insulinoma|8151/1
C0021670|T191|PT|10022498|MDR|Insulinoma|8151/1
C0021670|T191|PM|D007340|MSH|Adenoma, beta Cell|8151/1
C0021670|T191|ET|D007340|MSH|Adenoma, beta-Cell|8151/1
C0021670|T191|PM|D007340|MSH|Adenomas, beta-Cell|8151/1
C0021670|T191|PM|D007340|MSH|beta Cell Tumor|8151/1
C0021670|T191|PM|D007340|MSH|beta-Cell Adenoma|8151/1
C0021670|T191|PM|D007340|MSH|beta-Cell Adenomas|8151/1
C0021670|T191|ET|D007340|MSH|beta-Cell Tumor|8151/1
C0021670|T191|PM|D007340|MSH|beta-Cell Tumors|8151/1
C0021670|T191|MH|D007340|MSH|Insulinoma|8151/1
C0021670|T191|PM|D007340|MSH|Insulinomas|8151/1
C0021670|T191|ET|D007340|MSH|Insuloma|8151/1
C0021670|T191|PM|D007340|MSH|Insulomas|8151/1
C0021670|T191|PM|D007340|MSH|Tumor, beta-Cell|8151/1
C0021670|T191|PM|D007340|MSH|Tumors, beta-Cell|8151/1
C0021670|T191|PN|NOCODE|MTH|insulinoma|8151/1
C0021670|T191|SY|C3140|NCI|Beta Cell Tumor|8151/1
C0021670|T191|SY|C3140|NCI|Beta Cell Tumor of Pancreas|8151/1
C0021670|T191|SY|C3140|NCI|Beta Cell Tumor of the Pancreas|8151/1
C0021670|T191|SY|C3140|NCI|Insulin-Producing Islet Cell Tumor|8151/1
C0021670|T191|SY|C3140|NCI|Insulin-Producing Tumor of Islet Cells|8151/1
C0021670|T191|SY|C3140|NCI|Insulin-Producing Tumor of the Islet Cells|8151/1
C0021670|T191|SY|C95598|NCI|Insulinoma|8151/1
C0021670|T191|SY|C3140|NCI|Pancreatic Beta Cell Tumor|8151/1
C0021670|T191|SY|C3140|NCI|Pancreatic Insulin Producing Neoplasm|8151/1
C0021670|T191|SY|C3140|NCI|Pancreatic Insulin Producing NET|8151/1
C0021670|T191|SY|C3140|NCI|Pancreatic Insulin Producing Tumor|8151/1
C0021670|T191|PT|C3140|NCI|Pancreatic Insulin-Producing Neuroendocrine Tumor|8151/1
C0021670|T191|PT|C95598|NCI|Pancreatic Insulinoma|8151/1
C0021670|T191|DN|C3140|NCI_CTRP|Pancreatic Insulin-Producing Neuroendocrine Tumor|8151/1
C0021670|T191|DN|C95598|NCI_CTRP|Pancreatic Insulinoma|8151/1
C0021670|T191|PT|CDR0000657854|NCI_NCI-GLOSS|beta cell neoplasm|8151/1
C0021670|T191|PT|CDR0000657855|NCI_NCI-GLOSS|beta cell tumor of the pancreas|8151/1
C0021670|T191|PT|CDR0000657853|NCI_NCI-GLOSS|insulinoma|8151/1
C0021670|T191|PT|CDR0000657856|NCI_NCI-GLOSS|pancreatic insulin-producing tumor|8151/1
C0021670|T191|PT|C95598|NCI_NICHD|Insulinoma|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Neoplasm|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Neoplasm of Pancreas|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Neoplasm of the Pancreas|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Tumor|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Tumor of Pancreas|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Beta Cell Tumor of the Pancreas|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Islet Cell Neoplasm|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Islet Cell Tumor|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Neoplasm of Islet Cells|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Neoplasm of the Islet Cells|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Tumor of Islet Cells|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Insulin-Producing Tumor of the Islet Cells|8151/1
C0021670|T191|PSC|CDR0000038792|PDQ|insulinoma|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Insulinoma|8151/1
C0021670|T191|SY|CDR0000038792|PDQ|islet cell insulinoma|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Pancreatic Beta Cell Tumor|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Pancreatic Insulin Producing Neoplasm|8151/1
C0021670|T191|SY|CDR0000040018|PDQ|Pancreatic Insulin Producing Tumor|8151/1
C0021670|T191|SY|CDR0000038792|PDQ|pancreatic insulinoma|8151/1
C0021670|T191|PT|R0121652|QMR|INSULINOMA|8151/1
C0021670|T191|SY|Xa98M|RCD|Beta cell adenoma|8151/1
C0021670|T191|PT|Xa98M|RCD|Insulinoma|8151/1
C0021670|T191|PT|BB5B2|RCDSY|Insulinoma NOS|8151/1
C0021670|T191|OAS|25324008|SNOMEDCT_US|Beta cell adenoma|8151/1
C0021670|T191|OAS|302822000|SNOMEDCT_US|Beta cell adenoma|8151/1
C0021670|T191|OAP|302822000|SNOMEDCT_US|Insulinoma|8151/1
C0021670|T191|OAP|25324008|SNOMEDCT_US|Insulinoma|8151/1
C0021670|T191|IS|25324008|SNOMEDCT_US|Insulinoma, NOS|8151/1
C0334281|T191|PN|NOCODE|MTH|Insulinoma, malignant|8151/3
C4721412|T191|PN|NOCODE|MTH|Malignant Pancreatic Insulinoma|8151/3
C4721412|T191|SY|C65186|NCI|Malignant Insulinoma|8151/3
C4721412|T191|PT|C65186|NCI|Malignant Pancreatic Insulinoma|8151/3
C4721412|T191|SY|C65186|NCI|Pancreatic Beta Islet Cell Carcinoma|8151/3
C4721412|T191|SY|C65186|NCI|Pancreatic Insulin Producing Carcinoma|8151/3
C4721412|T191|DN|C65186|NCI_CTRP|Malignant Pancreatic Insulinoma|8151/3
C4721412|T191|SY|CDR0000040020|PDQ|beta islet cell carcinoma, pancreatic|8151/3
C4721412|T191|SY|CDR0000040020|PDQ|carcinoma, pancreatic beta islet cell|8151/3
C4721412|T191|SY|CDR0000040020|PDQ|insulin producing carcinoma|8151/3
C4721412|T191|SY|CDR0000040020|PDQ|insulin secreting carcinoma|8151/3
C4721412|T191|SY|CDR0000040020|PDQ|islet cell, beta, pancreatic carcinoma|8151/3
C4721412|T191|SY|CDR0000040020|PDQ|Malignant Insulinoma|8151/3
C4721412|T191|PT|CDR0000040020|PDQ|pancreatic beta islet cell carcinoma|8151/3
C4721412|T191|SY|CDR0000040020|PDQ|Pancreatic Insulin Producing Carcinoma|8151/3
C0334281|T191|SY|BB5B3|RCD|Malignant beta cell tumour|8151/3
C0334281|T191|PT|BB5B3|RCD|Malignant insulinoma|8151/3
C0334281|T191|SY|BB5B3|RCDAE|Malignant beta cell tumor|8151/3
C0334281|T191|SY|20955008|SNOMEDCT_US|Beta cell tumor, malignant|8151/3
C0334281|T191|SYGB|20955008|SNOMEDCT_US|Beta cell tumour, malignant|8151/3
C0334281|T191|PT|20955008|SNOMEDCT_US|Insulinoma, malignant|8151/3
C0334281|T191|SY|20955008|SNOMEDCT_US|Malignant beta cell tumor|8151/3
C0334281|T191|SYGB|20955008|SNOMEDCT_US|Malignant beta cell tumour|8151/3
C0334281|T191|PT|713189001|SNOMEDCT_US|Malignant insulinoma|8151/3
C0334281|T191|SY|20955008|SNOMEDCT_US|Malignant insulinoma|8151/3
C0017689|T191|PT|0000005553|CHV|glucagonoma|8152/1
C0017689|T191|SY|0000005553|CHV|glucagonomas|8152/1
C0017689|T191|SY|NOCODE|DXP|GLUCAGONOMA|8152/1
C0017689|T191|DI|U001398|DXP|PANCREAS, ISLET-CELL TUMOR, GLUCAGON-PRODUCING|8152/1
C0017689|T191|PT|HP:0030404|HPO|Glucagonoma|8152/1
C0017689|T191|PT|MTHU004942|ICPC2ICD10ENG|alpha cell; tumor, pancreas|8152/1
C0017689|T191|PT|MTHU004941|ICPC2ICD10ENG|alpha cell; tumor, unspecified site|8152/1
C0017689|T191|PT|MTHU032353|ICPC2ICD10ENG|glucagonoma; pancreas|8152/1
C0017689|T191|PT|MTHU032352|ICPC2ICD10ENG|glucagonoma; unspecified site|8152/1
C0017689|T191|PT|MTHU057092|ICPC2ICD10ENG|pancreas; alpha cell tumor|8152/1
C0017689|T191|PT|MTHU057124|ICPC2ICD10ENG|pancreas; glucagonoma|8152/1
C0017689|T191|PT|MTHU057158|ICPC2ICD10ENG|pancreas; tumor, alpha cell|8152/1
C0017689|T191|PT|MTHU077014|ICPC2ICD10ENG|tumor; alpha cell, pancreas|8152/1
C0017689|T191|PT|MTHU077013|ICPC2ICD10ENG|tumor; alpha cell, unspecified site|8152/1
C0017689|T191|PT|U001985|LCH|Glucagonoma|8152/1
C0017689|T191|PT|sh85055354|LCH_NW|Glucagonoma|8152/1
C0017689|T191|PT|10018404|MDR|Glucagonoma|8152/1
C0017689|T191|LLT|10018404|MDR|Glucagonoma|8152/1
C0017689|T191|PT|37609|MEDCIN|glucagonoma|8152/1
C0017689|T191|PT|31633|MEDCIN|glucagonoma of pancreas|8152/1
C0017689|T191|SY|31633|MEDCIN|pancreatic glucagonoma|8152/1
C0017689|T191|PM|D005935|MSH|Adenoma, alpha Cell|8152/1
C0017689|T191|ET|D005935|MSH|Adenoma, alpha-Cell|8152/1
C0017689|T191|PM|D005935|MSH|Adenomas, alpha-Cell|8152/1
C0017689|T191|PM|D005935|MSH|alpha Cell Tumor|8152/1
C0017689|T191|PM|D005935|MSH|alpha-Cell Adenoma|8152/1
C0017689|T191|PM|D005935|MSH|alpha-Cell Adenomas|8152/1
C0017689|T191|ET|D005935|MSH|alpha-Cell Tumor|8152/1
C0017689|T191|PM|D005935|MSH|alpha-Cell Tumors|8152/1
C0017689|T191|MH|D005935|MSH|Glucagonoma|8152/1
C0017689|T191|ET|D005935|MSH|Glucagonoma Syndrome|8152/1
C0017689|T191|PM|D005935|MSH|Glucagonoma Syndromes|8152/1
C0017689|T191|PM|D005935|MSH|Glucagonomas|8152/1
C0017689|T191|PM|D005935|MSH|Syndrome, Glucagonoma|8152/1
C0017689|T191|PM|D005935|MSH|Syndromes, Glucagonoma|8152/1
C0017689|T191|PM|D005935|MSH|Tumor, alpha-Cell|8152/1
C0017689|T191|PM|D005935|MSH|Tumors, alpha-Cell|8152/1
C0017689|T191|PN|NOCODE|MTH|Glucagonoma|8152/1
C0017689|T191|SY|C3062|NCI|Alpha Cell Tumor|8152/1
C0017689|T191|SY|C3062|NCI|Alpha Cell Tumor of Pancreas|8152/1
C0017689|T191|SY|C3062|NCI|Alpha Cell Tumor of the Pancreas|8152/1
C1266016|T191|OP|C66925|NCI|Enteroglucagonoma|8152/1
C1266016|T191|PT|C66925|NCI|Enteroglucagonoma|8152/1
C0017689|T191|SY|C3062|NCI|Glucagon-Producing Islet Cell Tumor|8152/1
C0017689|T191|SY|C3062|NCI|Glucagon-Producing Tumor of Islet Cells|8152/1
C0017689|T191|SY|C3062|NCI|Glucagon-Producing Tumor of the Islet Cells|8152/1
C0017689|T191|SY|C95597|NCI|Glucagonoma|8152/1
C3274140|T191|SY|C27448|NCI|L-Cell Glucagon-Like Peptide-Producing NET|8152/1
C3274140|T191|PT|C27448|NCI|L-Cell Glucagon-Like Peptide-Producing Neuroendocrine Tumor|8152/1
C0017689|T191|SY|C3062|NCI|Pancreatic Alpha Cell Tumor|8152/1
C0017689|T191|SY|C3062|NCI|Pancreatic Glucagon Producing NET|8152/1
C0017689|T191|SY|C3062|NCI|Pancreatic Glucagon Producing Neuroendocrine Tumor|8152/1
C0017689|T191|SY|C3062|NCI|Pancreatic Glucagon Producing Tumor|8152/1
C0017689|T191|PT|C3062|NCI|Pancreatic Glucagon-Producing Neuroendocrine Tumor|8152/1
C0017689|T191|PT|C95597|NCI|Pancreatic Glucagonoma|8152/1
C1882278|T191|OP|C67453|NCI|Pancreatic Polypeptide Neoplasm|8152/1
C1882278|T191|OP|C67453|NCI|Pancreatic Polypeptide Tumor|8152/1
C1882278|T191|PT|C67453|NCI|Pancreatic Polypeptide Tumor|8152/1
C1882278|T191|AB|C67453|NCI|PPoma|8152/1
C0017689|T191|DN|C95597|NCI_CTRP|Pancreatic Glucagonoma|8152/1
C1882278|T191|DN|C67453|NCI_CTRP|Pancreatic Polypeptide Tumor|8152/1
C0017689|T191|PT|CDR0000044280|NCI_NCI-GLOSS|glucagonoma|8152/1
C0017689|T191|PSC|CDR0000038989|PDQ|glucagonoma|8152/1
C1882278|T191|SY|CDR0000038988|PDQ|interacinar cell pancreatic polypeptide tumor|8152/1
C0017689|T191|SY|CDR0000038989|PDQ|islet cell glucagonoma|8152/1
C1882278|T191|SY|CDR0000038988|PDQ|multiple hormonal syndrome, pancreatic|8152/1
C0017689|T191|SY|CDR0000038989|PDQ|pancreatic glucagonoma|8152/1
C1882278|T191|SY|CDR0000038988|PDQ|pancreatic multiple hormonal syndrome|8152/1
C1882278|T191|PSC|CDR0000038988|PDQ|pancreatic polypeptide tumor|8152/1
C0017689|T191|PT|R0121611|QMR|GLUCAGONOMA|8152/1
C0017689|T191|SY|Xa98N|RCD|Alpha cell adenoma|8152/1
C0017689|T191|PT|Xa98N|RCD|Glucagonoma|8152/1
C0017689|T191|PT|X50GW|RCD|Glucagonoma syndrome|8152/1
C0017689|T191|PT|BB5B4|RCDSY|Glucagonoma NOS|8152/1
C0017689|T191|IS|48538009|SNOMEDCT_US|Alpha cell adenoma|8152/1
C0017689|T191|SY|302823005|SNOMEDCT_US|Alpha cell adenoma|8152/1
C0017689|T191|SY|128855009|SNOMEDCT_US|Alpha cell tumor|8152/1
C0017689|T191|SYGB|128855009|SNOMEDCT_US|Alpha cell tumour|8152/1
C1266016|T191|PT|128644006|SNOMEDCT_US|Enteroglucagonoma|8152/1
C0017689|T191|OAP|48538009|SNOMEDCT_US|Glucagonoma|8152/1
C0017689|T191|PT|128855009|SNOMEDCT_US|Glucagonoma|8152/1
C0017689|T191|PT|302823005|SNOMEDCT_US|Glucagonoma|8152/1
C0017689|T191|IS|48538009|SNOMEDCT_US|Glucagonoma -RETIRED-|8152/1
C0017689|T191|OF|48538009|SNOMEDCT_US|Glucagonoma -RETIRED-|8152/1
C0017689|T191|PT|16424000|SNOMEDCT_US|Glucagonoma syndrome|8152/1
C0017689|T191|IS|16424000|SNOMEDCT_US|Glucagonoma syndrome, NOS|8152/1
C0017689|T191|IS|48538009|SNOMEDCT_US|Glucagonoma, NOS|8152/1
C0334282|T191|PT|MTHU004940|ICPC2ICD10ENG|alpha cell; tumor, malignant, pancreas|8152/3
C0334282|T191|PT|MTHU004939|ICPC2ICD10ENG|alpha cell; tumor, malignant, unspecified site|8152/3
C0334282|T191|PT|MTHU032351|ICPC2ICD10ENG|glucagonoma; malignant, pancreas|8152/3
C0334282|T191|PT|MTHU032350|ICPC2ICD10ENG|glucagonoma; malignant, unspecified site|8152/3
C0334282|T191|PT|MTHU047287|ICPC2ICD10ENG|malignant; glucagonoma, pancreas|8152/3
C0334282|T191|PT|MTHU047286|ICPC2ICD10ENG|malignant; glucagonoma, unspecified site|8152/3
C0334282|T191|PT|MTHU057093|ICPC2ICD10ENG|pancreas; alpha cell tumor, malignant|8152/3
C0334282|T191|PT|MTHU057125|ICPC2ICD10ENG|pancreas; glucagonoma, malignant|8152/3
C0334282|T191|PT|MTHU057137|ICPC2ICD10ENG|pancreas; malignant glucagonoma|8152/3
C0334282|T191|PT|MTHU057159|ICPC2ICD10ENG|pancreas; tumor, alpha cell, malignant|8152/3
C0334282|T191|PT|MTHU077012|ICPC2ICD10ENG|tumor; alpha cell, malignant, pancreas|8152/3
C0334282|T191|PT|MTHU077011|ICPC2ICD10ENG|tumor; alpha cell, malignant, unspecified site|8152/3
C1266017|T191|PT|271426|MEDCIN|malignant enteroglucagonoma|8152/3
C0334282|T191|PT|35209|MEDCIN|malignant glucagonoma of pancreas|8152/3
C0334282|T191|SY|35209|MEDCIN|malignant pancreatic glucagonoma|8152/3
C1266017|T191|OP|C65191|NCI|Malignant Enteroglucagonoma|8152/3
C1266017|T191|PT|C65191|NCI|Malignant Enteroglucagonoma|8152/3
C0334282|T191|SY|C65187|NCI|Malignant Glucagonoma|8152/3
C0334282|T191|PT|C65187|NCI|Malignant Pancreatic Glucagonoma|8152/3
C0334282|T191|SY|C65187|NCI|Pancreatic Alpha Cell Carcinoma|8152/3
C0334282|T191|DN|C65187|NCI_CTRP|Malignant Pancreatic Glucagonoma|8152/3
C0334282|T191|SY|CDR0000040032|PDQ|carcinoma, alpha cell, pancreatic|8152/3
C0334282|T191|SY|CDR0000040032|PDQ|carcinoma, glucagon producing|8152/3
C0334282|T191|SY|CDR0000040032|PDQ|carcinoma, glucagon secreting|8152/3
C0334282|T191|SY|CDR0000040032|PDQ|carcinoma, pancreatic alpha cell|8152/3
C0334282|T191|SY|CDR0000040032|PDQ|glucagon producing carcinoma|8152/3
C0334282|T191|SY|CDR0000040032|PDQ|glucagon secreting carcinoma|8152/3
C0334282|T191|SY|CDR0000040032|PDQ|Malignant Glucagonoma|8152/3
C0334282|T191|PT|CDR0000040032|PDQ|pancreatic alpha cell carcinoma|8152/3
C0334282|T191|SY|BB5B5|RCD|Malignant alpha cell tumour|8152/3
C0334282|T191|PT|BB5B5|RCD|Malignant glucagonoma|8152/3
C0334282|T191|SY|BB5B5|RCDAE|Malignant alpha cell tumor|8152/3
C0334282|T191|SY|66515009|SNOMEDCT_US|Alpha cell tumor, malignant|8152/3
C0334282|T191|SYGB|66515009|SNOMEDCT_US|Alpha cell tumour, malignant|8152/3
C1266017|T191|OAP|128645007|SNOMEDCT_US|Enteroglucagonoma, malignant|8152/3
C0334282|T191|PT|66515009|SNOMEDCT_US|Glucagonoma, malignant|8152/3
C0334282|T191|SY|66515009|SNOMEDCT_US|Malignant alpha cell tumor|8152/3
C0334282|T191|SYGB|66515009|SNOMEDCT_US|Malignant alpha cell tumour|8152/3
C0334282|T191|SY|66515009|SNOMEDCT_US|Malignant glucagonoma|8152/3
C0017150|T191|SY|0000005374|CHV|gastrin producing tumor|8153/1
C0017150|T191|PT|0000005374|CHV|gastrinoma|8153/1
C0017150|T191|SY|0000005374|CHV|gastrinomas|8153/1
C0017150|T191|PT|MTHU030557|ICPC2ICD10ENG|G cell; tumor, unspecified site|8153/1
C0017150|T191|PT|MTHU030434|ICPC2ICD10ENG|gastrinoma; unspecified site|8153/1
C0017150|T191|PT|MTHU077060|ICPC2ICD10ENG|tumor; G cell, unspecified site|8153/1
C0017150|T191|LLT|10017852|MDR|Gastrinoma|8153/1
C0017150|T191|PT|10017852|MDR|Gastrinoma|8153/1
C0017150|T191|PT|352610|MEDCIN|gastrinoma|8153/1
C0017150|T191|SY|352610|MEDCIN|neuroendocrine tumor gastrinoma|8153/1
C0017150|T191|PM|D015408|MSH|Gastrin Producing Tumor|8153/1
C0017150|T191|ET|D015408|MSH|Gastrin-Producing Tumor|8153/1
C0017150|T191|PM|D015408|MSH|Gastrin-Producing Tumors|8153/1
C0017150|T191|MH|D015408|MSH|Gastrinoma|8153/1
C0017150|T191|PM|D015408|MSH|Gastrinomas|8153/1
C0017150|T191|ET|D015408|MSH|Islet Cell Tumor, Ulcerogenic|8153/1
C0017150|T191|PM|D015408|MSH|Tumor, Gastrin-Producing|8153/1
C0017150|T191|PM|D015408|MSH|Tumors, Gastrin-Producing|8153/1
C0017150|T191|ET|D015408|MSH|Ulcerogenic Islet Cell Tumor|8153/1
C0017150|T191|SY|C3050|NCI|G Cell Tumor|8153/1
C0017150|T191|SY|C3050|NCI|G-Cell Gastrin Producing Tumor|8153/1
C0017150|T191|SY|C3050|NCI|G-Cell Tumor|8153/1
C0017150|T191|SY|C3050|NCI|Gastrin Secreting Tumor|8153/1
C0017150|T191|SY|C3050|NCI|Gastrin-Producing NET|8153/1
C0017150|T191|PT|C3050|NCI|Gastrin-Producing Neuroendocrine Tumor|8153/1
C0017150|T191|SY|C3050|NCI|Gastrinoma|8153/1
C0017150|T191|DN|C3050|NCI_CTRP|Gastrin-Producing Neuroendocrine Tumor|8153/1
C0017150|T191|PT|CDR0000044239|NCI_NCI-GLOSS|gastrinoma|8153/1
C0017150|T191|PSC|CDR0000038718|PDQ|gastrinoma|8153/1
C0017150|T191|SY|Xa98O|RCD|G cell tumour|8153/1
C0017150|T191|PT|Xa98O|RCD|Gastrinoma|8153/1
C0017150|T191|SY|Xa98O|RCDAE|G cell tumor|8153/1
C0017150|T191|PT|BB5C0|RCDSY|Gastrinoma NOS|8153/1
C0017150|T191|SY|16189002|SNOMEDCT_US|G cell tumor|8153/1
C0017150|T191|SY|302824004|SNOMEDCT_US|G cell tumor|8153/1
C0017150|T191|IS|16189002|SNOMEDCT_US|G cell tumor, NOS|8153/1
C0017150|T191|SYGB|302824004|SNOMEDCT_US|G cell tumour|8153/1
C0017150|T191|SYGB|16189002|SNOMEDCT_US|G cell tumour|8153/1
C0017150|T191|SY|16189002|SNOMEDCT_US|Gastrin cell tumor|8153/1
C0017150|T191|SYGB|16189002|SNOMEDCT_US|Gastrin cell tumour|8153/1
C0017150|T191|PT|302824004|SNOMEDCT_US|Gastrinoma|8153/1
C0017150|T191|PT|16189002|SNOMEDCT_US|Gastrinoma|8153/1
C0017150|T191|IS|16189002|SNOMEDCT_US|Gastrinoma, NOS|8153/1
C0334283|T191|PT|MTHU030555|ICPC2ICD10ENG|G cell; tumor, malignant, unspecified site|8153/3
C0334283|T191|PT|MTHU030432|ICPC2ICD10ENG|gastrinoma; malignant, unspecified site|8153/3
C0334283|T191|PT|MTHU047282|ICPC2ICD10ENG|malignant; gastrinoma, unspecified site|8153/3
C0334283|T191|PT|MTHU077058|ICPC2ICD10ENG|tumor; G cell, malignant, unspecified site|8153/3
C0334283|T191|LLT|10051709|MDR|Gastrinoma malignant|8153/3
C0334283|T191|PT|10051709|MDR|Gastrinoma malignant|8153/3
C0334283|T191|PT|271424|MEDCIN|malignant gastrinoma|8153/3
C0334283|T191|PT|C65188|NCI|Malignant Gastrinoma|8153/3
C0334283|T191|DN|C65188|NCI_CTRP|Malignant Gastrinoma|8153/3
C0334283|T191|SY|BB5C1|RCD|Malignant G cell tumour|8153/3
C0334283|T191|PT|BB5C1|RCD|Malignant gastrinoma|8153/3
C0334283|T191|SY|BB5C1|RCDAE|Malignant G cell tumor|8153/3
C0334283|T191|SY|19756007|SNOMEDCT_US|G cell tumor, malignant|8153/3
C0334283|T191|SYGB|19756007|SNOMEDCT_US|G cell tumour, malignant|8153/3
C0334283|T191|SY|19756007|SNOMEDCT_US|Gastrin cell tumor, malignant|8153/3
C0334283|T191|SYGB|19756007|SNOMEDCT_US|Gastrin cell tumour, malignant|8153/3
C0334283|T191|PT|19756007|SNOMEDCT_US|Gastrinoma, malignant|8153/3
C0334283|T191|SY|19756007|SNOMEDCT_US|Malignant G cell tumor|8153/3
C0334283|T191|SYGB|19756007|SNOMEDCT_US|Malignant G cell tumour|8153/3
C0334283|T191|SY|19756007|SNOMEDCT_US|Malignant gastrinoma|8153/3
C1301048|T191|PN|NOCODE|MTH|Mixed Ductal-Endocrine Carcinoma|8154/3
C2987162|T191|PT|C95460|NCI|Mixed Acinar-Neuroendocrine-Ductal Carcinoma of the Pancreas|8154/3
C1301048|T191|SY|C6879|NCI|Mixed Ductal-Endocrine Carcinoma|8154/3
C1301048|T191|SY|C6879|NCI|Mixed Ductal-Endocrine Carcinoma of the Pancreas|8154/3
C1301048|T191|PT|C6879|NCI|Mixed Ductal-Neuroendocrine Carcinoma of the Pancreas|8154/3
C1301048|T191|SY|TCGA|NCI|Mixed Ductal-Neuroendocrine Carcinoma of the Pancreas|8154/3
C1709050|T191|SY|C45843|NCI|Mixed Exocrine-Endocrine Carcinoma of the Pancreas|8154/3
C1709050|T191|SY|C45843|NCI|Pancreatic Carcinoma with Mixed Differentiation|8154/3
C1709050|T191|PT|C45843|NCI|Pancreatic Mixed Adenoneuroendocrine Carcinoma|8154/3
C1709050|T191|SY|C45843|NCI|Pancreatic Mixed Neuroendocrine-Non-Neuroendocrine Carcinoma|8154/3
C0334284|T191|PT|BB5B6|RCD|Mixed islet cell and exocrine adenocarcinoma|8154/3
C0334284|T191|AB|BB5B6|RCD|Mixed islet cell+exocr adenoca|8154/3
C1301047|T191|PT|396891002|SNOMEDCT_US|Mixed acinar-endocrine carcinoma|8154/3
C1301047|T191|SY|999000|SNOMEDCT_US|Mixed acinar-endocrine carcinoma|8154/3
C5190873|T191|PT|783209004|SNOMEDCT_US|Mixed acinar-endocrine-ductal carcinoma|8154/3
C1301048|T191|PT|396892009|SNOMEDCT_US|Mixed ductal-endocrine carcinoma|8154/3
C1301048|T191|SY|999000|SNOMEDCT_US|Mixed ductal-endocrine carcinoma|8154/3
C0334284|T191|PT|999000|SNOMEDCT_US|Mixed islet cell and exocrine adenocarcinoma|8154/3
C0011993|T191|PT|0000003868|CHV|vipoma|8155/1
C0011993|T191|SY|0000003868|CHV|vipomas|8155/1
C0011993|T191|DI|U002005|DXP|VIPOMA|8155/1
C0011993|T191|PT|10047430|MDR|Vipoma|8155/1
C0011993|T191|LLT|10047430|MDR|Vipoma|8155/1
C0011993|T191|ET|D003969|MSH|Diarrheogenic Islet Cell Tumor|8155/1
C0011993|T191|ET|D003969|MSH|Diarrheogenic Tumor|8155/1
C0011993|T191|PM|D003969|MSH|Diarrheogenic Tumors|8155/1
C0011993|T191|ET|D003969|MSH|Pancreatic VIPoma|8155/1
C0011993|T191|PM|D003969|MSH|Pancreatic VIPomas|8155/1
C0011993|T191|PM|D003969|MSH|Tumor, Diarrheogenic|8155/1
C0011993|T191|PM|D003969|MSH|Tumors, Diarrheogenic|8155/1
C0011993|T191|PM|D003969|MSH|Vasoactive Intestinal Peptide Producing Tumor|8155/1
C0011993|T191|ET|D003969|MSH|Vasoactive Intestinal Peptide-Producing Tumor|8155/1
C0011993|T191|MH|D003969|MSH|Vipoma|8155/1
C0011993|T191|PM|D003969|MSH|VIPoma, Pancreatic|8155/1
C0011993|T191|PM|D003969|MSH|Vipomas|8155/1
C0011993|T191|PM|D003969|MSH|VIPomas, Pancreatic|8155/1
C0011993|T191|PN|NOCODE|MTH|Vipoma|8155/1
C0011993|T191|SY|C26749|NCI|Vasoactive Intestinal Peptide Producing Neoplasm|8155/1
C0011993|T191|SY|C26749|NCI|Vasoactive Intestinal Peptide Producing Tumor|8155/1
C0011993|T191|SY|C26749|NCI|Vasoactive Intestinal Peptide Secreting Neoplasm|8155/1
C0011993|T191|SY|C26749|NCI|VIP Producing Neoplasm|8155/1
C0011993|T191|SY|C26749|NCI|VIP- Secreting Neoplasm|8155/1
C0011993|T191|SY|C26749|NCI|VIP- Secreting Tumor|8155/1
C0011993|T191|SY|C26749|NCI|VIP-Producing NET|8155/1
C0011993|T191|PT|C26749|NCI|VIP-Producing Neuroendocrine Tumor|8155/1
C0011993|T191|SY|C26749|NCI|VIPoma|8155/1
C0011993|T191|OP|CDR0000040023|PDQ|pancreatic alpha-D islet cell adenoma|8155/1
C0011993|T191|AB|X77nW|RCD|Vasoact intes peptide-secr tum|8155/1
C0011993|T191|PT|X77nW|RCD|Vasoactive intestinal peptide-secreting tumour|8155/1
C0011993|T191|SY|X77nW|RCD|VIP-oma - Vasoactive intestinal peptide-secreting tumour|8155/1
C0011993|T191|AB|X77nW|RCD|VIP-oma - VIP-secreting tumour|8155/1
C0011993|T191|PT|X77nW|RCDAE|Vasoactive intestinal peptide-secreting tumor|8155/1
C0011993|T191|SY|X77nW|RCDAE|VIP-oma - Vasoactive intestinal peptide-secreting tumor|8155/1
C0011993|T191|AB|X77nW|RCDAE|VIP-oma - VIP-secreting tumor|8155/1
C0011993|T191|OP|BB5y1|RCDSY|Vipoma|8155/1
C0011993|T191|PT|253005002|SNOMEDCT_US|Vasoactive intestinal peptide-secreting tumor|8155/1
C0011993|T191|PTGB|253005002|SNOMEDCT_US|Vasoactive intestinal peptide-secreting tumour|8155/1
C0011993|T191|SY|253005002|SNOMEDCT_US|VIP-oma - Vasoactive intestinal peptide-secreting tumor|8155/1
C0011993|T191|SYGB|253005002|SNOMEDCT_US|VIP-oma - Vasoactive intestinal peptide-secreting tumour|8155/1
C0011993|T191|PT|447643008|SNOMEDCT_US|Vipoma|8155/1
C1881600|T191|PN|NOCODE|MTH|Malignant Vipoma|8155/3
C1881600|T191|PT|C65189|NCI|Malignant Vipoma|8155/3
C1881600|T191|SY|31131002|SNOMEDCT_US|Vipoma|8155/3
C1881600|T191|PT|31131002|SNOMEDCT_US|Vipoma, malignant|8155/3
C0037661|T191|PT|0000011525|CHV|somatostatinoma|8156/1
C0037661|T191|DI|U001759|DXP|SOMATOSTATINOMA|8156/1
C0037661|T191|LLT|10041329|MDR|Somatostatinoma|8156/1
C0037661|T191|PT|10041329|MDR|Somatostatinoma|8156/1
C0037661|T191|MH|D013005|MSH|Somatostatinoma|8156/1
C0037661|T191|PM|D013005|MSH|Somatostatinomas|8156/1
C0037661|T191|PN|NOCODE|MTH|Somatostatinoma|8156/1
C0037661|T191|SY|C3379|NCI|Delta Cell Tumor|8156/1
C0037661|T191|SY|C3379|NCI|Somatostatin Cell Tumor|8156/1
C0037661|T191|SY|C3379|NCI|Somatostatin Producing Tumor|8156/1
C0037661|T191|SY|C3379|NCI|Somatostatin-Producing NET|8156/1
C0037661|T191|PT|C3379|NCI|Somatostatin-Producing Neuroendocrine Tumor|8156/1
C0037661|T191|SY|C3379|NCI|Somatostatin-Producing Tumor|8156/1
C0037661|T191|SY|C3379|NCI|Somatostatinoma|8156/1
C0037661|T191|SY|C3379|NCI|Tumor of Delta Cells|8156/1
C0037661|T191|SY|C3379|NCI|Tumor of the Delta Cells|8156/1
C0037661|T191|DN|C3379|NCI_CTRP|Somatostatin-Producing Neuroendocrine Tumor|8156/1
C0037661|T191|SY|X77nX|RCD|Delta cell tumour|8156/1
C0037661|T191|PT|X77nX|RCD|Somatostatinoma|8156/1
C0037661|T191|SY|X77nX|RCDAE|Delta cell tumor|8156/1
C0037661|T191|SY|253006001|SNOMEDCT_US|Delta cell tumor|8156/1
C0037661|T191|SYGB|253006001|SNOMEDCT_US|Delta cell tumour|8156/1
C0037661|T191|SY|128642005|SNOMEDCT_US|Somatostatin cell tumor|8156/1
C0037661|T191|SYGB|128642005|SNOMEDCT_US|Somatostatin cell tumour|8156/1
C0037661|T191|PT|128642005|SNOMEDCT_US|Somatostatinoma|8156/1
C0037661|T191|PT|253006001|SNOMEDCT_US|Somatostatinoma|8156/1
C1266015|T191|PT|271425|MEDCIN|malignant somatostatinoma|8156/3
C1266015|T191|SY|C65190|NCI|Delta Cell Carcinoma|8156/3
C1266015|T191|PT|C65190|NCI|Malignant Somatostatinoma|8156/3
C1266015|T191|DN|C65190|NCI_CTRP|Malignant Somatostatinoma|8156/3
C1266015|T191|SY|128643000|SNOMEDCT_US|Somatostatin cell tumor, malignant|8156/3
C1266015|T191|SYGB|128643000|SNOMEDCT_US|Somatostatin cell tumour, malignant|8156/3
C1266015|T191|PT|128643000|SNOMEDCT_US|Somatostatinoma, malignant|8156/3
C1266016|T191|OP|C66925|NCI|Enteroglucagonoma|8157/1
C1266016|T191|PT|C66925|NCI|Enteroglucagonoma|8157/1
C1266016|T191|PT|128644006|SNOMEDCT_US|Enteroglucagonoma|8157/1
C1266017|T191|PT|271426|MEDCIN|malignant enteroglucagonoma|8157/3
C1266017|T191|PT|C65191|NCI|Malignant Enteroglucagonoma|8157/3
C1266017|T191|OP|C65191|NCI|Malignant Enteroglucagonoma|8157/3
C1266017|T191|OAP|128645007|SNOMEDCT_US|Enteroglucagonoma, malignant|8157/3
C1335300|T191|SY|C27466|NCI|Ectopic ACTH-Producing Pancreatic Neuroendocrine Tumor|8158/1
C2986655|T191|PT|C94759|NCI|Functioning Endocrine Neoplasm|8158/1
C1335300|T191|SY|C27466|NCI|Pancreatic ACTH Producing NET|8158/1
C1335300|T191|SY|C27466|NCI|Pancreatic ACTH Producing Neuroendocrine Tumor|8158/1
C1335300|T191|SY|C27466|NCI|Pancreatic ACTH Producing Tumor|8158/1
C1335300|T191|PT|C27466|NCI|Pancreatic ACTH-Producing Neuroendocrine Tumor|8158/1
C1335300|T191|SY|C27466|NCI|Pancreatic ACTH-Producing Neuroendocrine Tumor With Cushing Syndrome|8158/1
C1335300|T191|SY|C27466|NCI|Pancreatic Adrenocorticotropic Hormone Producing Tumor|8158/1
C2986655|T191|PT|CDR0000458094|NCI_NCI-GLOSS|functioning tumor|8158/1
C3472604|T191|PT|450891001|SNOMEDCT_US|Functioning endocrine tumor|8158/1
C3472604|T191|PTGB|450891001|SNOMEDCT_US|Functioning endocrine tumour|8158/1
C0008309|T191|SY|0000002856|CHV|adenoma bile duct|8160/0
C0008309|T191|SY|0000002856|CHV|bile duct adenoma|8160/0
C0008309|T191|SY|0000002856|CHV|bile duct adenomas|8160/0
C0008309|T191|PT|0000002856|CHV|cholangioma|8160/0
C0008309|T191|SY|0000002856|CHV|cholangiomas|8160/0
C0008309|T191|PT|MTHU003501|ICPC2ICD10ENG|adenoma; bile duct|8160/0
C0008309|T191|PT|MTHU030173|ICPC2ICD10ENG|bile duct; adenoma|8160/0
C0008309|T191|PT|MTHU016244|ICPC2ICD10ENG|cholangioma|8160/0
C0008309|T191|LLT|10008592|MDR|Cholangioadenoma|8160/0
C0008309|T191|PT|10008592|MDR|Cholangioadenoma|8160/0
C0008309|T191|MH|D002759|MSH|Adenoma, Bile Duct|8160/0
C0008309|T191|PM|D002759|MSH|Adenomas, Bile Duct|8160/0
C0008309|T191|PM|D002759|MSH|Bile Duct Adenoma|8160/0
C0008309|T191|PM|D002759|MSH|Bile Duct Adenomas|8160/0
C0008309|T191|ET|D002759|MSH|Cholangioma|8160/0
C0008309|T191|PM|D002759|MSH|Cholangiomas|8160/0
C0008309|T191|PN|NOCODE|MTH|Bile duct adenoma|8160/0
C0008309|T191|SY|C2942|NCI|Adenoma of Bile Duct|8160/0
C0008309|T191|SY|C2942|NCI|Adenoma of the Bile Duct|8160/0
C0008309|T191|PT|C2942|NCI|Bile Duct Adenoma|8160/0
C0008309|T191|SY|C2942|NCI|Cholangioadenoma|8160/0
C0008309|T191|SY|C2942|NCI|Cholangioma|8160/0
C0008309|T191|SY|C2942|NCI_CDISC|Adenoma of Bile Duct|8160/0
C0008309|T191|SY|C2942|NCI_CDISC|Adenoma of the Bile Duct|8160/0
C0008309|T191|SY|C2942|NCI_CDISC|Cholangioadenoma|8160/0
C0008309|T191|SY|C2942|NCI_CDISC|Cholangioma|8160/0
C0008309|T191|PT|C2942|NCI_CDISC|CHOLANGIOMA, BENIGN|8160/0
C0008309|T191|SY|C2942|NCI_CDISC|Hepatocholangiocellular Adenoma|8160/0
C0008309|T191|SY|C2942|NCI_CDISC|Hepatocholangioma|8160/0
C0008309|T191|PT|XM1FD|RCD|Bile duct adenoma|8160/0
C0008309|T191|SY|XM1FD|RCD|Cholangioma|8160/0
C0008309|T191|OP|BB5D0|RCDSY|Bile duct adenoma|8160/0
C0008309|T191|PT|39471001|SNOMEDCT_US|Bile duct adenoma|8160/0
C0008309|T191|PT|424091006|SNOMEDCT_US|Cholangioadenoma|8160/0
C0008309|T191|SY|39471001|SNOMEDCT_US|Cholangioma|8160/0
C0206698|T191|PT|0000021030|CHV|cholangiocarcinoma|8160/3
C0206698|T191|SY|0000021030|CHV|cholangiocarcinomas|8160/3
C0206698|T191|SY|0000021030|CHV|cholangiocellular carcinoma|8160/3
C0206698|T191|SY|HP:0030153|HPO|Bile duct cancer|8160/3
C0206698|T191|PT|HP:0030153|HPO|Cholangiocarcinoma|8160/3
C0206698|T191|ET|C22.1|ICD10CM|Cholangiocarcinoma|8160/3
C0206698|T191|PT|MTHU016239|ICPC2ICD10ENG|cholangiocarcinoma; unspecified site|8160/3
C0206698|T191|PT|10008593|MDR|Cholangiocarcinoma|8160/3
C0206698|T191|LLT|10008593|MDR|Cholangiocarcinoma|8160/3
C0206698|T191|LLT|10008595|MDR|Cholangiocarcinoma NOS|8160/3
C0206698|T191|PT|10077861|MDR|Cholangiosarcoma|8160/3
C0206698|T191|LLT|10077861|MDR|Cholangiosarcoma|8160/3
C0206698|T191|PT|353455|MEDCIN|Cholangiocarcinoma of biliary tract|8160/3
C0206698|T191|SY|353455|MEDCIN|malignant neoplasm of biliary tract cholangiocarcinoma|8160/3
C0206698|T191|SY|5905|MEDLINEPLUS|Cholangiocarcinoma|8160/3
C0206698|T191|ET|5905|MEDLINEPLUS|Cholangiocarcinoma|8160/3
C0206698|T191|PM|D018281|MSH|Carcinoma, Cholangiocellular|8160/3
C0206698|T191|PM|D018281|MSH|Carcinomas, Cholangiocellular|8160/3
C0206698|T191|MH|D018281|MSH|Cholangiocarcinoma|8160/3
C0206698|T191|PM|D018281|MSH|Cholangiocarcinomas|8160/3
C0206698|T191|ET|D018281|MSH|Cholangiocellular Carcinoma|8160/3
C0206698|T191|PM|D018281|MSH|Cholangiocellular Carcinomas|8160/3
C0206698|T191|PN|NOCODE|MTH|Cholangiocarcinoma|8160/3
C0206698|T191|AB|C4436|NCI|CC|8160/3
C0206698|T191|PT|C4436|NCI|Cholangiocarcinoma|8160/3
C0206698|T191|SY|TCGA|NCI|Cholangiocarcinoma|8160/3
C0206698|T191|OP|C4436|NCI|Cholangiocellular Carcinoma|8160/3
C0206698|T191|PT|C4436|NCI_CDISC|CHOLANGIOCARCINOMA, MALIGNANT|8160/3
C0206698|T191|SY|C4436|NCI_CDISC|Cholangiocellular Carcinoma|8160/3
C0206698|T191|PT|C4436|NCI_CPTAC|Cholangiocarcinoma|8160/3
C0206698|T191|SY|10004669|NCI_CTEP-SDC|Cholangiocar.- intra/extrahepatic|8160/3
C0206698|T191|PT|C4436|NCI_CTRP|Cholangiocarcinoma|8160/3
C0206698|T191|PT|CDR0000335064|NCI_NCI-GLOSS|cholangiocarcinoma|8160/3
C0206698|T191|PT|CDR0000046473|NCI_NCI-GLOSS|cholangiosarcoma|8160/3
C0206698|T191|AB|XaDbr|RCD|Cholangiocarcin biliary tract|8160/3
C0206698|T191|PT|BB5D1|RCD|Cholangiocarcinoma|8160/3
C0206698|T191|PT|XaDbr|RCD|Cholangiocarcinoma of biliary tract|8160/3
C0206698|T191|PT|70179006|SNOMEDCT_US|Cholangiocarcinoma|8160/3
C0206698|T191|PT|312104005|SNOMEDCT_US|Cholangiocarcinoma of biliary tract|8160/3
C0206698|T191|SY|70179006|SNOMEDCT_US|Cholangiocellular carcinoma|8160/3
C0334285|T191|PT|MTHU030194|ICPC2ICD10ENG|bile duct; cystadenoma|8161/0
C0334285|T191|PT|MTHU020308|ICPC2ICD10ENG|cystadenoma; bile duct|8161/0
C0334285|T191|SY|C4129|NCI|Bile Duct Cystadenoma|8161/0
C0334285|T191|PT|C4129|NCI|Bile Duct Mucinous Cystic Neoplasm|8161/0
C0334285|T191|SY|C4129|NCI|Cystadenoma of Bile Duct|8161/0
C0334285|T191|SY|C4129|NCI|Cystadenoma of the Bile Duct|8161/0
C0334285|T191|PT|BB5D2|RCD|Bile duct cystadenoma|8161/0
C0334285|T191|PT|83025009|SNOMEDCT_US|Bile duct cystadenoma|8161/0
C0334286|T191|PT|MTHU030193|ICPC2ICD10ENG|bile duct; cystadenocarcinoma|8161/3
C0334286|T191|PT|MTHU020291|ICPC2ICD10ENG|cystadenocarcinoma; bile duct|8161/3
C0334286|T191|PT|217840|MEDCIN|cystadenocarcinoma of bile duct|8161/3
C0334286|T191|SY|217840|MEDCIN|liver neoplasm malignant bile duct cystadenocarcinoma|8161/3
C0334286|T191|SY|C4130|NCI|Bile Duct Cystadenocarcinoma|8161/3
C0334286|T191|PT|C4130|NCI|Bile Duct Mucinous Cystic Neoplasm with an Associated Invasive Carcinoma|8161/3
C0334286|T191|SY|C4130|NCI|Biliary Cystadenocarcinoma|8161/3
C0334286|T191|SY|C4130|NCI|Cystadenocarcinoma of Bile Duct|8161/3
C0334286|T191|SY|C4130|NCI|Cystadenocarcinoma of the Bile Duct|8161/3
C0334286|T191|PT|BB5D3|RCD|Bile duct cystadenocarcinoma|8161/3
C0334286|T191|PT|50422007|SNOMEDCT_US|Bile duct cystadenocarcinoma|8161/3
C0206702|T191|PT|0000021033|CHV|klatskin tumor|8162/3
C0206702|T191|SY|0000021033|CHV|klatskin tumors|8162/3
C0206702|T191|SY|0000021033|CHV|klatskin's tumor|8162/3
C0206702|T191|SY|0000021033|CHV|klatskin's tumour|8162/3
C0206702|T191|SY|0000021033|CHV|klatskins tumor|8162/3
C0206702|T191|SY|0000021033|CHV|klatzkin tumor|8162/3
C0206702|T191|PT|MTHU041472|ICPC2ICD10ENG|Klatskin|8162/3
C0206702|T191|PT|MTHU041473|ICPC2ICD10ENG|Klatskin; tumor|8162/3
C0206702|T191|PT|MTHU077078|ICPC2ICD10ENG|tumor; Klatskin|8162/3
C0206702|T191|LLT|10074878|MDR|Hilar cholangiocarcinoma|8162/3
C0206702|T191|LLT|10074874|MDR|Klatskin tumor|8162/3
C0206702|T191|LLT|10074877|MDR|Klatskin tumour|8162/3
C0206702|T191|PM|D018285|MSH|Cholangiocarcinoma, Hilar|8162/3
C0206702|T191|PM|D018285|MSH|Cholangiocarcinomas, Hilar|8162/3
C0206702|T191|ET|D018285|MSH|Hilar Cholangiocarcinoma|8162/3
C0206702|T191|PM|D018285|MSH|Hilar Cholangiocarcinomas|8162/3
C0206702|T191|MH|D018285|MSH|Klatskin Tumor|8162/3
C0206702|T191|ET|D018285|MSH|Klatskin's Tumor|8162/3
C0206702|T191|PM|D018285|MSH|Klatskins Tumor|8162/3
C0206702|T191|PM|D018285|MSH|Tumor, Klatskin|8162/3
C0206702|T191|PM|D018285|MSH|Tumor, Klatskin's|8162/3
C0206702|T191|SY|C36077|NCI|Hilar CC|8162/3
C0206702|T191|PT|C36077|NCI|Hilar Cholangiocarcinoma|8162/3
C0206702|T191|SY|C36077|NCI|Klatskin Tumor|8162/3
C3273047|T191|SY|C96804|NCI|Perihilar Bile Duct Carcinoma|8162/3
C3273047|T191|SY|C96804|NCI|Perihilar ICC|8162/3
C3273047|T191|PT|C96804|NCI|Perihilar Intrahepatic Cholangiocarcinoma|8162/3
C0206702|T191|DN|C36077|NCI_CTRP|Hilar Cholangiocarcinoma|8162/3
C0206702|T191|PT|CDR0000335074|NCI_NCI-GLOSS|Klatskin tumor|8162/3
C0206702|T191|SY|CDR0000040913|PDQ|Klatskin tumor|8162/3
C0206702|T191|PT|X77nj|RCD|Klatskin's tumour|8162/3
C0206702|T191|OP|BB5y2|RCD|Klatskin's tumour morphology|8162/3
C0206702|T191|PT|X77nj|RCDAE|Klatskin's tumor|8162/3
C0206702|T191|OP|BB5y2|RCDAE|Klatskin's tumor morphology|8162/3
C0206702|T191|IS|BB5y2|RCDSA|Klatskin's tumor|8162/3
C0206702|T191|IS|BB5y2|RCDSY|Klatskin's tumour|8162/3
C0206702|T191|SY|6492006|SNOMEDCT_US|Klatskin tumor|8162/3
C0206702|T191|SY|253017000|SNOMEDCT_US|Klatskin tumor|8162/3
C0206702|T191|SYGB|253017000|SNOMEDCT_US|Klatskin tumour|8162/3
C0206702|T191|SYGB|6492006|SNOMEDCT_US|Klatskin tumour|8162/3
C0206702|T191|PT|6492006|SNOMEDCT_US|Klatskin's tumor|8162/3
C0206702|T191|PT|253017000|SNOMEDCT_US|Klatskin's tumor|8162/3
C0206702|T191|SY|6492006|SNOMEDCT_US|Klatskin's tumor morphology|8162/3
C0206702|T191|PTGB|6492006|SNOMEDCT_US|Klatskin's tumour|8162/3
C0206702|T191|PTGB|253017000|SNOMEDCT_US|Klatskin's tumour|8162/3
C0206702|T191|SYGB|6492006|SNOMEDCT_US|Klatskin's tumour morphology|8162/3
C3272434|T191|SY|C95914|NCI|Ampullary Low Grade Intraepithelial Neoplasia|8163/0
C3272434|T191|PT|C95914|NCI|Ampullary Noninvasive Pancreatobiliary Papillary Neoplasm with Low Grade Dysplasia|8163/0
C3272433|T191|PT|C95913|NCI|Ampullary Noninvasive Papillary Neoplasm, Pancreatobiliary Type|8163/0
C3272433|T191|SY|C95913|NCI|Noninvasive Papillary Neoplasm, Pancreatobiliary Type|8163/0
C3472605|T191|PT|450892008|SNOMEDCT_US|Non-invasive pancreatobiliary neoplasm|8163/0
C3272435|T191|SY|C95915|NCI|Ampullary High Grade Intraepithelial Neoplasia|8163/2
C3272435|T191|PT|C95915|NCI|Ampullary Noninvasive Pancreatobiliary Papillary Neoplasm with High Grade Dysplasia|8163/2
C3472606|T191|PT|450893003|SNOMEDCT_US|Papillary neoplasm, pancreatobiliary-type, with high grade intraepithelial neoplasia|8163/2
C3272461|T191|PT|C95963|NCI|Ampulla of Vater Pancreatobiliary Type Adenocarcinoma|8163/3
C3472607|T191|SY|450894009|SNOMEDCT_US|Adenocarcinoma, pancreatobiliary-type|8163/3
C3472607|T191|PT|450894009|SNOMEDCT_US|Pancreatobiliary-type carcinoma|8163/3
C0206669|T191|PT|0047129|CCPSS|LIVER ADENOMA|8170/0
C0206669|T191|PT|0047124|CCPSS|LIVER CELL ADENOMA|8170/0
C0206669|T191|SY|0000038513|CHV|adenoma liver|8170/0
C0206669|T191|SY|0000038513|CHV|adenomas hepatic|8170/0
C0206669|T191|SY|0000038513|CHV|adenomas liver|8170/0
C0206669|T191|PT|0000038513|CHV|hepatic adenoma|8170/0
C0206669|T191|PT|0000021008|CHV|hepatocellular adenoma|8170/0
C0206669|T191|SY|0000021008|CHV|hepatocellular adenomas|8170/0
C0206669|T191|SY|0000038513|CHV|liver adenoma|8170/0
C0206669|T191|SY|0000021008|CHV|liver cell adenoma|8170/0
C0206669|T191|GT|NEOPL LIVER|CST|ADENOMA LIVER|8170/0
C0206669|T191|SY|HP:0012028|HPO|Hepatic adenoma|8170/0
C0206669|T191|PT|HP:0012028|HPO|Hepatocellular adenoma|8170/0
C0206669|T191|SY|HP:0012028|HPO|Liver cell adenoma|8170/0
C0206669|T191|PT|MTHU003508|ICPC2ICD10ENG|adenoma; hepatocellular|8170/0
C0206669|T191|PT|MTHU003511|ICPC2ICD10ENG|adenoma; liver cell|8170/0
C0206669|T191|PT|MTHU010316|ICPC2ICD10ENG|benign; hepatoma|8170/0
C0206669|T191|PT|MTHU034361|ICPC2ICD10ENG|hepatocellular; adenoma|8170/0
C0206669|T191|PT|MTHU034385|ICPC2ICD10ENG|hepatoma; benign|8170/0
C0206669|T191|PT|MTHU045062|ICPC2ICD10ENG|liver cell; adenoma|8170/0
C0206669|T191|PT|D78013|ICPC2P|Adenoma;hepatic|8170/0
C0206669|T191|PTN|D78013|ICPC2P|hepatic adenoma|8170/0
C0206669|T191|LLT|10001235|MDR|Adenoma liver|8170/0
C0206669|T191|LLT|10019629|MDR|Hepatic adenoma|8170/0
C0206669|T191|PT|10019629|MDR|Hepatic adenoma|8170/0
C0206669|T191|LLT|10019827|MDR|Hepatocellular adenoma|8170/0
C0206669|T191|PT|31585|MEDCIN|benign adenoma of liver|8170/0
C0206669|T191|SY|31585|MEDCIN|hepatic adenoma|8170/0
C0206669|T191|ET|D018248|MSH|Adenoma, Hepatocellular|8170/0
C0206669|T191|MH|D018248|MSH|Adenoma, Liver Cell|8170/0
C0206669|T191|PM|D018248|MSH|Adenomas, Hepatocellular|8170/0
C0206669|T191|PM|D018248|MSH|Adenomas, Liver Cell|8170/0
C0206669|T191|PM|D018248|MSH|Benign Hepatoma|8170/0
C0206669|T191|PM|D018248|MSH|Benign Hepatomas|8170/0
C0206669|T191|PM|D018248|MSH|Hepatocellular Adenoma|8170/0
C0206669|T191|PM|D018248|MSH|Hepatocellular Adenomas|8170/0
C0206669|T191|ET|D018248|MSH|Hepatoma, Benign|8170/0
C0206669|T191|PM|D018248|MSH|Hepatomas, Benign|8170/0
C0206669|T191|PM|D018248|MSH|Liver Cell Adenoma|8170/0
C0206669|T191|PM|D018248|MSH|Liver Cell Adenomas|8170/0
C0206669|T191|PN|NOCODE|MTH|Hepatocellular Adenoma|8170/0
C0206669|T191|SY|C3758|NCI|Adenoma of Liver Cells|8170/0
C0206669|T191|SY|C3758|NCI|Adenoma of the Liver Cells|8170/0
C0206669|T191|AB|C3758|NCI|HCA|8170/0
C0206669|T191|PT|C3758|NCI|Hepatocellular Adenoma|8170/0
C0206669|T191|SY|C3758|NCI|Liver Cell Adenoma|8170/0
C0206669|T191|SY|C3758|NCI_CDISC|Adenoma of Liver Cells|8170/0
C0206669|T191|SY|C3758|NCI_CDISC|Adenoma of the Liver Cells|8170/0
C0206669|T191|PT|C3758|NCI_CDISC|ADENOMA, HEPATOCELLULAR, BENIGN|8170/0
C0206669|T191|SY|C3758|NCI_CDISC|HCA|8170/0
C0206669|T191|SY|C3758|NCI_CDISC|Liver Cell Adenoma|8170/0
C0206669|T191|PT|R0121629|QMR|HEPATOCELLULAR ADENOMA <S>|8170/0
C0206669|T191|SY|BB5D4|RCD|Benign hepatoma|8170/0
C0206669|T191|SY|BB5D4|RCD|HCA - Hepatocellular adenoma|8170/0
C0206669|T191|SY|BB5D4|RCD|Hepatocellular adenoma|8170/0
C0206669|T191|PT|BB5D4|RCD|Liver cell adenoma|8170/0
C0206669|T191|PT|424263008|SNOMEDCT_US|Adenoma of liver|8170/0
C0206669|T191|SY|78058005|SNOMEDCT_US|Benign hepatoma|8170/0
C0206669|T191|SY|78058005|SNOMEDCT_US|HCA - Hepatocellular adenoma|8170/0
C0206669|T191|SY|78058005|SNOMEDCT_US|Hepatocellular adenoma|8170/0
C0206669|T191|SY|78058005|SNOMEDCT_US|Hepatoma, benign|8170/0
C0206669|T191|PT|78058005|SNOMEDCT_US|Liver cell adenoma|8170/0
C2239176|T191|ET|0000004597|AOD|hepatocellular carcinoma|8170/3
C2239176|T191|ET|0000004595|AOD|hepatoma|8170/3
C2239176|T191|NP|0000023073|AOD|liver cell carcinoma|8170/3
C2239176|T191|PT|1017965|CCPSS|HEPATOCELLULAR CARCINOMA|8170/3
C2239176|T191|SY|0000006061|CHV|hepatic carcinoma|8170/3
C2239176|T191|SY|0000006061|CHV|hepatocarcinoma|8170/3
C2239176|T191|SY|0000006061|CHV|hepatocellular carcinoma|8170/3
C2239176|T191|SY|0000006061|CHV|hepatoma|8170/3
C2239176|T191|SY|0000006061|CHV|hepatomas|8170/3
C2239176|T191|SY|0000006061|CHV|liver carcinoma|8170/3
C2239176|T191|PT|0000006061|CHV|liver cell cancer|8170/3
C2239176|T191|SY|0000006061|CHV|liver cell carcinoma|8170/3
C2239176|T191|PT|144|COSTAR|CARCINOMA OF LIVER|8170/3
C2239176|T191|PT|NOCODE|COSTAR|Hepatic Carcinoma|8170/3
C2239176|T191|PT|NOCODE|COSTAR|Hepatoma|8170/3
C2239176|T191|PT|2003-4684|CSP|hepatocellular carcinoma|8170/3
C2239176|T191|ET|2003-4684|CSP|hepatoma|8170/3
C2239176|T191|GT|CARCINOMA LIVER|CST|CARCINOMA LIVER|8170/3
C2239176|T191|PT|CARCINOMA LIVER|CST|CARCINOMA OF LIVER|8170/3
C2239176|T191|PT|HEPATOMA|CST|HEPATOMA|8170/3
C2239176|T191|GT|CARCINOMA LIVER|CST|LIVER CARCINOMA|8170/3
C2239176|T191|DI|U000820|DXP|HEPATOCARCINOMA|8170/3
C2239176|T191|SY|NOCODE|DXP|HEPATOCELLULAR CARCINOMA|8170/3
C2239176|T191|SY|NOCODE|DXP|HEPATOMA|8170/3
C2239176|T191|SY|NOCODE|DXP|LIVER CANCER, HEPATOCARCINOMA|8170/3
C2239176|T191|SY|NOCODE|DXP|LIVER CELL CARCINOMA|8170/3
C2239176|T191|SY|NOCODE|DXP|LIVER, CARCINOMA, PRIMARY|8170/3
C2239176|T191|PT|HP:0001402|HPO|Hepatocellular carcinoma|8170/3
C2239176|T191|PT|C22.0|ICD10|Liver cell carcinoma|8170/3
C2239176|T191|ET|C22.0|ICD10CM|Hepatocellular carcinoma|8170/3
C2239176|T191|PT|C22.0|ICD10CM|Liver cell carcinoma|8170/3
C2239176|T191|AB|C22.0|ICD10CM|Liver cell carcinoma|8170/3
C2239176|T191|PT|MTHU014785|ICPC2ICD10ENG|carcinoma; hepatic cell|8170/3
C2239176|T191|PT|MTHU014763|ICPC2ICD10ENG|carcinoma; hepatocellular|8170/3
C2239176|T191|PT|MTHU045063|ICPC2ICD10ENG|hepatic cell; carcinoma|8170/3
C2239176|T191|PT|MTHU034360|ICPC2ICD10ENG|hepatocarcinoma|8170/3
C2239176|T191|PT|MTHU034362|ICPC2ICD10ENG|hepatocellular; carcinoma|8170/3
C2239176|T191|PT|MTHU034384|ICPC2ICD10ENG|hepatoma|8170/3
C2239176|T191|PT|D77001|ICPC2P|Hepatoma|8170/3
C2239176|T191|PTN|D77001|ICPC2P|hepatoma|8170/3
C2239176|T191|PT|U002176|LCH|Hepatoma|8170/3
C2239176|T191|PT|sh85060302|LCH_NW|Hepatoma|8170/3
C2239176|T191|LLT|10049010|MDR|Carcinoma hepatocellular|8170/3
C2239176|T191|LLT|10007416|MDR|Carcinoma liver|8170/3
C2239176|T191|LLT|10048491|MDR|Carcinoma of liver|8170/3
C2239176|T191|LLT|10073071|MDR|Hepatocellular carcinoma|8170/3
C2239176|T191|PT|10073071|MDR|Hepatocellular carcinoma|8170/3
C2239176|T191|LLT|10019838|MDR|Hepatoma|8170/3
C2239176|T191|LLT|10024658|MDR|Liver carcinoma|8170/3
C2239176|T191|PT|217827|MEDCIN|carcinoma of liver|8170/3
C2239176|T191|PT|31588|MEDCIN|hepatocellular carcinoma of liver|8170/3
C2239176|T191|SY|217827|MEDCIN|liver neoplasm malignant carcinoma|8170/3
C2239176|T191|SY|353786|MEDCIN|liver neoplasm malignant carcinoma primary|8170/3
C2239176|T191|PT|353786|MEDCIN|Primary carcinoma of liver|8170/3
C2239176|T191|SY|309|MEDLINEPLUS|Hepatocellular carcinoma|8170/3
C2239176|T191|ET|309|MEDLINEPLUS|Hepatocellular Carcinoma|8170/3
C2239176|T191|PM|D006528|MSH|Adult Liver Cancer|8170/3
C2239176|T191|PM|D006528|MSH|Adult Liver Cancers|8170/3
C2239176|T191|PM|D006528|MSH|Cancer, Adult Liver|8170/3
C2239176|T191|PM|D006528|MSH|Cancers, Adult Liver|8170/3
C2239176|T191|MH|D006528|MSH|Carcinoma, Hepatocellular|8170/3
C2239176|T191|PM|D006528|MSH|Carcinoma, Liver Cell|8170/3
C2239176|T191|PM|D006528|MSH|Carcinomas, Hepatocellular|8170/3
C2239176|T191|PM|D006528|MSH|Carcinomas, Liver Cell|8170/3
C2239176|T191|PM|D006528|MSH|Cell Carcinoma, Liver|8170/3
C2239176|T191|PM|D006528|MSH|Cell Carcinomas, Liver|8170/3
C2239176|T191|ET|D006528|MSH|Hepatocellular Carcinoma|8170/3
C2239176|T191|PM|D006528|MSH|Hepatocellular Carcinomas|8170/3
C2239176|T191|ET|D006528|MSH|Hepatoma|8170/3
C2239176|T191|PM|D006528|MSH|Hepatomas|8170/3
C2239176|T191|ET|D006528|MSH|Liver Cancer, Adult|8170/3
C2239176|T191|PM|D006528|MSH|Liver Cancers, Adult|8170/3
C2239176|T191|ET|D006528|MSH|Liver Cell Carcinoma|8170/3
C2239176|T191|ET|D006528|MSH|Liver Cell Carcinoma, Adult|8170/3
C2239176|T191|PM|D006528|MSH|Liver Cell Carcinomas|8170/3
C2239176|T191|PN|NOCODE|MTH|Liver carcinoma|8170/3
C2239176|T191|ET|155.0|MTHICD9|Carcinoma of liver cell|8170/3
C2239176|T191|ET|155.0|MTHICD9|Carcinoma of liver, specified as primary|8170/3
C2239176|T191|ET|155.0|MTHICD9|Hepatocellular carcinoma|8170/3
C2239176|T191|SY|C3099|NCI|Carcinoma of Liver Cells|8170/3
C2239176|T191|SY|C3099|NCI|Carcinoma of the Liver Cells|8170/3
C2239176|T191|AB|C3099|NCI|HCC|8170/3
C2239176|T191|PT|C3099|NCI|Hepatocellular Carcinoma|8170/3
C2239176|T191|SY|TCGA|NCI|Hepatocellular Carcinoma|8170/3
C2239176|T191|SY|C3099|NCI|Hepatoma|8170/3
C2239176|T191|SY|C3099|NCI|Liver Cell Carcinoma|8170/3
C2239176|T191|SY|C3099|NCI|Primary Carcinoma of Liver Cells|8170/3
C2239176|T191|SY|C3099|NCI|Primary Carcinoma of the Liver Cells|8170/3
C2239176|T191|SY|C3099|NCI_CDISC|Carcinoma of Liver Cells|8170/3
C2239176|T191|SY|C3099|NCI_CDISC|Carcinoma of the Liver Cells|8170/3
C2239176|T191|PT|C3099|NCI_CDISC|CARCINOMA, HEPATOCELLULAR, MALIGNANT|8170/3
C2239176|T191|SY|C3099|NCI_CDISC|HCC|8170/3
C2239176|T191|SY|C3099|NCI_CDISC|Hepatoma|8170/3
C2239176|T191|SY|C3099|NCI_CDISC|Liver Cell Carcinoma|8170/3
C2239176|T191|SY|C3099|NCI_CDISC|Primary Carcinoma of Liver Cells|8170/3
C2239176|T191|SY|C3099|NCI_CDISC|Primary Carcinoma of the Liver Cells|8170/3
C2239176|T191|PT|C3099|NCI_CPTAC|Hepatocellular Carcinoma|8170/3
C2239176|T191|PT|10049010|NCI_CTEP-SDC|Hepatocellular carcinoma|8170/3
C2239176|T191|DN|C3099|NCI_CTRP|Hepatocellular Cancer|8170/3
C2239176|T191|PT|C3099|NCI_CTRP|Hepatocellular Carcinoma|8170/3
C2239176|T191|PT|CDR0000046363|NCI_NCI-GLOSS|hepatocellular carcinoma|8170/3
C2239176|T191|PT|CDR0000046661|NCI_NCI-GLOSS|hepatoma|8170/3
C2239176|T191|PT|R0121630|QMR|HEPATOCELLULAR CARCINOMA|8170/3
C2239176|T191|SY|B1503|RCD|HCC - Hepatocellular carcinoma|8170/3
C2239176|T191|SY|B1503|RCD|Hepatocarcinoma|8170/3
C2239176|T191|PT|B1503|RCD|Hepatocellular carcinoma|8170/3
C2239176|T191|SY|B1503|RCD|LCC - Liver cell carcinoma|8170/3
C2239176|T191|SY|B1503|RCD|Liver carcinoma|8170/3
C2239176|T191|SY|B1503|RCD|Liver cell carcinoma|8170/3
C2239176|T191|SY|B1503|RCD|Malignant hepatoma|8170/3
C2239176|T191|OP|B1500|RCD|Primary carcinoma of liver|8170/3
C2239176|T191|OA|BB5D5|RCDSY|Hepatocellular ca. NOS|8170/3
C2239176|T191|OP|BB5D5|RCDSY|Hepatocellular carcinoma NOS|8170/3
C2239176|T191|SY|109841003|SNOMEDCT_US|HCC - Hepatocellular carcinoma|8170/3
C2239176|T191|SY|25370001|SNOMEDCT_US|Hepatocarcinoma|8170/3
C2239176|T191|SY|109841003|SNOMEDCT_US|Hepatocarcinoma|8170/3
C2239176|T191|PT|25370001|SNOMEDCT_US|Hepatocellular carcinoma|8170/3
C2239176|T191|SY|109841003|SNOMEDCT_US|Hepatocellular carcinoma|8170/3
C2239176|T191|IS|25370001|SNOMEDCT_US|Hepatocellular carcinoma, NOS|8170/3
C2239176|T191|SY|25370001|SNOMEDCT_US|Hepatoma|8170/3
C2239176|T191|SY|25370001|SNOMEDCT_US|Hepatoma, malignant|8170/3
C2239176|T191|IS|25370001|SNOMEDCT_US|Hepatoma, NOS|8170/3
C2239176|T191|SY|109841003|SNOMEDCT_US|LCC - Liver cell carcinoma|8170/3
C2239176|T191|OAS|269547001|SNOMEDCT_US|Liver carcinoma|8170/3
C2239176|T191|SY|109841003|SNOMEDCT_US|Liver carcinoma|8170/3
C2239176|T191|OAS|154469006|SNOMEDCT_US|Liver carcinoma|8170/3
C2239176|T191|PT|109841003|SNOMEDCT_US|Liver cell carcinoma|8170/3
C2239176|T191|SY|25370001|SNOMEDCT_US|Liver cell carcinoma|8170/3
C2239176|T191|SY|109841003|SNOMEDCT_US|Malignant hepatoma|8170/3
C2239176|T191|PT|187769009|SNOMEDCT_US|Primary carcinoma of liver|8170/3
C2239176|T191|IT|1023|WHO|HEPATOMA|8170/3
C0334287|T191|PT|MTHU014764|ICPC2ICD10ENG|carcinoma; hepatocellular, fibrolamellar|8171/3
C0334287|T191|PT|MTHU028192|ICPC2ICD10ENG|fibrolamellar; hepatocellular carcinoma|8171/3
C0334287|T191|PT|MTHU034363|ICPC2ICD10ENG|hepatocellular; carcinoma, fibrolamellar|8171/3
C0334287|T191|PT|217841|MEDCIN|fibrolamellar hepatocellular carcinoma of liver|8171/3
C0334287|T191|NM|C537258|MSH|Fibrolamellar hepatocellular carcinoma|8171/3
C0334287|T191|CE|C537258|MSH|Fibrolamellar variant of hepatocellular carcinoma|8171/3
C0334287|T191|PN|NOCODE|MTH|Fibrolamellar Hepatocellular Carcinoma|8171/3
C0334287|T191|PT|C4131|NCI|Fibrolamellar Carcinoma|8171/3
C0334287|T191|SY|TCGA|NCI|Fibrolamellar Carcinoma|8171/3
C0334287|T191|SY|C4131|NCI|Fibrolamellar Carcinoma of Liver Cells|8171/3
C0334287|T191|SY|C4131|NCI|Fibrolamellar Carcinoma of the Liver Cells|8171/3
C0334287|T191|SY|C4131|NCI|Fibrolamellar Hepatocellular Carcinoma|8171/3
C0334287|T191|AB|C4131|NCI|FLC|8171/3
C0334287|T191|SY|C4131|NCI|Hepatocellular Fibrolamellar Carcinoma|8171/3
C0334287|T191|SY|C4131|NCI|Liver Cell Fibrolamellar Carcinoma|8171/3
C0334287|T191|SY|C4131|NCI|Oncocytic Hepatocellular Tumor|8171/3
C0334287|T191|SY|C4131|NCI|Polygonal Cell Type Hepatocellular Carcinoma with Fibrous Stroma|8171/3
C0334287|T191|PT|C4131|NCI_CPTAC|Fibrolamellar Carcinoma|8171/3
C0334287|T191|DN|C4131|NCI_CTRP|Fibrolamellar Cancer|8171/3
C0334287|T191|AB|X77nk|RCD|Fibrolamellar hepatocell ca|8171/3
C0334287|T191|PT|X77nk|RCD|Fibrolamellar hepatocellular carcinoma|8171/3
C0334287|T191|OA|BB5D8|RCDSY|Hepatocell carcin, fibrolam|8171/3
C0334287|T191|OP|BB5D8|RCDSY|Hepatocellular carcinoma, fibrolamellar|8171/3
C0334287|T191|PT|253018005|SNOMEDCT_US|Fibrolamellar hepatocellular carcinoma|8171/3
C0334287|T191|PT|15619004|SNOMEDCT_US|Hepatocellular carcinoma, fibrolamellar|8171/3
C1266018|T191|PT|C27388|NCI|Scirrhous Hepatocellular Carcinoma|8172/3
C1266018|T191|SY|C27388|NCI|Sclerosing Hepatic Carcinoma|8172/3
C1266018|T191|SY|C27388|NCI|Sclerosing Hepatocellular Carcinoma|8172/3
C1266018|T191|DN|C27388|NCI_CTRP|Scirrhous Hepatocellular Cancer|8172/3
C1266018|T191|PT|128646008|SNOMEDCT_US|Hepatocellular carcinoma, scirrhous|8172/3
C1266018|T191|SY|128646008|SNOMEDCT_US|Sclerosing hepatic carcinoma|8172/3
C1266019|T191|PT|217843|MEDCIN|spindle cell hepatocellular carcinoma of liver|8173/3
C1710014|T191|PT|C43627|NCI|Sarcomatoid Hepatocellular Carcinoma|8173/3
C1710014|T191|SY|C43627|NCI|Sarcomatous Hepatocellular Carcinoma|8173/3
C1710014|T191|DN|C43627|NCI_CTRP|Sarcomatoid Hepatocellular Cancer|8173/3
C1266019|T191|SY|128648009|SNOMEDCT_US|Hepatocellular carcinoma, sarcomatoid|8173/3
C1266019|T191|PT|128648009|SNOMEDCT_US|Hepatocellular carcinoma, spindle cell variant|8173/3
C1266020|T191|PT|217844|MEDCIN|clear cell hepatocellular carcinoma of liver|8174/3
C1333067|T191|SY|C5754|NCI|Clear Cell Carcinoma of Liver Cells|8174/3
C1333067|T191|SY|C5754|NCI|Clear Cell Carcinoma of the Liver Cells|8174/3
C1333067|T191|PT|C5754|NCI|Clear Cell Hepatocellular Carcinoma|8174/3
C1333067|T191|SY|C5754|NCI|Hepatocellular Clear Cell Carcinoma|8174/3
C1333067|T191|SY|C5754|NCI|Liver Cell Clear Cell Carcinoma|8174/3
C1333067|T191|DN|C5754|NCI_CTRP|Clear Cell Hepatocellular Cancer|8174/3
C1266020|T191|PT|128649001|SNOMEDCT_US|Hepatocellular carcinoma, clear cell type|8174/3
C1709568|T191|PN|NOCODE|MTH|Pleomorphic Hepatocellular Carcinoma|8175/3
C1709568|T191|PT|C43625|NCI|Pleomorphic Hepatocellular Carcinoma|8175/3
C1709568|T191|DN|C43625|NCI_CTRP|Pleomorphic Hepatocellular Cancer|8175/3
C1266021|T191|PT|128650001|SNOMEDCT_US|Hepatocellular carcinoma, pleomorphic type|8175/3
C0476108|T191|OP|BB5D6|RCDSY|Hepatocholangioma, benign|8180/0
C0476108|T191|PT|110456001|SNOMEDCT_US|Hepatocholangioma, benign|8180/0
C0221287|T191|SY|NOCODE|DXP|CHOLANGIOHEPATOMA|8180/3
C0221287|T191|SY|NOCODE|DXP|HEPATOCELLULAR, CHOLANGIOCARCINOMA COMBINED|8180/3
C0221287|T191|DI|U000821|DXP|HEPATOCHOLANGIOCARCINOMA|8180/3
C0221287|T191|PT|MTHU016238|ICPC2ICD10ENG|cholangiocarcinoma; with hepatocellular carcinoma|8180/3
C0221287|T191|PT|MTHU016240|ICPC2ICD10ENG|cholangiohepatoma|8180/3
C0221287|T191|PT|MTHU034365|ICPC2ICD10ENG|hepatocellular carcinoma; cholangiocarcinoma|8180/3
C0221287|T191|PT|MTHU034366|ICPC2ICD10ENG|hepatocholangiocarcinoma|8180/3
C0221287|T191|LLT|10073076|MDR|Combined hepatocellular and cholangiocarcinoma|8180/3
C0221287|T191|PT|10027761|MDR|Mixed hepatocellular cholangiocarcinoma|8180/3
C0221287|T191|LLT|10027761|MDR|Mixed hepatocellular cholangiocarcinoma|8180/3
C0221287|T191|PT|39426|MEDCIN|hepatocellular carcinoma and cholangiocarcinoma|8180/3
C0221287|T191|SY|39426|MEDCIN|liver neoplasm hepatocellular carcinoma & cholangiocarcinoma|8180/3
C0221287|T191|PN|NOCODE|MTH|Combined Hepatocellular Carcinoma and Cholangiocarcinoma|8180/3
C0221287|T191|SY|C3828|NCI|Carcinoma of Liver and Intrahepatic Biliary Tract|8180/3
C0221287|T191|SY|C3828|NCI|Carcinoma of the Liver and Intrahepatic Biliary Tract|8180/3
C0221287|T191|SY|C3828|NCI|Cholangiohepatoma|8180/3
C0221287|T191|PT|C3828|NCI|Combined Hepatocellular Carcinoma and Cholangiocarcinoma|8180/3
C0221287|T191|SY|C3828|NCI|Hepatocholangiocarcinoma|8180/3
C0221287|T191|SY|C3828|NCI|Liver and Intrahepatic Biliary Tract Carcinoma|8180/3
C0221287|T191|SY|C3828|NCI|Mixed Hepatocellular Cholangiocarcinoma|8180/3
C0221287|T191|PT|CDR0000752915|PDQ|adult primary mixed hepatocellular cholangiocarcinoma|8180/3
C0221287|T191|SY|CDR0000752915|PDQ|carcinoma of liver and intrahepatic biliary tract|8180/3
C0221287|T191|SY|CDR0000752915|PDQ|carcinoma of the liver and intrahepatic biliary tract|8180/3
C0221287|T191|SY|CDR0000752915|PDQ|cholangiohepatoma|8180/3
C0221287|T191|SY|CDR0000752915|PDQ|combined hepatocellular carcinoma and cholangiocarcinoma|8180/3
C0221287|T191|SY|CDR0000752915|PDQ|hepatocholangiocarcinoma|8180/3
C0221287|T191|SY|CDR0000752915|PDQ|liver and intrahepatic biliary tract carcinoma|8180/3
C0221287|T191|AB|XM1FE|RCD|Comb hepatocell ca+cholangioca|8180/3
C0221287|T191|PT|XM1FE|RCD|Combined hepatocellular carcinoma and cholangiocarcinoma|8180/3
C0221287|T191|SY|XM1FE|RCD|Hepatocholangiocarcinoma|8180/3
C0221287|T191|AB|XM1FE|RCD|Mixed hepatocell+bile duct ca|8180/3
C0221287|T191|SY|XM1FE|RCD|Mixed hepatocellular and bile duct carcinoma|8180/3
C0221287|T191|OA|BB5D7|RCDSY|Comb.hepatocell./cholang.ca|8180/3
C0221287|T191|OP|BB5D7|RCDSY|Combined hepatocellular carcinoma and cholangiocarcinoma|8180/3
C0221287|T191|PT|52178006|SNOMEDCT_US|Combined hepatocellular carcinoma and cholangiocarcinoma|8180/3
C0221287|T191|PT|274902006|SNOMEDCT_US|Combined hepatocellular carcinoma and cholangiocarcinoma|8180/3
C0221287|T191|SY|52178006|SNOMEDCT_US|Hepatocholangiocarcinoma|8180/3
C0221287|T191|SY|274902006|SNOMEDCT_US|Hepatocholangiocarcinoma|8180/3
C0221287|T191|SY|52178006|SNOMEDCT_US|Mixed hepatocellular and bile duct carcinoma|8180/3
C0221287|T191|SY|274902006|SNOMEDCT_US|Mixed hepatocellular and bile duct carcinoma|8180/3
C0205651|T191|PEP|D000236|MSH|Adenoma, Trabecular|8190/0
C0205651|T191|PM|D000236|MSH|Adenomas, Trabecular|8190/0
C0205651|T191|PM|D000236|MSH|Trabecular Adenoma|8190/0
C0205651|T191|PM|D000236|MSH|Trabecular Adenomas|8190/0
C0205651|T191|PT|C3688|NCI|Trabecular Adenoma|8190/0
C0205651|T191|PT|BB5E.|RCD|Trabecular adenoma|8190/0
C0205651|T191|PT|21930005|SNOMEDCT_US|Trabecular adenoma|8190/0
C0302182|T191|PT|271476|MEDCIN|trabecular adenocarcinoma|8190/3
C0302182|T191|PT|C4068|NCI|Trabecular Adenocarcinoma|8190/3
C0302182|T191|SY|C4068|NCI|Trabecular Carcinoma|8190/3
C0302182|T191|PT|BB5F.|RCD|Trabecular adenocarcinoma|8190/3
C0302182|T191|SY|BB5F.|RCD|Trabecular carcinoma|8190/3
C0302182|T191|PT|29792007|SNOMEDCT_US|Trabecular adenocarcinoma|8190/3
C0302182|T191|SY|29792007|SNOMEDCT_US|Trabecular carcinoma|8190/3
C1266045|T191|SY|C27253|NCI|Kidney Embryonal Adenoma|8191/0
C1266045|T191|PT|C27253|NCI|Metanephric Adenoma|8191/0
C0334288|T191|PT|BB5G.|RCD|Embryonal adenoma|8191/0
C0334288|T191|PT|59120003|SNOMEDCT_US|Embryonal adenoma|8191/0
C1266045|T191|PT|128670007|SNOMEDCT_US|Metanephric adenoma|8191/0
C1851526|T046|SY|0000056370|CHV|cylindromas dermal|8200/0
C1851526|T046|SY|0000056370|CHV|tumors turban|8200/0
C1851526|T046|SY|0000057839|CHV|tumors turban|8200/0
C1851526|T046|PT|0000056370|CHV|turban tumor|8200/0
C1851526|T046|PT|0000057839|CHV|turban tumor|8200/0
C1305968|T191|PT|HP:0031024|HPO|Cylindroma|8200/0
C1851526|T046|PT|MTHU077165|ICPC2ICD10ENG|tumor; turban|8200/0
C1851526|T046|PT|MTHU077004|ICPC2ICD10ENG|turban tumor|8200/0
C1851526|T046|PT|MTHU077003|ICPC2ICD10ENG|turban; tumor|8200/0
C1305968|T191|LLT|10012425|MDR|Dermal cylindroma|8200/0
C1851526|T046|PT|6380|MEDCIN|turban tumor|8200/0
C1305968|T191|CE|C536611|MSH|Ancell-Spiegler cylindromas|8200/0
C1305968|T191|CE|C536611|MSH|Cylindromas, Dermal Eccrine|8200/0
C1305968|T191|CE|C536611|MSH|Cylindromatosis, familial|8200/0
C1305968|T191|CE|C536611|MSH|Dermal Eccrine Cylindroma|8200/0
C1305968|T191|NM|C536611|MSH|Familial cylindromatosis|8200/0
C1305968|T191|CE|C536611|MSH|Familial Trichoepithelioma|8200/0
C1305968|T191|CE|C536611|MSH|Turban tumor syndrome|8200/0
C1305968|T191|CE|C536611|MSH|Turban tumors|8200/0
C1851526|T046|PN|NOCODE|MTH|Ancell-Spiegler cylindromas|8200/0
C1305968|T191|PN|NOCODE|MTH|Eccrine dermal cylindroma|8200/0
C1851526|T046|SY|C43352|NCI|Ancell-Spiegler Syndrome|8200/0
C1305968|T191|PT|C27094|NCI|Cylindroma|8200/0
C1305968|T191|SY|C27094|NCI|Cylindroma of Skin|8200/0
C1305968|T191|SY|C27094|NCI|Cylindroma of the Skin|8200/0
C1305968|T191|SY|C27094|NCI|Dermal Cylindroma|8200/0
C1851526|T046|PT|C43352|NCI|Turban Tumor|8200/0
C1851526|T046|SY|C43352|NCI|Turban Tumor Syndrome|8200/0
C1305968|T191|SY|XM1FF|RCD|Cylindroma of skin|8200/0
C1305968|T191|SY|XM1FF|RCD|Dermal cylindroma|8200/0
C1305968|T191|PT|XM1FF|RCD|Eccrine dermal cylindroma|8200/0
C1305968|T191|SY|XM1FF|RCD|Spiegler's tumour|8200/0
C1305968|T191|SY|XM1FF|RCD|Turban tumour|8200/0
C1305968|T191|SY|XM1FF|RCDAE|Spiegler's tumor|8200/0
C1305968|T191|SY|XM1FF|RCDAE|Turban tumor|8200/0
C1305968|T191|OP|BB5H.|RCDSY|Eccrine dermal cylindroma|8200/0
C3839386|T191|PT|703550009|SNOMEDCT_US|Cylindroma of breast|8200/0
C1851526|T046|OAS|212546007|SNOMEDCT_US|Cylindroma of skin|8200/0
C1851526|T046|PT|447147008|SNOMEDCT_US|Cylindroma of skin|8200/0
C1851526|T046|SY|64773009|SNOMEDCT_US|Cylindroma of skin|8200/0
C1305968|T191|SY|274903001|SNOMEDCT_US|Cylindroma of skin|8200/0
C1305968|T191|SY|274903001|SNOMEDCT_US|Dermal cylindroma|8200/0
C1305968|T191|PT|274903001|SNOMEDCT_US|Eccrine dermal cylindroma|8200/0
C1851526|T046|OAP|212546007|SNOMEDCT_US|Eccrine dermal cylindroma|8200/0
C1851526|T046|PT|64773009|SNOMEDCT_US|Eccrine dermal cylindroma|8200/0
C1305968|T191|SY|274903001|SNOMEDCT_US|Eccrine dermal cylindroma of skin|8200/0
C1305968|T191|SY|274903001|SNOMEDCT_US|Spiegler's tumor|8200/0
C1305968|T191|SYGB|274903001|SNOMEDCT_US|Spiegler's tumour|8200/0
C1305968|T191|SY|274903001|SNOMEDCT_US|Turban tumor|8200/0
C1851526|T046|SY|64773009|SNOMEDCT_US|Turban tumor|8200/0
C1851526|T046|IS|211710004|SNOMEDCT_US|turban tumor|8200/0
C1851526|T046|PT|211710004|SNOMEDCT_US|Turban tumor|8200/0
C1851526|T046|IS|211710004|SNOMEDCT_US|turban tumour|8200/0
C1851526|T046|PTGB|211710004|SNOMEDCT_US|Turban tumour|8200/0
C1851526|T046|SYGB|64773009|SNOMEDCT_US|Turban tumour|8200/0
C1305968|T191|SYGB|274903001|SNOMEDCT_US|Turban tumour|8200/0
C0010606|T191|SY|0000003536|CHV|adenocystic carcinoma|8200/3
C0010606|T191|SY|0000003536|CHV|adenoid cystic cancer|8200/3
C0010606|T191|PT|0000003536|CHV|adenoid cystic carcinoma|8200/3
C0010606|T191|SY|0000003536|CHV|adenoid cystic carcinomas|8200/3
C0010606|T191|SY|0000003536|CHV|carcinoma adenoid cystic|8200/3
C0010606|T191|SY|0000003536|CHV|cylindroma|8200/3
C0010606|T191|SY|0000003536|CHV|cylindromas|8200/3
C0010606|T191|PT|sh91002009|LCH_NW|Adenoid cystic carcinoma|8200/3
C0010606|T191|PT|10053231|MDR|Adenoid cystic carcinoma|8200/3
C0010606|T191|LLT|10053231|MDR|Adenoid cystic carcinoma|8200/3
C0010606|T191|LLT|10011729|MDR|Cylindroma|8200/3
C0010606|T191|PT|271437|MEDCIN|adenoid cystic carcinoma|8200/3
C0346017|T191|PT|231615|MEDCIN|adenoid cystic carcinoma of skin|8200/3
C0346017|T191|PT|357601|MEDCIN|Adenoid cystic eccrine carcinoma of skin|8200/3
C0346017|T191|SY|357601|MEDCIN|skin neop malignant adnexa w/ eccrine differentiation adenoid cystic carcinoma|8200/3
C0010606|T191|ET|D003528|MSH|Adenocystic Carcinoma|8200/3
C0010606|T191|PM|D003528|MSH|Adenocystic Carcinomas|8200/3
C0010606|T191|PM|D003528|MSH|Adenoid Cystic Carcinoma|8200/3
C0010606|T191|PM|D003528|MSH|Adenoid Cystic Carcinomas|8200/3
C0010606|T191|PM|D003528|MSH|Carcinoma, Adenocystic|8200/3
C0010606|T191|MH|D003528|MSH|Carcinoma, Adenoid Cystic|8200/3
C0010606|T191|PM|D003528|MSH|Carcinomas, Adenocystic|8200/3
C0010606|T191|PM|D003528|MSH|Carcinomas, Adenoid Cystic|8200/3
C0010606|T191|ET|D003528|MSH|Cylindroma|8200/3
C0010606|T191|PM|D003528|MSH|Cylindromas|8200/3
C0010606|T191|PM|D003528|MSH|Cystic Carcinoma, Adenoid|8200/3
C0010606|T191|PM|D003528|MSH|Cystic Carcinomas, Adenoid|8200/3
C0010606|T191|PN|NOCODE|MTH|Adenoid Cystic Carcinoma|8200/3
C0010606|T191|SY|C2970|NCI|Adenocystic Carcinoma|8200/3
C0010606|T191|SY|TCGA|NCI|Adenoid Cystic Carcinoma|8200/3
C0010606|T191|PT|C2970|NCI|Adenoid Cystic Carcinoma|8200/3
C0346017|T191|SY|C4471|NCI|Adenoid Cystic Carcinoma of Skin|8200/3
C0346017|T191|SY|C4471|NCI|Adenoid Cystic Carcinoma of the Skin|8200/3
C0346017|T191|SY|C4471|NCI|Adenoid Cystic Cutaneous Carcinoma|8200/3
C0346017|T191|PT|C4471|NCI|Adenoid Cystic Skin Carcinoma|8200/3
C0010606|T191|SY|C2970|NCI|Cylindroid Adenocarcinoma|8200/3
C0346017|T191|SY|C4471|NCI|Primary Cutaneous Adenocystic Carcinoma|8200/3
C0010606|T191|PT|C2970|NCI_CPTAC|Adenoid Cystic Carcinoma|8200/3
C0010606|T191|PT|CDR0000046022|NCI_NCI-GLOSS|adenoid cystic cancer|8200/3
C0010606|T191|SY|Xa98T|RCD|Adenocystic carcinoma|8200/3
C0346017|T191|AB|X78Sh|RCD|Adenoid cystc eccrin carcinoma|8200/3
C0010606|T191|OP|XE1wT|RCD|Adenoid cystic carcinoma|8200/3
C0346017|T191|AB|X78Sh|RCD|Adenoid cystic eccrine carcin|8200/3
C0346017|T191|PT|X78Sh|RCD|Adenoid cystic eccrine carcinoma|8200/3
C0346017|T191|SY|X78Sh|RCD|Adenoid cystic eccrine carcinoma of skin|8200/3
C0010606|T191|SY|Xa98T|RCD|Cylindroid adenocarcinoma|8200/3
C0010606|T191|SY|Xa98T|RCD|Cylindroid bronchial adenoma|8200/3
C0010606|T191|PT|Xa98T|RCD|Cylindroma|8200/3
C0346017|T191|AB|X78Sh|RCD|Prim cut adenocystic carcinoma|8200/3
C0346017|T191|SY|X78Sh|RCD|Primary cutaneous adenocystic carcinoma|8200/3
C0010606|T191|SY|11671000|SNOMEDCT_US|Adenocarcinoma, cylindroid|8200/3
C0010606|T191|SY|11671000|SNOMEDCT_US|Adenocystic carcinoma|8200/3
C0010606|T191|IS|302827006|SNOMEDCT_US|Adenocystic carcinoma|8200/3
C0010606|T191|PT|11671000|SNOMEDCT_US|Adenoid cystic carcinoma|8200/3
C0346017|T191|PT|399968001|SNOMEDCT_US|Adenoid cystic eccrine carcinoma|8200/3
C0346017|T191|PT|254711000|SNOMEDCT_US|Adenoid cystic eccrine carcinoma|8200/3
C0346017|T191|SY|254711000|SNOMEDCT_US|Adenoid cystic eccrine carcinoma of skin|8200/3
C0010606|T191|IS|11671000|SNOMEDCT_US|Bronchial adenoma, cylindroid|8200/3
C0010606|T191|IS|302827006|SNOMEDCT_US|Cylindroid adenocarcinoma|8200/3
C0010606|T191|IS|302827006|SNOMEDCT_US|Cylindroid bronchial adenoma|8200/3
C0010606|T191|PT|302827006|SNOMEDCT_US|Cylindroma|8200/3
C0346017|T191|SY|254711000|SNOMEDCT_US|Primary cutaneous adenocystic carcinoma|8200/3
C4511178|T191|PT|725504002|SNOMEDCT_US|Thymic carcinoma with adenoid cystic carcinoma-like features|8200/3
C1266022|T191|PT|271390|MEDCIN|cribriform carcinoma in situ|8201/2
C1334248|T191|SY|C5138|NCI|Cribriform DCIS of Breast|8201/2
C1334248|T191|SY|C5138|NCI|Cribriform DCIS of the Breast|8201/2
C1334248|T191|SY|C5138|NCI|Cribriform Ductal Breast Carcinoma in situ|8201/2
C1334248|T191|SY|C5138|NCI|Cribriform Ductal Carcinoma in situ of Breast|8201/2
C1334248|T191|SY|C5138|NCI|Cribriform Ductal Carcinoma in situ of the Breast|8201/2
C1334248|T191|SY|C5138|NCI|DCIS of Breast with Cribriform Pattern|8201/2
C1334248|T191|SY|C5138|NCI|DCIS of the Breast with Cribriform Pattern|8201/2
C1334248|T191|SY|C5138|NCI|Ductal Carcinoma in situ of Breast with Cribriform Pattern|8201/2
C1334248|T191|SY|C5138|NCI|Ductal Carcinoma in situ of the Breast with Cribriform Pattern|8201/2
C1334248|T191|PT|C5138|NCI|Intraductal Cribriform Breast Adenocarcinoma|8201/2
C1334248|T191|SY|C5138|NCI|Non-Infiltrating Cribriform Ductal Breast Carcinoma|8201/2
C1334248|T191|SY|C5138|NCI|Non-Invasive Cribriform Ductal Breast Carcinoma|8201/2
C1266022|T191|PT|128879006|SNOMEDCT_US|Cribriform carcinoma in situ|8201/2
C1266022|T191|SY|128879006|SNOMEDCT_US|Ductal carcinoma in situ, cribriform type|8201/2
C0205643|T191|PT|0000020664|CHV|cribriform carcinoma|8201/3
C4296895|T191|LA|LA26494-7|LNC|Cribriform comedo-type adenocarcinoma|8201/3
C0205643|T191|PT|271438|MEDCIN|cribriform carcinoma|8201/3
C0205643|T191|PEP|D000230|MSH|Carcinoma, Cribriform|8201/3
C0205643|T191|PM|D000230|MSH|Carcinomas, Cribriform|8201/3
C0205643|T191|PM|D000230|MSH|Cribriform Carcinoma|8201/3
C0205643|T191|PM|D000230|MSH|Cribriform Carcinomas|8201/3
C3272812|T191|PT|C96488|NCI|Colorectal Cribriform Comedo-Type Adenocarcinoma|8201/3
C0205643|T191|PT|C3680|NCI|Cribriform Carcinoma|8201/3
C0205643|T191|PT|C3680|NCI_CPTAC|Cribriform Carcinoma|8201/3
C0205643|T191|PT|BB5K.|RCD|Cribriform carcinoma|8201/3
C0205643|T191|PT|30156004|SNOMEDCT_US|Cribriform carcinoma|8201/3
C4296895|T191|PT|733838009|SNOMEDCT_US|Cribriform comedo-type adenocarcinoma|8201/3
C0205643|T191|SY|30156004|SNOMEDCT_US|Ductal carcinoma, cribriform type|8201/3
C0205648|T191|PEP|D000236|MSH|Adenoma, Microcystic|8202/0
C0205648|T191|PM|D000236|MSH|Adenomas, Microcystic|8202/0
C0205648|T191|PM|D000236|MSH|Microcystic Adenoma|8202/0
C0205648|T191|PM|D000236|MSH|Microcystic Adenomas|8202/0
C0205648|T191|PT|C3685|NCI|Microcystic Adenoma|8202/0
C0205648|T191|PT|X77nI|RCD|Microcystic adenoma|8202/0
C0205648|T191|PT|79494009|SNOMEDCT_US|Microcystic adenoma|8202/0
C0205648|T191|OAP|189580001|SNOMEDCT_US|Microcystic adenoma|8202/0
C0205648|T191|OF|189580001|SNOMEDCT_US|Microcystic adenoma|8202/0
C1266023|T191|SY|0000056676|CHV|lactate adenoma|8204/0
C1266023|T191|PT|0000056676|CHV|lactating adenoma|8204/0
C1266023|T191|PT|C9473|NCI|Lactating Adenoma|8204/0
C1266023|T191|SY|C9473|NCI|Pregnancy Adenoma|8204/0
C1266023|T191|PT|128651002|SNOMEDCT_US|Lactating adenoma|8204/0
C0206677|T191|PT|0062825|CCPSS|POLYP ADENOMATOUS|8210/0
C0206677|T191|PT|0000021014|CHV|adenomatous polyp|8210/0
C0206677|T191|SY|0000021014|CHV|adenomatous polyps|8210/0
C0206677|T191|PT|4005-0002|CSP|adenomatous polyp|8210/0
C0206677|T191|ET|4005-0002|CSP|polypoid adenoma|8210/0
C0206677|T191|ET|D28|ICD10CM|adenomatous polyp|8210/0
C0206677|T191|PM|D018256|MSH|Adenomatous Polyp|8210/0
C0206677|T191|MH|D018256|MSH|Adenomatous Polyps|8210/0
C0206677|T191|PM|D018256|MSH|Polyp, Adenomatous|8210/0
C0206677|T191|PM|D018256|MSH|Polyps, Adenomatous|8210/0
C0206677|T191|PN|NOCODE|MTH|Adenomatous Polyps|8210/0
C0206677|T191|PT|C3764|NCI|Adenomatous Polyp|8210/0
C0206677|T191|SY|C3764|NCI|Polypoid Adenoma|8210/0
C0206677|T191|DN|C3764|NCI_CTRP|Adenomatous Polyp|8210/0
C0206677|T191|PT|CDR0000590650|PDQ|adenomatous polyp|8210/0
C0206677|T191|SY|CDR0000590650|PDQ|Polypoid Adenoma|8210/0
C0206677|T191|PT|Xa98W|RCD|Adenomatous polyp|8210/0
C0206677|T191|SY|Xa98W|RCD|Polypoid adenoma|8210/0
C0206677|T191|OP|BB5L0|RCDSY|Adenomatous polyp NOS|8210/0
C0206677|T191|PT|82375006|SNOMEDCT_US|Adenomatous polyp|8210/0
C0206677|T191|IS|82375006|SNOMEDCT_US|Adenomatous polyp, NOS|8210/0
C0206677|T191|SY|82375006|SNOMEDCT_US|Polypoid adenoma|8210/0
C0334290|T191|PT|271387|MEDCIN|adenocarcinoma in situ in adenomatous polyp|8210/2
C1377630|T191|PN|NOCODE|MTH|Adenocarcinoma in situ in a polyp|8210/2
C0334290|T191|PN|NOCODE|MTH|Adenocarcinoma in situ in adenomatous polyp|8210/2
C1377630|T191|PT|C7680|NCI|Adenocarcinoma In Situ in a Polyp|8210/2
C0334290|T191|PT|C7678|NCI|Adenocarcinoma In Situ in Adenomatous Polyp|8210/2
C1377630|T191|OA|BB5L1|RCD|Adenoca in situ in a polyp|8210/2
C0334290|T191|AB|BB5L2|RCD|Adenoca situ in adenom polyp|8210/2
C0334290|T191|AB|BB5L2|RCD|Adenoca situ in polyp adenoma|8210/2
C1377630|T191|OP|BB5L1|RCD|Adenocarcinoma in situ in a polyp|8210/2
C0334290|T191|PT|BB5L2|RCD|Adenocarcinoma in situ in adenomatous polyp|8210/2
C0334290|T191|SY|BB5L2|RCD|Adenocarcinoma in situ in polypoid adenoma|8210/2
C0334290|T191|AB|BB5L2|RCD|Ca in situ in adenomat polyp|8210/2
C0334290|T191|SY|BB5L2|RCD|Carcinoma in situ in adenomatous polyp|8210/2
C0334290|T191|AB|BB5L2|RCDSY|Adencar in situ,adeno polyp|8210/2
C1377630|T191|IS|60286009|SNOMEDCT_US|Adenocarcinoma in situ in a polyp|8210/2
C1377630|T191|PT|189598002|SNOMEDCT_US|Adenocarcinoma in situ in a polyp|8210/2
C1377630|T191|IS|60286009|SNOMEDCT_US|Adenocarcinoma in situ in a polyp, NOS|8210/2
C0334290|T191|PT|60286009|SNOMEDCT_US|Adenocarcinoma in situ in adenomatous polyp|8210/2
C0334290|T191|SY|60286009|SNOMEDCT_US|Adenocarcinoma in situ in polypoid adenoma|8210/2
C0334290|T191|SY|60286009|SNOMEDCT_US|Carcinoma in situ in adenomatous polyp|8210/2
C1321861|T191|PT|271473|MEDCIN|adenocarcinoma in adenomatous polyp|8210/3
C1321861|T191|PT|C7676|NCI|Adenocarcinoma in Adenomatous Polyp|8210/3
C1321861|T191|AB|X77nK|RCD|Adenoca in adenomatous polyp|8210/3
C1321861|T191|AB|X77nK|RCD|Adenoca in polypoid adenoma|8210/3
C1321861|T191|SY|X77nK|RCD|Adenocarcinoma in a polyp|8210/3
C1321861|T191|PT|X77nK|RCD|Adenocarcinoma in adenomatous polyp|8210/3
C1321861|T191|SY|X77nK|RCD|Adenocarcinoma in polypoid adenoma|8210/3
C1321861|T191|SY|X77nK|RCD|Carcinoma in adenomatous polyp|8210/3
C1321861|T191|SY|43233001|SNOMEDCT_US|Adenocarcinoma in a polyp|8210/3
C1321861|T191|IS|43233001|SNOMEDCT_US|Adenocarcinoma in a polyp, NOS|8210/3
C1321861|T191|PT|29421000119105|SNOMEDCT_US|Adenocarcinoma in adenomatous polyp|8210/3
C1321861|T191|PT|43233001|SNOMEDCT_US|Adenocarcinoma in adenomatous polyp|8210/3
C1321861|T191|SY|43233001|SNOMEDCT_US|Adenocarcinoma in polypoid adenoma|8210/3
C1321861|T191|SY|43233001|SNOMEDCT_US|Carcinoma in adenomatous polyp|8210/3
C0334292|T191|PT|0049870|CCPSS|ADENOMA TUBULAR|8211/0
C0334292|T191|SY|0000029953|CHV|adenoma tubular|8211/0
C0334292|T191|SY|0000029953|CHV|adenomas tubular|8211/0
C0334292|T191|PT|0000029953|CHV|tubular adenoma|8211/0
C0334292|T191|LA|LA15387-6|LNC|Tubular adenoma|8211/0
C0334292|T191|LA|LA26485-5|LNC|Tubular adenoma, NOS|8211/0
C0334292|T191|PT|C4133|NCI|Tubular Adenoma|8211/0
C0334292|T191|PT|C4133|NCI_CDISC|ADENOMA, TUBULAR CELL, BENIGN|8211/0
C0334292|T191|PT|Xa98X|RCD|Tubular adenoma|8211/0
C0334292|T191|OP|BB5M0|RCDSY|Tubular adenoma NOS|8211/0
C0334292|T191|PT|444408007|SNOMEDCT_US|Tubular adenoma|8211/0
C0334292|T191|SY|19665009|SNOMEDCT_US|Tubular adenoma|8211/0
C2733364|T191|PT|443897009|SNOMEDCT_US|Tubular adenoma - category|8211/0
C0334292|T191|PT|19665009|SNOMEDCT_US|Tubular adenoma, no ICD-O subtype|8211/0
C0334292|T191|SY|19665009|SNOMEDCT_US|Tubular adenoma, no International Classification of Diseases for Oncology subtype|8211/0
C0334292|T191|IS|19665009|SNOMEDCT_US|Tubular adenoma, NOS|8211/0
C0205645|T191|SY|0000020665|CHV|carcinoma tubular|8211/3
C0205645|T191|SY|0000020665|CHV|tubular adenocarcinoma|8211/3
C0205645|T191|PT|0000020665|CHV|tubular carcinoma|8211/3
C0205645|T191|SY|0000020665|CHV|tubular carcinomas|8211/3
C0205645|T191|LA|LA26094-5|LNC|Tubular adenocarcinoma|8211/3
C0205645|T191|PT|271474|MEDCIN|tubular adenocarcinoma|8211/3
C0205645|T191|PEP|D000230|MSH|Adenocarcinoma, Tubular|8211/3
C0205645|T191|PM|D000230|MSH|Adenocarcinomas, Tubular|8211/3
C0205645|T191|ET|D000230|MSH|Carcinoma, Tubular|8211/3
C0205645|T191|PM|D000230|MSH|Carcinomas, Tubular|8211/3
C0205645|T191|PM|D000230|MSH|Tubular Adenocarcinoma|8211/3
C0205645|T191|PM|D000230|MSH|Tubular Adenocarcinomas|8211/3
C0205645|T191|PM|D000230|MSH|Tubular Carcinoma|8211/3
C0205645|T191|PM|D000230|MSH|Tubular Carcinomas|8211/3
C0205645|T191|PN|NOCODE|MTH|Adenocarcinoma, Tubular|8211/3
C0205645|T191|PT|C65192|NCI|Tubular Adenocarcinoma|8211/3
C0205645|T191|PT|C65192|NCI_CDISC|CARCINOMA, TUBULAR CELL, MALIGNANT|8211/3
C0205645|T191|PT|BB5M1|RCD|Tubular adenocarcinoma|8211/3
C0205645|T191|SY|BB5M1|RCD|Tubular carcinoma|8211/3
C0205645|T191|PT|4631006|SNOMEDCT_US|Tubular adenocarcinoma|8211/3
C0205645|T191|SY|4631006|SNOMEDCT_US|Tubular carcinoma|8211/3
C1266024|T191|PN|NOCODE|MTH|Flat adenoma|8212/0
C1266024|T191|PT|C65193|NCI|Flat Adenoma|8212/0
C1266024|T191|PT|128652009|SNOMEDCT_US|Flat adenoma|8212/0
C1266025|T191|SY|0000056677|CHV|adenomas serrated|8213/0
C1266025|T191|PT|0000056677|CHV|serrated adenoma|8213/0
C2732618|T191|LA|LA27155-3|LNC|Sessile serrated adenoma|8213/0
C2732618|T191|LA|LA26490-5|LNC|Sessile serrated adenoma/polyp|8213/0
C1266025|T191|LA|LA26492-1|LNC|Traditional serrated adenoma|8213/0
C2732618|T191|PN|NOCODE|MTH|Sessile Serrated Adenoma/Polyp|8213/0
C1266025|T191|PN|NOCODE|MTH|Traditional Serrated Adenoma|8213/0
C1266025|T191|SY|C38458|NCI|Serrated Adenoma|8213/0
C2732618|T191|SY|C96414|NCI|Serrated Adenoma Type I|8213/0
C1266025|T191|SY|C38458|NCI|Serrated Adenoma Type II|8213/0
C2732618|T191|SY|C96414|NCI|Serrated Polyp with Abnormal Proliferation|8213/0
C2732618|T191|SY|C96414|NCI|Sessile Serrated Adenoma|8213/0
C2732618|T191|PT|C96414|NCI|Sessile Serrated Adenoma/Polyp|8213/0
C2732618|T191|SY|C96414|NCI|Sessile Serrated Polyp|8213/0
C2732618|T191|SY|C96414|NCI|Sessile Serrated Polyp/Adenoma|8213/0
C2732618|T191|AB|C96414|NCI|SSA|8213/0
C2732618|T191|AB|C96414|NCI|SSA/P|8213/0
C2732618|T191|AB|C96414|NCI|SSP|8213/0
C1266025|T191|PT|C38458|NCI|Traditional Serrated Adenoma|8213/0
C1266025|T191|AB|C38458|NCI|TSA|8213/0
C1266025|T191|SY|128653004|SNOMEDCT_US|Mixed adenomatous and hyperplastic polyp|8213/0
C1266025|T191|PT|128653004|SNOMEDCT_US|Serrated adenoma|8213/0
C2732618|T191|PT|443157008|SNOMEDCT_US|Sessile serrated adenoma|8213/0
C5190874|T191|PT|783210009|SNOMEDCT_US|Sessile serrated adenoma with dysplasia|8213/0
C2732618|T191|SY|443157008|SNOMEDCT_US|Sessile serrated polyp|8213/0
C1266025|T191|PT|443734007|SNOMEDCT_US|Traditional serrated adenoma|8213/0
C3838988|T191|PT|703843001|SNOMEDCT_US|Traditional sessile serrated adenoma|8213/0
C3472623|T191|LA|LA26498-8|LNC|Serrated adenocarcinoma|8213/3
C3272809|T191|PT|C96485|NCI|Colorectal Serrated Adenocarcinoma|8213/3
C3472623|T191|PT|450948005|SNOMEDCT_US|Serrated adenocarcinoma|8213/3
C1266026|T191|PT|C65194|NCI|Gastric Parietal Cell Adenocarcinoma|8214/3
C1266026|T191|SY|C65194|NCI|Parietal Cell Adenocarcinoma|8214/3
C1266026|T191|SY|128654005|SNOMEDCT_US|Parietal cell adenocarcinoma|8214/3
C1266026|T191|PT|128654005|SNOMEDCT_US|Parietal cell carcinoma|8214/3
C1266027|T191|PT|39205|MEDCIN|adenocarcinoma of anal glands|8215/3
C1266027|T191|SY|C5609|NCI|Adenocarcinoma of Anal Gland|8215/3
C1266027|T191|SY|C5609|NCI|Adenocarcinoma of the Anal Gland|8215/3
C1266027|T191|PT|C5609|NCI|Anal Glands Adenocarcinoma|8215/3
C1266027|T191|SY|128655006|SNOMEDCT_US|Adenocarcinoma of anal ducts|8215/3
C1266027|T191|PT|128655006|SNOMEDCT_US|Adenocarcinoma of anal glands|8215/3
C0032580|T191|PT|0011401|CCPSS|COLON NOS POLYPOSIS|8220/0
C0032580|T191|SY|0000009935|CHV|adenomatous coli polyposis|8220/0
C0032580|T191|SY|0000009935|CHV|adenomatous polyposis|8220/0
C0032580|T191|SY|0000009935|CHV|adenomatous polyposis coli|8220/0
C0032580|T191|SY|0000009935|CHV|familial adenomatous polyposis|8220/0
C0032580|T191|SY|0000009935|CHV|familial intestinal polyposis|8220/0
C0032580|T191|SY|0000009935|CHV|familial polyposis|8220/0
C0032580|T191|SY|0000009935|CHV|familial polyposis coli|8220/0
C0032580|T191|SY|0000009935|CHV|familial polyposis syndrome|8220/0
C0032580|T191|PT|0000009935|CHV|fap|8220/0
C0032580|T191|SY|0000009935|CHV|polyposis coli|8220/0
C0032580|T191|SY|0000009935|CHV|polyposis familial|8220/0
C0032580|T191|PT|U000281|COSTAR|FAMILIAL POLYPOSIS|8220/0
C0032580|T191|ET|4005-0002|CSP|familial adenomatous polyposis|8220/0
C0032580|T191|ET|4006-0027|CSP|familial adenomatous polyposis|8220/0
C0032580|T191|ET|2010-0350|CSP|familial polyposis coli|8220/0
C0032580|T191|DI|U000383|DXP|COLON, POLYPOSIS, FAMILIAL ADENOMATOUS|8220/0
C0032580|T191|PT|MTHU017127|ICPC2ICD10ENG|colon; polyposis coli|8220/0
C0032580|T191|PT|MTHU027706|ICPC2ICD10ENG|familial; polyposis|8220/0
C0032580|T191|PT|MTHU061091|ICPC2ICD10ENG|polyposis; colon|8220/0
C0032580|T191|PT|MTHU061092|ICPC2ICD10ENG|polyposis; familial|8220/0
C0032580|T191|PT|D78004|ICPC2P|Polyposis Coli|8220/0
C0032580|T191|PTN|D78004|ICPC2P|Polyposis Coli|8220/0
C0032580|T191|PT|10056981|MDR|Adenomatous polyposis coli|8220/0
C0032580|T191|LLT|10056981|MDR|Adenomatous polyposis coli|8220/0
C0032580|T191|LLT|10059327|MDR|Familial adenomatous polyposis|8220/0
C0032580|T191|LLT|10057848|MDR|Familial polyposis|8220/0
C0032580|T191|LLT|10036135|MDR|Polyposis coli|8220/0
C0032580|T191|SY|312779|MEDCIN|adenomatous polyposis coli|8220/0
C0032580|T191|PT|312779|MEDCIN|adenomatous polyposis coli of large intestine|8220/0
C0032580|T191|PM|D011125|MSH|Adenomatous Polyposes, Familial|8220/0
C0032580|T191|MH|D011125|MSH|Adenomatous Polyposis Coli|8220/0
C0032580|T191|ET|D011125|MSH|Adenomatous Polyposis Coli, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Adenomatous Polyposis Colus|8220/0
C0032580|T191|ET|D011125|MSH|Adenomatous Polyposis of the Colon|8220/0
C0032580|T191|PM|D011125|MSH|Adenomatous Polyposis, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Coli, Adenomatous Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Coli, Familial Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Coli, Hereditary Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Coli, Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Colus, Adenomatous Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Colus, Familial Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Colus, Hereditary Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Colus, Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Familial Adenomatous Polyposes|8220/0
C0032580|T191|ET|D011125|MSH|Familial Adenomatous Polyposis|8220/0
C0032580|T191|ET|D011125|MSH|Familial Adenomatous Polyposis Coli|8220/0
C0032580|T191|ET|D011125|MSH|Familial Adenomatous Polyposis of the Colon|8220/0
C0032580|T191|PM|D011125|MSH|Familial Multiple Polyposes|8220/0
C0032580|T191|ET|D011125|MSH|Familial Multiple Polyposi|8220/0
C0032580|T191|ET|D011125|MSH|Familial Multiple Polyposis|8220/0
C0032580|T191|ET|D011125|MSH|Familial Multiple Polyposis Syndrome|8220/0
C0032580|T191|PM|D011125|MSH|Familial Multiple Polyposus|8220/0
C0032580|T191|ET|D011125|MSH|Familial Polyposis Coli|8220/0
C0032580|T191|PM|D011125|MSH|Familial Polyposis Colus|8220/0
C0032580|T191|ET|D011125|MSH|Familial Polyposis of the Colon|8220/0
C0032580|T191|ET|D011125|MSH|Familial Polyposis Syndrome|8220/0
C0032580|T191|PM|D011125|MSH|Familial Polyposis Syndromes|8220/0
C0032580|T191|ET|D011125|MSH|Hereditary Polyposis Coli|8220/0
C0032580|T191|PM|D011125|MSH|Hereditary Polyposis Colus|8220/0
C0032580|T191|PM|D011125|MSH|Multiple Polyposes, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Multiple Polyposi, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Multiple Polyposis, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Multiple Polyposus, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Myh Associated Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Myh-Associated Polyposes|8220/0
C0032580|T191|ET|D011125|MSH|Myh-Associated Polyposis|8220/0
C0032580|T191|PM|D011125|MSH|Polyposes, Familial Adenomatous|8220/0
C0032580|T191|PM|D011125|MSH|Polyposes, Familial Multiple|8220/0
C0032580|T191|PM|D011125|MSH|Polyposes, Myh-Associated|8220/0
C0032580|T191|PM|D011125|MSH|Polyposi, Familial Multiple|8220/0
C0032580|T191|ET|D011125|MSH|Polyposis Coli|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis Coli, Adenomatous|8220/0
C0032580|T191|ET|D011125|MSH|Polyposis Coli, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis Coli, Hereditary|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis Colus|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis Colus, Adenomatous|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis Colus, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis Colus, Hereditary|8220/0
C0032580|T191|ET|D011125|MSH|Polyposis Syndrome, Familial|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis, Familial Adenomatous|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis, Familial Multiple|8220/0
C0032580|T191|PM|D011125|MSH|Polyposis, Myh-Associated|8220/0
C0032580|T191|PM|D011125|MSH|Polyposus, Familial Multiple|8220/0
C0032580|T191|PN|NOCODE|MTH|Adenomatous Polyposis Coli|8220/0
C0032580|T191|SY|C3339|NCI|Adenomatous Polyposis Coli|8220/0
C0032580|T191|SY|C3339|NCI|APC - Adenomatous Polyposis Coli|8220/0
C0032580|T191|PT|C3339|NCI|Familial Adenomatous Polyposis|8220/0
C0032580|T191|SY|C3339|NCI|Familial Adenomatous Polyposis Coli|8220/0
C0032580|T191|SY|C3339|NCI|Familial Adenomatous Polyposis Syndrome|8220/0
C0032580|T191|AB|C3339|NCI|FAP|8220/0
C0032580|T191|SY|C3339|NCI|Hereditary Adenomatous Polyposis Coli|8220/0
C0032580|T191|SY|C3339|NCI|Polyposis Coli|8220/0
C0032580|T191|DN|C3339|NCI_CTRP|Familial Adenomatous Polyposis|8220/0
C0032580|T191|PT|CDR0000045100|NCI_NCI-GLOSS|familial adenomatous polyposis|8220/0
C0032580|T191|PT|CDR0000045688|NCI_NCI-GLOSS|familial polyposis|8220/0
C0032580|T191|PT|CDR0000044777|NCI_NCI-GLOSS|FAP|8220/0
C0032580|T191|SY|CDR0000042839|PDQ|adenomatous polyposis coli|8220/0
C0032580|T191|SY|CDR0000042839|PDQ|APC - adenomatous polyposis coli|8220/0
C0032580|T191|PT|CDR0000042839|PDQ|familial adenomatous polyposis|8220/0
C0032580|T191|SY|CDR0000042839|PDQ|familial adenomatous polyposis coli|8220/0
C0032580|T191|SY|CDR0000042839|PDQ|familial adenomatous polyposis syndrome|8220/0
C0032580|T191|ACR|CDR0000042839|PDQ|FAP|8220/0
C0032580|T191|SY|CDR0000042839|PDQ|hereditary adenomatous polyposis coli|8220/0
C0032580|T191|PT|CDR0000725405|PDQ|MYH-associated polyposis|8220/0
C0032580|T191|SY|CDR0000042839|PDQ|polyposis coli|8220/0
C0032580|T191|SY|CDR0000042839|PDQ|polyposis, familial adenomatous|8220/0
C0032580|T191|SY|CDR0000725405|PDQ|polyposis, MYH-associated|8220/0
C0032580|T191|SY|XE2xj|RCD|Adenomatous polyposis|8220/0
C0032580|T191|PT|XE2xj|RCD|Adenomatous polyposis coli|8220/0
C0032580|T191|AB|XE2xj|RCD|APC - Adenoma polyposis coli|8220/0
C0032580|T191|SY|XE2xj|RCD|APC - Adenomatous polyposis coli|8220/0
C0032580|T191|SY|XE2xj|RCD|Familial adenomatous polyposis|8220/0
C0032580|T191|SY|XE2xj|RCD|Familial polyposis coli|8220/0
C0032580|T191|AB|XE2xj|RCD|FAP - Fam adenoma polyposis|8220/0
C0032580|T191|SY|XE2xj|RCD|FAP - Familial adenomatous polyposis|8220/0
C0032580|T191|SY|XE2xj|RCD|FPC - Familial polyposis coli|8220/0
C0032580|T191|SY|XE2xj|RCD|Polyposis coli|8220/0
C0032580|T191|PT|BB5N0|RCDSY|Adenomatous polyposis coli|8220/0
C0032580|T191|SY|BB5N0|RCDSY|Familial polyposis coli|8220/0
C0032580|T191|SY|72900001|SNOMEDCT_US|Adenomatous polyposis|8220/0
C0032580|T191|PT|70921007|SNOMEDCT_US|Adenomatous polyposis coli|8220/0
C0032580|T191|SY|72900001|SNOMEDCT_US|Adenomatous polyposis coli|8220/0
C0032580|T191|SY|72900001|SNOMEDCT_US|APC - Adenomatous polyposis coli|8220/0
C0032580|T191|SY|72900001|SNOMEDCT_US|Familial adenomatous polyposis|8220/0
C0032580|T191|PT|72900001|SNOMEDCT_US|Familial multiple polyposis syndrome|8220/0
C0032580|T191|SY|72900001|SNOMEDCT_US|Familial polyposis coli|8220/0
C0032580|T191|SY|70921007|SNOMEDCT_US|Familial polyposis coli|8220/0
C0032580|T191|SY|72900001|SNOMEDCT_US|FAP - Familial adenomatous polyposis|8220/0
C0032580|T191|SY|72900001|SNOMEDCT_US|FPC - Familial polyposis coli|8220/0
C0032580|T191|SY|423471004|SNOMEDCT_US|MAP - MYH associated polyposis|8220/0
C0032580|T191|PT|423471004|SNOMEDCT_US|MYH-associated polyposis|8220/0
C0032580|T191|OAS|188828009|SNOMEDCT_US|Polyposis coli|8220/0
C0032580|T191|OAS|269636003|SNOMEDCT_US|Polyposis coli|8220/0
C0032580|T191|SY|72900001|SNOMEDCT_US|Polyposis coli|8220/0
C0032580|T191|OAS|154609001|SNOMEDCT_US|Polyposis coli|8220/0
C0032580|T191|SY|70921007|SNOMEDCT_US|Polyposis coli|8220/0
C0334293|T191|PT|C4134|NCI|Adenocarcinoma in Adenomatous Polyposis Coli|8220/3
C0334293|T191|AB|BB5N1|RCD|Adenoca in adenom polypos coli|8220/3
C0334293|T191|PT|BB5N1|RCD|Adenocarcinoma in adenomatous polyposis coli|8220/3
C0334293|T191|PT|57513006|SNOMEDCT_US|Adenocarcinoma in adenomatous polyposis coli|8220/3
C0334294|T191|PT|0003345|CCPSS|POLYP ADENOMATOUS MULTIPLE|8221/0
C0334294|T191|PT|0000000718|CHV|adenomatosis|8221/0
C0334294|T191|PT|MTHU003464|ICPC2ICD10ENG|adenomatosis; unspecified site|8221/0
C0334294|T191|PT|C4135|NCI|Multiple Adenomatous Polyps|8221/0
C0334294|T191|PT|BB5N2|RCD|Multiple adenomatous polyps|8221/0
C0334294|T191|SY|70921007|SNOMEDCT_US|Adenomatosis|8221/0
C0334294|T191|IS|70921007|SNOMEDCT_US|Adenomatosis, NOS|8221/0
C0334294|T191|PT|6379007|SNOMEDCT_US|Multiple adenomatous polyps|8221/0
C0334295|T191|PT|C4136|NCI|Adenocarcinoma in Multiple Adenomatous Polyps|8221/3
C0334295|T191|AB|X77nN|RCD|Adenoca in mult adenom polyps|8221/3
C0334295|T191|PT|X77nN|RCD|Adenocarcinoma in multiple adenomatous polyps|8221/3
C0334295|T191|AB|X77nN|RCDSY|Adencarc multp adenom polyp|8221/3
C0334295|T191|OAP|189599005|SNOMEDCT_US|Adenocarcinoma in multiple adenomatous polyps|8221/3
C0334295|T191|OF|189599005|SNOMEDCT_US|Adenocarcinoma in multiple adenomatous polyps|8221/3
C0334295|T191|PT|47299001|SNOMEDCT_US|Adenocarcinoma in multiple adenomatous polyps|8221/3
C1266028|T191|SY|271391|MEDCIN|duct carcinoma in situ, solid type|8230/2
C1266028|T191|PT|271391|MEDCIN|solid type ductal carcinoma in situ|8230/2
C1880424|T191|PT|232267|MEDCIN|solid type ductal carcinoma in situ of breast|8230/2
C1880424|T191|PT|C66933|NCI|Ductal Breast Carcinoma In Situ, Solid Type|8230/2
C1880424|T191|SY|C66933|NCI|Ductal Breast Carcinoma in Situ, Solid Type|8230/2
C1266028|T191|PT|128880009|SNOMEDCT_US|Ductal carcinoma in situ, solid type|8230/2
C1266028|T191|SY|128880009|SNOMEDCT_US|Intraductal carcinoma, solid type|8230/2
C0334296|T191|PT|271427|MEDCIN|solid carcinoma|8230/3
C0334296|T191|PT|C4137|NCI|Solid Carcinoma|8230/3
C0334296|T191|PT|C4137|NCI_CPTAC|Solid Carcinoma|8230/3
C0334296|T191|PT|Xa98Y|RCD|Solid carcinoma|8230/3
C0334296|T191|OP|BB5P.|RCDSY|Solid carcinoma NOS|8230/3
C0334296|T191|SY|81920005|SNOMEDCT_US|Solid adenocarcinoma with mucin formation|8230/3
C0334296|T191|PT|81920005|SNOMEDCT_US|Solid carcinoma|8230/3
C0334296|T191|SY|81920005|SNOMEDCT_US|Solid carcinoma with mucin formation|8230/3
C0334296|T191|IS|81920005|SNOMEDCT_US|Solid carcinoma, NOS|8230/3
C0334297|T191|PT|271428|MEDCIN|carcinoma simplex|8231/3
C0334297|T191|OP|C65195|NCI|Carcinoma Simplex|8231/3
C0334297|T191|PT|C65195|NCI|Carcinoma Simplex|8231/3
C0334297|T191|PT|BB5Q.|RCD|Carcinoma simplex|8231/3
C0334297|T191|PT|45881000|SNOMEDCT_US|Carcinoma simplex|8231/3
C0334297|T191|SY|403939009|SNOMEDCT_US|Carcinoma simplex|8231/3
C0334298|T191|SY|0000029954|CHV|appendix carcinoid|8240/1
C0334298|T191|SY|0000029954|CHV|appendix carcinoid tumors|8240/1
C0334298|T191|SY|0000029954|CHV|appendix carcinoids|8240/1
C0334298|T191|SY|0000029954|CHV|carcinoid appendix|8240/1
C0334298|T191|SY|0000029954|CHV|carcinoid of appendix|8240/1
C0334298|T191|SY|0000029954|CHV|carcinoid tumor appendix|8240/1
C0334298|T191|PT|0000029954|CHV|carcinoid tumor of appendix|8240/1
C0600176|T191|ET|2010-0179|CSP|argentaffinoma|8240/1
C0600176|T191|ET|1025-5693|CSP|argentaffinoma|8240/1
C0334298|T191|PT|MTHU007630|ICPC2ICD10ENG|appendix; carcinoid|8240/1
C0334298|T191|PT|MTHU014699|ICPC2ICD10ENG|carcinoid; appendix|8240/1
C0334298|T191|MTH_LLT|10003015|MDR|Appendix carcinoid tumor|8240/1
C0334298|T191|LLT|10003015|MDR|Appendix carcinoid tumour|8240/1
C0600176|T191|LLT|10003089|MDR|Argentaffinoma|8240/1
C0334298|T191|LLT|10007272|MDR|Carcinoid tumor of the appendix|8240/1
C0334298|T191|MTH_PT|10007277|MDR|Carcinoid tumor of the appendix|8240/1
C0334298|T191|LLT|10007277|MDR|Carcinoid tumour of the appendix|8240/1
C0334298|T191|PT|10007277|MDR|Carcinoid tumour of the appendix|8240/1
C0600176|T191|PEP|D002276|MSH|Argentaffinoma|8240/1
C0600176|T191|PM|D002276|MSH|Argentaffinomas|8240/1
C0600176|T191|PN|NOCODE|MTH|Argentaffinoma|8240/1
C0334298|T191|PN|NOCODE|MTH|Carcinoid tumor of appendix|8240/1
C0334298|T191|SY|C4138|NCI|Appendiceal Carcinoid Tumor|8240/1
C0334298|T191|SY|C4138|NCI|Appendix Carcinoid Tumor|8240/1
C0334298|T191|SY|C4138|NCI|Appendix NET G1|8240/1
C0334298|T191|PT|C4138|NCI|Appendix Neuroendocrine Tumor G1|8240/1
C0334298|T191|SY|C4138|NCI|Carcinoid Tumor of Appendix|8240/1
C0334298|T191|SY|C4138|NCI|Carcinoid Tumor of the Appendix|8240/1
C0600176|T191|OP|C65196|NCI|Carcinoid Tumor of Uncertain Malignant Potential|8240/1
C0600176|T191|PT|C65196|NCI|Carcinoid Tumor of Uncertain Malignant Potential|8240/1
C0334298|T191|PT|C4138|NCI_CPTAC|Appendix Neuroendocrine Tumor G1|8240/1
C0600176|T191|SY|XM1FG|RCD|Argentaffinoma|8240/1
C0334298|T191|SY|X77nS|RCD|Carcinoid of appendix|8240/1
C0600176|T191|PT|XM1FG|RCD|Carcinoid tumour - argentaffin|8240/1
C0334298|T191|PT|X77nS|RCD|Carcinoid tumour of appendix|8240/1
C0600176|T191|PT|XM1FG|RCDAE|Carcinoid tumor - argentaffin|8240/1
C0334298|T191|PT|X77nS|RCDAE|Carcinoid tumor of appendix|8240/1
C0600176|T191|SY|XM1FG|RCDSA|Carcinoid tumor, argentaffin, NOS|8240/1
C0600176|T191|SY|XM1FG|RCDSY|Carcinoid tumour, argentaffin, NOS|8240/1
C0600176|T191|AB|XM1FG|RCDSY|Carcinoid, argentaffin NOS|8240/1
C0600176|T191|SY|274904007|SNOMEDCT_US|Argentaffinoma|8240/1
C0600176|T191|IS|15005003|SNOMEDCT_US|Argentaffinoma, NOS|8240/1
C0334298|T191|SY|253002004|SNOMEDCT_US|Carcinoid of appendix|8240/1
C0600176|T191|OAP|189610004|SNOMEDCT_US|Carcinoid tumor - argentaffin|8240/1
C0600176|T191|PT|274904007|SNOMEDCT_US|Carcinoid tumor - argentaffin|8240/1
C0334298|T191|PT|253002004|SNOMEDCT_US|Carcinoid tumor of appendix|8240/1
C0334298|T191|PT|22228003|SNOMEDCT_US|Carcinoid tumor of uncertain malignant potential|8240/1
C0334298|T191|SY|22228003|SNOMEDCT_US|Carcinoid tumor, argentaffin|8240/1
C0600176|T191|OAP|15005003|SNOMEDCT_US|Carcinoid tumor, argentaffin|8240/1
C0600176|T191|IS|15005003|SNOMEDCT_US|Carcinoid tumor, argentaffin -RETIRED-|8240/1
C0600176|T191|OF|15005003|SNOMEDCT_US|Carcinoid tumor, argentaffin -RETIRED-|8240/1
C0600176|T191|IS|15005003|SNOMEDCT_US|Carcinoid tumor, argentaffin, NOS|8240/1
C0334298|T191|IS|22228003|SNOMEDCT_US|Carcinoid tumor, NOS, of appendix|8240/1
C0334298|T191|SY|22228003|SNOMEDCT_US|Carcinoid tumor, of appendix|8240/1
C0600176|T191|OAP|189610004|SNOMEDCT_US|Carcinoid tumour - argentaffin|8240/1
C0600176|T191|OF|189610004|SNOMEDCT_US|Carcinoid tumour - argentaffin|8240/1
C0600176|T191|PTGB|274904007|SNOMEDCT_US|Carcinoid tumour - argentaffin|8240/1
C0334298|T191|PTGB|253002004|SNOMEDCT_US|Carcinoid tumour of appendix|8240/1
C0334298|T191|PTGB|22228003|SNOMEDCT_US|Carcinoid tumour of uncertain malignant potential|8240/1
C0334298|T191|SYGB|22228003|SNOMEDCT_US|Carcinoid tumour, argentaffin|8240/1
C0600176|T191|OAP|15005003|SNOMEDCT_US|Carcinoid tumour, argentaffin|8240/1
C0600176|T191|IS|15005003|SNOMEDCT_US|Carcinoid tumour, argentaffin -RETIRED-|8240/1
C0334298|T191|SYGB|22228003|SNOMEDCT_US|Carcinoid tumour, of appendix|8240/1
C0334298|T191|IS|22228003|SNOMEDCT_US|Carcinoid, NOS, of appendix|8240/1
C0334298|T191|SY|22228003|SNOMEDCT_US|Carcinoid, of appendix|8240/1
C0007095|T191|PT|0050269|CCPSS|CARCINOID TUMOR|8240/3
C0007095|T191|SY|0000002415|CHV|carcinoid|8240/3
C0220620|T191|SY|0000021166|CHV|carcinoid gastrointestinal tumors|8240/3
C0007095|T191|PT|0000002415|CHV|carcinoid tumor|8240/3
C0007095|T191|SY|0000002415|CHV|carcinoid tumors|8240/3
C0007095|T191|SY|0000002415|CHV|carcinoid tumour|8240/3
C0007095|T191|SY|0000002415|CHV|carcinoid tumours|8240/3
C0007095|T191|SY|0000002415|CHV|carcinoids|8240/3
C0220620|T191|PT|0000021166|CHV|gastrointestinal carcinoid tumor|8240/3
C0007095|T191|PT|U000102|COSTAR|CARCINOID|8240/3
C0007095|T191|SY|HP:0100570|HPO|Carcinoid|8240/3
C0007095|T191|PT|HP:0100570|HPO|Carcinoid tumor|8240/3
C0007095|T191|ET|HP:0100570|HPO|Carcinoid tumors|8240/3
C0007095|T191|ET|D3A.00|ICD10CM|Carcinoid tumor NOS|8240/3
C0007095|T191|PT|sh85020159|LCH_NW|Carcinoid|8240/3
C0007095|T191|LLT|10007271|MDR|Carcinoid tumor|8240/3
C0007095|T191|MTH_PT|10007275|MDR|Carcinoid tumor|8240/3
C0007095|T191|MTH_LLT|10007276|MDR|Carcinoid tumor NOS|8240/3
C0220620|T191|LLT|10062391|MDR|Carcinoid tumor of the gastrointestinal tract|8240/3
C0220620|T191|MTH_PT|10007279|MDR|Carcinoid tumor of the gastrointestinal tract|8240/3
C0007095|T191|MTH_HT|10007283|MDR|Carcinoid tumors|8240/3
C0007095|T191|LLT|10007275|MDR|Carcinoid tumour|8240/3
C0007095|T191|PT|10007275|MDR|Carcinoid tumour|8240/3
C0007095|T191|LLT|10007276|MDR|Carcinoid tumour NOS|8240/3
C0220620|T191|PT|10007279|MDR|Carcinoid tumour of the gastrointestinal tract|8240/3
C0220620|T191|LLT|10007279|MDR|Carcinoid tumour of the gastrointestinal tract|8240/3
C0007095|T191|HT|10007283|MDR|Carcinoid tumours|8240/3
C0220620|T191|LLT|10062426|MDR|Gastrointestinal carcinoid tumor|8240/3
C0220620|T191|LLT|10017939|MDR|Gastrointestinal carcinoid tumour|8240/3
C0007095|T191|PT|1277|MEDLINEPLUS|Carcinoid Tumors|8240/3
C0007095|T191|ET|D002276|MSH|Carcinoid|8240/3
C0007095|T191|MH|D002276|MSH|Carcinoid Tumor|8240/3
C0007095|T191|PM|D002276|MSH|Carcinoid Tumors|8240/3
C0007095|T191|PM|D002276|MSH|Carcinoids|8240/3
C0007095|T191|PM|D002276|MSH|Tumor, Carcinoid|8240/3
C0007095|T191|PM|D002276|MSH|Tumors, Carcinoid|8240/3
C0007095|T191|PN|NOCODE|MTH|Carcinoid Tumor|8240/3
C0334299|T191|PN|NOCODE|MTH|Carcinoid tumor no ICD-O subtype|8240/3
C0220620|T191|PN|NOCODE|MTH|Gastrointestinal Carcinoid Tumor|8240/3
C0007095|T191|ET|209.60|MTHICD9|Carcinoid tumor NOS|8240/3
C0007095|T191|SY|C2915|NCI|Carcinoid|8240/3
C0007095|T191|SY|TCGA|NCI|Carcinoid Tumor|8240/3
C0007095|T191|PT|C2915|NCI|Carcinoid Tumor|8240/3
C0220620|T191|SY|C7709|NCI|Carcinoid Tumor of Digestive System|8240/3
C0220620|T191|SY|C7709|NCI|Carcinoid Tumor of Gastrointestinal System|8240/3
C0220620|T191|SY|C7709|NCI|Carcinoid Tumor of GI System|8240/3
C0220620|T191|SY|C7709|NCI|Carcinoid Tumor of the Digestive System|8240/3
C0220620|T191|SY|C7709|NCI|Carcinoid Tumor of the Gastrointestinal System|8240/3
C0220620|T191|SY|C7709|NCI|Carcinoid Tumor of the GI System|8240/3
C0220620|T191|SY|C7709|NCI|Digestive Carcinoid Tumor|8240/3
C0220620|T191|SY|C7709|NCI|Digestive System Carcinoid Tumor|8240/3
C0220620|T191|PT|C7709|NCI|Digestive System Neuroendocrine Tumor G1|8240/3
C0220620|T191|SY|C7709|NCI|Gastrointestinal Carcinoid Tumor|8240/3
C0220620|T191|SY|C7709|NCI|Gastrointestinal NET G1|8240/3
C0220620|T191|SY|C7709|NCI|Gastrointestinal Neuroendocrine Tumor G1|8240/3
C0220620|T191|SY|C7709|NCI|Gastrointestinal System Carcinoid Tumor|8240/3
C0220620|T191|AB|C7709|NCI|GCT|8240/3
C0220620|T191|SY|C7709|NCI|GI Carcinoid Tumor|8240/3
C1266147|T191|OP|C35727|NCI|Grade I Neuroendocrine Carcinoma|8240/3
C1266147|T191|PT|C35727|NCI|Grade I Neuroendocrine Carcinoma|8240/3
C0007095|T191|PT|C2915|NCI_CPTAC|Carcinoid Tumor|8240/3
C0007095|T191|PT|10007276|NCI_CTEP-SDC|Carcinoid tumor|8240/3
C0007095|T191|DN|C2915|NCI_CTRP|Carcinoid Tumor|8240/3
C0220620|T191|DN|C7709|NCI_CTRP|Gastrointestinal Neuroendocrine Tumor G1|8240/3
C0007095|T191|PT|CDR0000044233|NCI_NCI-GLOSS|carcinoid|8240/3
C0220620|T191|PT|CDR0000446559|NCI_NCI-GLOSS|gastrointestinal carcinoid tumor|8240/3
C0007095|T191|PT|CDR0000665198|PDQ|carcinoid tumor|8240/3
C0220620|T191|SY|CDR0000038092|PDQ|carcinoid tumor, gastrointestinal|8240/3
C0220620|T191|ET|CDR0000038092|PDQ|Gastrointestinal carcinoid tumor|8240/3
C0220620|T191|PSC|CDR0000038092|PDQ|gastrointestinal carcinoid tumor|8240/3
C0220620|T191|SY|CDR0000038092|PDQ|GCT|8240/3
C0220620|T191|SY|CDR0000038092|PDQ|GI carcinoid tumor|8240/3
C0007095|T191|SY|BB5R.|RCD|Carcinoid|8240/3
C0007095|T191|SY|BB5R.|RCD|Carcinoid tumour|8240/3
C0007095|T191|PT|BB5R.|RCD|Carcinoid tumour - morphology|8240/3
C0007095|T191|SY|BB5R.|RCDAE|Carcinoid tumor|8240/3
C0007095|T191|PT|BB5R.|RCDAE|Carcinoid tumor - morphology|8240/3
C0007095|T191|OP|BB5R0|RCDSA|Carcinoid tumor NOS|8240/3
C0007095|T191|SY|BB5R.|RCDSA|Carcinoid tumors|8240/3
C0007095|T191|OP|BB5Rz|RCDSA|Carcinoid tumors NOS|8240/3
C0007095|T191|OP|BB5R0|RCDSY|Carcinoid tumour NOS|8240/3
C0007095|T191|SY|BB5R.|RCDSY|Carcinoid tumours|8240/3
C0007095|T191|OP|BB5Rz|RCDSY|Carcinoid tumours NOS|8240/3
C0007095|T191|SY|189607006|SNOMEDCT_US|Carcinoid|8240/3
C0334299|T191|SY|81622000|SNOMEDCT_US|Carcinoid|8240/3
C0334299|T191|PT|81622000|SNOMEDCT_US|Carcinoid tumor|8240/3
C0007095|T191|PT|443492008|SNOMEDCT_US|Carcinoid tumor|8240/3
C0007095|T191|SY|189607006|SNOMEDCT_US|Carcinoid tumor|8240/3
C0007095|T191|PT|189607006|SNOMEDCT_US|Carcinoid tumor - morphology|8240/3
C0334299|T191|SY|81622000|SNOMEDCT_US|Carcinoid tumor no ICD-O subtype|8240/3
C0334299|T191|SY|81622000|SNOMEDCT_US|Carcinoid tumor no International Classification of Diseases for Oncology subtype|8240/3
C0220620|T191|PT|428701004|SNOMEDCT_US|Carcinoid tumor of gastrointestinal tract|8240/3
C0334299|T191|PTGB|81622000|SNOMEDCT_US|Carcinoid tumour|8240/3
C0007095|T191|PTGB|443492008|SNOMEDCT_US|Carcinoid tumour|8240/3
C0007095|T191|SYGB|189607006|SNOMEDCT_US|Carcinoid tumour|8240/3
C0007095|T191|PTGB|189607006|SNOMEDCT_US|Carcinoid tumour - morphology|8240/3
C0334299|T191|SYGB|81622000|SNOMEDCT_US|Carcinoid tumour no ICD-O subtype|8240/3
C0220620|T191|PTGB|428701004|SNOMEDCT_US|Carcinoid tumour of gastrointestinal tract|8240/3
C1266147|T191|SY|127572005|SNOMEDCT_US|Grade 1 neuroendocrine carcinoma|8240/3
C1266147|T191|SY|127572005|SNOMEDCT_US|Neuroendocrine carcinoma, grade 1|8240/3
C1266147|T191|PT|127572005|SNOMEDCT_US|Neuroendocrine tumor grade 1|8240/3
C1266147|T191|PTGB|127572005|SNOMEDCT_US|Neuroendocrine tumour grade 1|8240/3
C0334299|T191|SY|81622000|SNOMEDCT_US|Typical carcinoid|8240/3
C1266147|T191|SY|127572005|SNOMEDCT_US|Well-differentiated neuroendocrine carcinoma|8240/3
C0007095|T191|PT|0050269|CCPSS|CARCINOID TUMOR|8241/3
C0007095|T191|SY|0000002415|CHV|carcinoid|8241/3
C0007095|T191|PT|0000002415|CHV|carcinoid tumor|8241/3
C0007095|T191|SY|0000002415|CHV|carcinoid tumors|8241/3
C0007095|T191|SY|0000002415|CHV|carcinoid tumour|8241/3
C0007095|T191|SY|0000002415|CHV|carcinoid tumours|8241/3
C0007095|T191|SY|0000002415|CHV|carcinoids|8241/3
C0007095|T191|PT|U000102|COSTAR|CARCINOID|8241/3
C0007095|T191|SY|HP:0100570|HPO|Carcinoid|8241/3
C0007095|T191|PT|HP:0100570|HPO|Carcinoid tumor|8241/3
C0007095|T191|ET|HP:0100570|HPO|Carcinoid tumors|8241/3
C0007095|T191|ET|D3A.00|ICD10CM|Carcinoid tumor NOS|8241/3
C0007095|T191|PT|sh85020159|LCH_NW|Carcinoid|8241/3
C0007095|T191|LLT|10007271|MDR|Carcinoid tumor|8241/3
C0007095|T191|MTH_PT|10007275|MDR|Carcinoid tumor|8241/3
C0007095|T191|MTH_LLT|10007276|MDR|Carcinoid tumor NOS|8241/3
C0007095|T191|MTH_HT|10007283|MDR|Carcinoid tumors|8241/3
C0007095|T191|LLT|10007275|MDR|Carcinoid tumour|8241/3
C0007095|T191|PT|10007275|MDR|Carcinoid tumour|8241/3
C0007095|T191|LLT|10007276|MDR|Carcinoid tumour NOS|8241/3
C0007095|T191|HT|10007283|MDR|Carcinoid tumours|8241/3
C0334300|T191|SY|271482|MEDCIN|enterochromaffin cell carcinoid tumor|8241/3
C0334300|T191|PT|271482|MEDCIN|malignant enterochromaffin cell carcinoid tumor|8241/3
C0007095|T191|PT|1277|MEDLINEPLUS|Carcinoid Tumors|8241/3
C0007095|T191|ET|D002276|MSH|Carcinoid|8241/3
C0007095|T191|MH|D002276|MSH|Carcinoid Tumor|8241/3
C0007095|T191|PM|D002276|MSH|Carcinoid Tumors|8241/3
C0007095|T191|PM|D002276|MSH|Carcinoids|8241/3
C0007095|T191|PM|D002276|MSH|Tumor, Carcinoid|8241/3
C0007095|T191|PM|D002276|MSH|Tumors, Carcinoid|8241/3
C0007095|T191|PN|NOCODE|MTH|Carcinoid Tumor|8241/3
C0007095|T191|ET|209.60|MTHICD9|Carcinoid tumor NOS|8241/3
C0007095|T191|SY|C2915|NCI|Carcinoid|8241/3
C0007095|T191|SY|TCGA|NCI|Carcinoid Tumor|8241/3
C0007095|T191|PT|C2915|NCI|Carcinoid Tumor|8241/3
C0007095|T191|PT|C2915|NCI_CPTAC|Carcinoid Tumor|8241/3
C0007095|T191|PT|10007276|NCI_CTEP-SDC|Carcinoid tumor|8241/3
C0007095|T191|DN|C2915|NCI_CTRP|Carcinoid Tumor|8241/3
C0007095|T191|PT|CDR0000044233|NCI_NCI-GLOSS|carcinoid|8241/3
C0007095|T191|PT|CDR0000665198|PDQ|carcinoid tumor|8241/3
C0007095|T191|SY|BB5R.|RCD|Carcinoid|8241/3
C0007095|T191|SY|BB5R.|RCD|Carcinoid tumour|8241/3
C0007095|T191|PT|BB5R.|RCD|Carcinoid tumour - morphology|8241/3
C0334300|T191|AB|BB5R3|RCD|Malig carcinoid tum-argentaff|8241/3
C0334300|T191|SY|BB5R3|RCD|Malignant argentaffinoma|8241/3
C0334300|T191|SY|BB5R3|RCD|Malignant carcinoid tumour - argentaffin|8241/3
C0007095|T191|SY|BB5R.|RCDAE|Carcinoid tumor|8241/3
C0007095|T191|PT|BB5R.|RCDAE|Carcinoid tumor - morphology|8241/3
C0334300|T191|SY|BB5R3|RCDAE|Malignant carcinoid tumor - argentaffin|8241/3
C0007095|T191|OP|BB5R0|RCDSA|Carcinoid tumor NOS|8241/3
C0334300|T191|PT|BB5R3|RCDSA|Carcinoid tumor, argentaffin, malignant|8241/3
C0007095|T191|SY|BB5R.|RCDSA|Carcinoid tumors|8241/3
C0007095|T191|OP|BB5Rz|RCDSA|Carcinoid tumors NOS|8241/3
C0007095|T191|OP|BB5R0|RCDSY|Carcinoid tumour NOS|8241/3
C0334300|T191|PT|BB5R3|RCDSY|Carcinoid tumour, argentaffin, malignant|8241/3
C0007095|T191|SY|BB5R.|RCDSY|Carcinoid tumours|8241/3
C0007095|T191|OP|BB5Rz|RCDSY|Carcinoid tumours NOS|8241/3
C0334300|T191|AB|BB5R3|RCDSY|Carcinoid,argentaffin,malig|8241/3
C0334300|T191|SY|48554007|SNOMEDCT_US|Argentaffinoma, malignant|8241/3
C0007095|T191|SY|189607006|SNOMEDCT_US|Carcinoid|8241/3
C0007095|T191|PT|443492008|SNOMEDCT_US|Carcinoid tumor|8241/3
C0007095|T191|SY|189607006|SNOMEDCT_US|Carcinoid tumor|8241/3
C0007095|T191|PT|189607006|SNOMEDCT_US|Carcinoid tumor - morphology|8241/3
C0334300|T191|SY|48554007|SNOMEDCT_US|Carcinoid tumor, argentaffin, malignant|8241/3
C0007095|T191|PTGB|443492008|SNOMEDCT_US|Carcinoid tumour|8241/3
C0007095|T191|SYGB|189607006|SNOMEDCT_US|Carcinoid tumour|8241/3
C0007095|T191|PTGB|189607006|SNOMEDCT_US|Carcinoid tumour - morphology|8241/3
C0334300|T191|SYGB|48554007|SNOMEDCT_US|Carcinoid tumour, argentaffin, malignant|8241/3
C0334300|T191|SY|48554007|SNOMEDCT_US|EC cell carcinoid|8241/3
C0334300|T191|PT|48554007|SNOMEDCT_US|Enterochromaffin cell carcinoid|8241/3
C0334300|T191|SY|48554007|SNOMEDCT_US|Malignant argentaffinoma|8241/3
C0334300|T191|SY|48554007|SNOMEDCT_US|Malignant carcinoid tumor - argentaffin|8241/3
C0334300|T191|SYGB|48554007|SNOMEDCT_US|Malignant carcinoid tumour - argentaffin|8241/3
C0334300|T191|SY|48554007|SNOMEDCT_US|Serotonin producing carcinoid|8241/3
C1333401|T191|SY|C27252|NCI|ECL Cell NET G1|8242/1
C1333401|T191|SY|C27252|NCI|Enterochromaffin-Like Cell Carcinoid Tumor|8242/1
C1333401|T191|SY|C27252|NCI|Enterochromaffin-Like Cell NET G1|8242/1
C1333401|T191|SY|C27252|NCI|Enterochromaffin-Like Cell Neuroendocrine Tumor|8242/1
C1333401|T191|PT|C27252|NCI|Enterochromaffin-Like Cell Neuroendocrine Tumor G1|8242/1
C1266029|T191|SY|128656007|SNOMEDCT_US|ECL cell carcinoid|8242/1
C1266029|T191|PT|128656007|SNOMEDCT_US|Enterochromaffin-like cell carcinoid|8242/1
C1333401|T191|SY|C27252|NCI|ECL Cell NET G1|8242/3
C1333401|T191|SY|C27252|NCI|Enterochromaffin-Like Cell Carcinoid Tumor|8242/3
C1333401|T191|SY|C27252|NCI|Enterochromaffin-Like Cell NET G1|8242/3
C1333401|T191|SY|C27252|NCI|Enterochromaffin-Like Cell Neuroendocrine Tumor|8242/3
C1333401|T191|PT|C27252|NCI|Enterochromaffin-Like Cell Neuroendocrine Tumor G1|8242/3
C1266030|T191|SY|128657003|SNOMEDCT_US|ECL cell carcinoid, malignant|8242/3
C1266030|T191|PT|128657003|SNOMEDCT_US|Enterochromaffin-like cell tumor, malignant|8242/3
C1266030|T191|PTGB|128657003|SNOMEDCT_US|Enterochromaffin-like cell tumour, malignant|8242/3
C0205695|T191|PT|MTHU014700|ICPC2ICD10ENG|carcinoid; goblet cell|8243/3
C0205695|T191|PT|MTHU010082|ICPC2ICD10ENG|goblet cell; carcinoid|8243/3
C0205695|T191|PT|MTHU050456|ICPC2ICD10ENG|mucocarcinoid; tumor, unspecified site|8243/3
C0205695|T191|PT|MTHU077102|ICPC2ICD10ENG|tumor; mucocarcinoid, unspecified site|8243/3
C0205695|T191|PT|217269|MEDCIN|adenocarcinoid tumor of appendix|8243/3
C0205695|T191|PT|271484|MEDCIN|goblet cell carcinoid|8243/3
C0205695|T191|PT|217267|MEDCIN|goblet cell carcinoid of appendix|8243/3
C0205695|T191|SY|271484|MEDCIN|goblet cell carcinoid tumor|8243/3
C0205695|T191|PEP|D002276|MSH|Carcinoid, Goblet Cell|8243/3
C0205695|T191|PM|D002276|MSH|Carcinoids, Goblet Cell|8243/3
C0205695|T191|PM|D002276|MSH|Goblet Cell Carcinoid|8243/3
C0205695|T191|PM|D002276|MSH|Goblet Cell Carcinoids|8243/3
C0205695|T191|SY|C3689|NCI|Appendix Adenocarcinoid Tumor|8243/3
C0205695|T191|PT|C3689|NCI|Appendix Goblet Cell Carcinoid|8243/3
C0205695|T191|SY|C3689|NCI|Appendix Goblet Cell Carcinoid Tumor|8243/3
C0205695|T191|SY|C3689|NCI|Appendix Mixed Carcinoid-Adenocarcinoma|8243/3
C0205695|T191|SY|C3689|NCI|Goblet Cell Carcinoid Tumor|8243/3
C0205695|T191|SY|C3689|NCI|Mucinous Carcinoid Tumor|8243/3
C0205695|T191|PT|Xa98Z|RCD|Goblet cell carcinoid|8243/3
C0205695|T191|SY|Xa98Z|RCD|Mucinous carcinoid|8243/3
C0205695|T191|SY|Xa98Z|RCD|Mucocarcinoid tumour|8243/3
C0205695|T191|SY|Xa98Z|RCDAE|Mucocarcinoid tumor|8243/3
C0205695|T191|SY|Xa98Z|RCDSA|Mucocarcinoid tumor, malignant|8243/3
C0205695|T191|AB|Xa98Z|RCDSA|Mucocarcinoid tumor,malig.|8243/3
C0205695|T191|SY|Xa98Z|RCDSY|Mucocarcinoid tumour, malignant|8243/3
C0205695|T191|AB|Xa98Z|RCDSY|Mucocarcinoid tumour,malig.|8243/3
C0205695|T191|OF|189613002|SNOMEDCT_US|Goblet cell carcinoid|8243/3
C0205695|T191|PT|31396002|SNOMEDCT_US|Goblet cell carcinoid|8243/3
C0205695|T191|OAP|189613002|SNOMEDCT_US|Goblet cell carcinoid|8243/3
C0205695|T191|SY|31396002|SNOMEDCT_US|Mucinous carcinoid|8243/3
C0205695|T191|SY|31396002|SNOMEDCT_US|Mucocarcinoid tumor|8243/3
C0205695|T191|SY|31396002|SNOMEDCT_US|Mucocarcinoid tumor, malignant|8243/3
C0205695|T191|SYGB|31396002|SNOMEDCT_US|Mucocarcinoid tumour|8243/3
C0205695|T191|SYGB|31396002|SNOMEDCT_US|Mucocarcinoid tumour, malignant|8243/3
C0334302|T191|PT|0000029955|CHV|adenocarcinoid tumor|8244/3
C0334302|T191|LA|LA26102-6|LNC|Mixed adenoneuroendocrine carcinoma|8244/3
C0334302|T191|LLT|10076748|MDR|Mixed adenoneuroendocrine carcinoma|8244/3
C0334302|T191|PT|10076748|MDR|Mixed adenoneuroendocrine carcinoma|8244/3
C0334302|T191|PT|271486|MEDCIN|adenocarcinoid tumor|8244/3
C0334302|T191|PT|271485|MEDCIN|composite carcinoid tumor|8244/3
C0334302|T191|NM|C538230|MSH|Adenocarcinoid tumor|8244/3
C0334302|T191|PN|NOCODE|MTH|Adenocarcinoid tumor|8244/3
C2987129|T191|PN|NOCODE|MTH|Gastrointestinal Mixed Adenoneuroendocrine Carcinoma|8244/3
C0334302|T191|SY|C4139|NCI|Adenocarcinoid Neoplasm|8244/3
C0334302|T191|SY|C4139|NCI|Adenocarcinoid Tumor|8244/3
C0334302|T191|PT|C4139|NCI|Combined Carcinoid and Adenocarcinoma|8244/3
C0334302|T191|SY|C4139|NCI|Combined Carcinoid Neoplasm and Adenocarcinoma|8244/3
C0334302|T191|SY|C4139|NCI|Combined Carcinoid Tumor and Adenocarcinoma|8244/3
C0334302|T191|SY|C4139|NCI|Composite Carcinoid|8244/3
C0334302|T191|SY|C4139|NCI|Composite Carcinoid Neoplasm|8244/3
C0334302|T191|SY|C4139|NCI|Composite Carcinoid Tumor|8244/3
C2987129|T191|PT|C95406|NCI|Digestive System Mixed Adenoneuroendocrine Carcinoma|8244/3
C2987129|T191|SY|C95406|NCI|Gastrointestinal MANEC|8244/3
C2987129|T191|SY|C95406|NCI|Gastrointestinal Mixed Adenoneuroendocrine Carcinoma|8244/3
C2987129|T191|AB|C95406|NCI|MANEC|8244/3
C2987129|T191|SY|C95406|NCI|Mixed Adenoneuroendocrine Carcinoma|8244/3
C0334302|T191|SY|C4139|NCI|Mixed Carcinoid Neoplasm|8244/3
C0334302|T191|SY|C4139|NCI|Mixed Carcinoid Tumor|8244/3
C0334302|T191|PT|C4139|NCI_CPTAC|Combined Carcinoid and Adenocarcinoma|8244/3
C2987129|T191|DN|C95406|NCI_CTRP|Digestive System Mixed Adenoneuroendocrine Cancer|8244/3
C0334302|T191|PT|X77nU|RCD|Adenocarcinoid tumour|8244/3
C0334302|T191|AB|BB5R7|RCD|Combined carcinoid + adenoca|8244/3
C0334302|T191|SY|BB5R7|RCD|Combined carcinoid and adenocarcinoma|8244/3
C0334302|T191|PT|BB5R7|RCD|Composite carcinoid|8244/3
C0334302|T191|PT|X77nU|RCDAE|Adenocarcinoid tumor|8244/3
C0334302|T191|OAP|189614008|SNOMEDCT_US|Adenocarcinoid tumor|8244/3
C0334302|T191|PT|86293007|SNOMEDCT_US|Adenocarcinoid tumor|8244/3
C0334302|T191|OAP|189614008|SNOMEDCT_US|Adenocarcinoid tumour|8244/3
C0334302|T191|OF|189614008|SNOMEDCT_US|Adenocarcinoid tumour|8244/3
C0334302|T191|PTGB|86293007|SNOMEDCT_US|Adenocarcinoid tumour|8244/3
C0334302|T191|SY|51465000|SNOMEDCT_US|Combined carcinoid and adenocarcinoma|8244/3
C0334302|T191|SY|51465000|SNOMEDCT_US|Composite carcinoid|8244/3
C0334302|T191|SY|51465000|SNOMEDCT_US|MANEC|8244/3
C0334302|T191|PT|51465000|SNOMEDCT_US|Mixed adenoneuroendocrine carcinoma|8244/3
C0334302|T191|SY|51465000|SNOMEDCT_US|Mixed carcinoid-adenocarcinoma|8244/3
C1706835|T191|PT|C43565|NCI|Appendix Tubular Carcinoid|8245/1
C1706835|T191|SY|C43565|NCI|Appendix Tubular Carcinoid Tumor|8245/1
C1266031|T191|PT|128889005|SNOMEDCT_US|Tubular carcinoid|8245/1
C0334302|T191|PT|0000029955|CHV|adenocarcinoid tumor|8245/3
C0334302|T191|LA|LA26102-6|LNC|Mixed adenoneuroendocrine carcinoma|8245/3
C0334302|T191|LLT|10076748|MDR|Mixed adenoneuroendocrine carcinoma|8245/3
C0334302|T191|PT|10076748|MDR|Mixed adenoneuroendocrine carcinoma|8245/3
C0334302|T191|PT|271486|MEDCIN|adenocarcinoid tumor|8245/3
C0334302|T191|PT|271485|MEDCIN|composite carcinoid tumor|8245/3
C0334302|T191|NM|C538230|MSH|Adenocarcinoid tumor|8245/3
C0334302|T191|PN|NOCODE|MTH|Adenocarcinoid tumor|8245/3
C0334302|T191|SY|C4139|NCI|Adenocarcinoid Neoplasm|8245/3
C0334302|T191|SY|C4139|NCI|Adenocarcinoid Tumor|8245/3
C0334302|T191|PT|C4139|NCI|Combined Carcinoid and Adenocarcinoma|8245/3
C0334302|T191|SY|C4139|NCI|Combined Carcinoid Neoplasm and Adenocarcinoma|8245/3
C0334302|T191|SY|C4139|NCI|Combined Carcinoid Tumor and Adenocarcinoma|8245/3
C0334302|T191|SY|C4139|NCI|Composite Carcinoid|8245/3
C0334302|T191|SY|C4139|NCI|Composite Carcinoid Neoplasm|8245/3
C0334302|T191|SY|C4139|NCI|Composite Carcinoid Tumor|8245/3
C0334302|T191|SY|C4139|NCI|Mixed Carcinoid Neoplasm|8245/3
C0334302|T191|SY|C4139|NCI|Mixed Carcinoid Tumor|8245/3
C0334302|T191|PT|C4139|NCI_CPTAC|Combined Carcinoid and Adenocarcinoma|8245/3
C0334302|T191|PT|X77nU|RCD|Adenocarcinoid tumour|8245/3
C0334302|T191|AB|BB5R7|RCD|Combined carcinoid + adenoca|8245/3
C0334302|T191|SY|BB5R7|RCD|Combined carcinoid and adenocarcinoma|8245/3
C0334302|T191|PT|BB5R7|RCD|Composite carcinoid|8245/3
C0334302|T191|PT|X77nU|RCDAE|Adenocarcinoid tumor|8245/3
C0334302|T191|OAP|189614008|SNOMEDCT_US|Adenocarcinoid tumor|8245/3
C0334302|T191|PT|86293007|SNOMEDCT_US|Adenocarcinoid tumor|8245/3
C0334302|T191|PTGB|86293007|SNOMEDCT_US|Adenocarcinoid tumour|8245/3
C0334302|T191|OAP|189614008|SNOMEDCT_US|Adenocarcinoid tumour|8245/3
C0334302|T191|OF|189614008|SNOMEDCT_US|Adenocarcinoid tumour|8245/3
C0334302|T191|SY|51465000|SNOMEDCT_US|Combined carcinoid and adenocarcinoma|8245/3
C0334302|T191|SY|51465000|SNOMEDCT_US|Composite carcinoid|8245/3
C0334302|T191|SY|51465000|SNOMEDCT_US|MANEC|8245/3
C0334302|T191|PT|51465000|SNOMEDCT_US|Mixed adenoneuroendocrine carcinoma|8245/3
C0334302|T191|SY|51465000|SNOMEDCT_US|Mixed carcinoid-adenocarcinoma|8245/3
C0206695|T191|SY|0000021027|CHV|carcinoma neuroendocrine|8246/3
C0206754|T191|SY|0000056678|CHV|neoplasms neuroendocrine|8246/3
C0206695|T191|PT|0000021027|CHV|neuroendocrine carcinoma|8246/3
C0206695|T191|SY|0000021027|CHV|neuroendocrine carcinomas|8246/3
C0206754|T191|PT|0000056678|CHV|neuroendocrine neoplasm|8246/3
C0206754|T191|PT|0000021067|CHV|neuroendocrine tumor|8246/3
C0206754|T191|SY|0000021067|CHV|neuroendocrine tumors|8246/3
C0206754|T191|SY|0000021067|CHV|neuroendocrine tumour|8246/3
C0206754|T191|SY|0000021067|CHV|neuroendocrine tumours|8246/3
C0206754|T191|SY|HP:0100634|HPO|Neuroendocrine neoplasia|8246/3
C0206754|T191|PT|HP:0100634|HPO|Neuroendocrine neoplasm|8246/3
C0206754|T191|ET|D3A.8|ICD10CM|Neuroendocrine tumor NOS|8246/3
C0206754|T191|HT|209-209.99|ICD9CM|NEUROENDOCRINE TUMORS|8246/3
C0206754|T191|HT|209|ICD9CM|Neuroendocrine tumors|8246/3
C0206754|T191|PT|sh94005134|LCH_NW|Neuroendocrine tumors|8246/3
C0206695|T191|LA|LA26099-4|LNC|Neuroendocrine carcinoma|8246/3
C0206695|T191|LA|LA26506-8|LNC|Neuroendocrine carcinoma, NOS|8246/3
C0206695|T191|LLT|10057270|MDR|Neuroendocrine carcinoma|8246/3
C0206695|T191|PT|10057270|MDR|Neuroendocrine carcinoma|8246/3
C0206754|T191|LLT|10062476|MDR|Neuroendocrine tumor|8246/3
C0206754|T191|MTH_PT|10052399|MDR|Neuroendocrine tumor|8246/3
C0206754|T191|LLT|10052399|MDR|Neuroendocrine tumour|8246/3
C0206754|T191|PT|10052399|MDR|Neuroendocrine tumour|8246/3
C0206695|T191|PT|271448|MEDCIN|neuroendocrine carcinoma|8246/3
C0206754|T191|PT|352608|MEDCIN|Neuroendocrine tumor|8246/3
C0206695|T191|MH|D018278|MSH|Carcinoma, Neuroendocrine|8246/3
C0206695|T191|PM|D018278|MSH|Carcinomas, Neuroendocrine|8246/3
C0206695|T191|PM|D018278|MSH|Neuroendocrine Carcinoma|8246/3
C0206695|T191|PM|D018278|MSH|Neuroendocrine Carcinomas|8246/3
C0206754|T191|PM|D018358|MSH|Neuroendocrine Tumor|8246/3
C0206754|T191|MH|D018358|MSH|Neuroendocrine Tumors|8246/3
C0206754|T191|PM|D018358|MSH|Tumor, Neuroendocrine|8246/3
C0206754|T191|PM|D018358|MSH|Tumors, Neuroendocrine|8246/3
C0206695|T191|PN|NOCODE|MTH|Carcinoma, Neuroendocrine|8246/3
C0206754|T191|ET|209.60|MTHICD9|Neuroendocrine tumor NOS|8246/3
C1266149|T191|OP|C35726|NCI|Grade III Neuroendocrine Carcinoma|8246/3
C1266149|T191|PT|C35726|NCI|Grade III Neuroendocrine Carcinoma|8246/3
C0206695|T191|AB|C3773|NCI|NEC|8246/3
C0206695|T191|PT|C3773|NCI|Neuroendocrine Carcinoma|8246/3
C0206754|T191|PT|C3809|NCI|Neuroendocrine Neoplasm|8246/3
C0206695|T191|PT|C3773|NCI_CPTAC|Neuroendocrine Carcinoma|8246/3
C0206754|T191|PT|C3809|NCI_CPTAC|Neuroendocrine Neoplasm|8246/3
C0206695|T191|PT|10057270|NCI_CTEP-SDC|Neuroendocrine cancer, NOS|8246/3
C0206695|T191|DN|C3773|NCI_CTRP|Neuroendocrine Cancer|8246/3
C0206695|T191|PT|C3773|NCI_CTRP|Neuroendocrine Cancer|8246/3
C0206695|T191|SY|C3773|NCI_CTRP|Neuroendocrine Carcinoma|8246/3
C0206754|T191|SY|C3809|NCI_CTRP|Neuroendocrine Neoplasm|8246/3
C0206754|T191|DN|C3809|NCI_CTRP|Neuroendocrine Tumor|8246/3
C0206754|T191|PT|C3809|NCI_CTRP|Neuroendocrine Tumor|8246/3
C0206754|T191|PT|CDR0000044904|NCI_NCI-GLOSS|neuroendocrine tumor|8246/3
C0206754|T191|PT|C3809|NCI_NICHD|Neuroendocrine Tumor|8246/3
C0206695|T191|SY|CDR0000038259|PDQ|carcinoma, neuroendocrine|8246/3
C0206695|T191|ET|CDR0000038259|PDQ|Neuroendocrine carcinoma|8246/3
C0206695|T191|PSC|CDR0000038259|PDQ|neuroendocrine carcinoma|8246/3
C0206754|T191|PT|CDR0000550683|PDQ|neuroendocrine neoplasm|8246/3
C0206754|T191|SY|CDR0000550683|PDQ|neuroendocrine tumor|8246/3
C0206695|T191|PT|X77nQ|RCD|Neuroendocrine carcinoma|8246/3
C0206754|T191|PT|X78dr|RCD|Neuroendocrine tumour|8246/3
C0457185|T191|AB|Xa0aO|RCD|Olfact neuroendocrine carcinom|8246/3
C0457185|T191|PT|Xa0aO|RCD|Olfactory neuroendocrine carcinoma|8246/3
C0206754|T191|PT|X78dr|RCDAE|Neuroendocrine tumor|8246/3
C0206695|T191|OP|BB5R9|RCDSY|Neuroendocrine carcinoma|8246/3
C1266150|T191|PT|127575007|SNOMEDCT_US|Malignant neuroendocrine neoplasm, epithelial|8246/3
C5191660|T191|SY|785766008|SNOMEDCT_US|MiNEN - mixed neuroendocrine-non neuroendocrine neoplasm|8246/3
C5191660|T191|PT|785766008|SNOMEDCT_US|Mixed neuroendocrine-non neuroendocrine neoplasm|8246/3
C0206695|T191|PT|253000007|SNOMEDCT_US|Neuroendocrine carcinoma|8246/3
C0206695|T191|SY|55937004|SNOMEDCT_US|Neuroendocrine carcinoma|8246/3
C1266149|T191|SY|127574006|SNOMEDCT_US|Neuroendocrine carcinoma, grade 3|8246/3
C0206754|T191|PT|128928004|SNOMEDCT_US|Neuroendocrine neoplasm|8246/3
C0206754|T191|PT|55937004|SNOMEDCT_US|Neuroendocrine tumor|8246/3
C0206754|T191|PT|255046005|SNOMEDCT_US|Neuroendocrine tumor|8246/3
C1266149|T191|PT|127574006|SNOMEDCT_US|Neuroendocrine tumor grade 3|8246/3
C0206754|T191|PTGB|55937004|SNOMEDCT_US|Neuroendocrine tumour|8246/3
C0206754|T191|PTGB|255046005|SNOMEDCT_US|Neuroendocrine tumour|8246/3
C1266149|T191|PTGB|127574006|SNOMEDCT_US|Neuroendocrine tumour grade 3|8246/3
C0457185|T191|PT|277993001|SNOMEDCT_US|Olfactory neuroendocrine carcinoma|8246/3
C0007129|T191|SY|0000002431|CHV|carcinoma cell merkels|8247/3
C0007129|T191|SY|0000002431|CHV|carcinoma neuroendocrine skin|8247/3
C0007129|T191|SY|0000002431|CHV|cell merkel tumors|8247/3
C0007129|T191|SY|0000002431|CHV|mcc|8247/3
C0007129|T191|SY|0000002431|CHV|merkel cell cancer|8247/3
C0007129|T191|PT|0000002431|CHV|merkel cell carcinoma|8247/3
C0007129|T191|SY|0000002431|CHV|merkel cell tumor|8247/3
C0007129|T191|SY|0000002431|CHV|merkel cell tumour|8247/3
C0007129|T191|SY|HP:0030447|HPO|Anaplastic carcinoma of the skin|8247/3
C0007129|T191|SY|HP:0030447|HPO|Cutaneous APUDoma|8247/3
C0007129|T191|SY|HP:0030447|HPO|Merkel cell cancer of the skin|8247/3
C0007129|T191|PT|HP:0030447|HPO|Merkel cell skin cancer|8247/3
C0007129|T191|SY|HP:0030447|HPO|Neuroendocrine carcinoma of the skin|8247/3
C0007129|T191|SY|HP:0030447|HPO|Neuroendocrine tumor of the skin|8247/3
C0007129|T191|SY|HP:0030447|HPO|Primary small cell carcinoma of the skin|8247/3
C0007129|T191|SY|HP:0030447|HPO|Primary undifferentiated carcinoma of the skin|8247/3
C0007129|T191|AB|C4A|ICD10CM|Merkel cell carcinoma|8247/3
C0007129|T191|HT|C4A|ICD10CM|Merkel cell carcinoma|8247/3
C0007129|T191|ET|C4A.9|ICD10CM|Merkel cell carcinoma NOS|8247/3
C0007129|T191|PT|sh00000069|LCH_NW|Merkel cell carcinoma|8247/3
C0007129|T191|LLT|10064025|MDR|Merkel cell carcinoma|8247/3
C0007129|T191|LLT|10029266|MDR|Neuroendocrine carcinoma of the skin|8247/3
C0007129|T191|PT|10029266|MDR|Neuroendocrine carcinoma of the skin|8247/3
C0007129|T191|PT|355432|MEDCIN|Apudoma of skin|8247/3
C0007129|T191|SY|355432|MEDCIN|neuroendocrine tumor apudoma of skin|8247/3
C0007129|T191|ET|405|MEDLINEPLUS|Merkel Cell Cancer|8247/3
C0007129|T191|PM|D015266|MSH|Cancer, Merkel Cell|8247/3
C0007129|T191|MH|D015266|MSH|Carcinoma, Merkel Cell|8247/3
C0007129|T191|PM|D015266|MSH|Cell Cancer, Merkel|8247/3
C0007129|T191|ET|D015266|MSH|Merkel Cell Cancer|8247/3
C0007129|T191|ET|D015266|MSH|Merkel Cell Carcinoma|8247/3
C0007129|T191|ET|D015266|MSH|Merkel Cell Tumor|8247/3
C0007129|T191|ET|D015266|MSH|Merkle Tumors|8247/3
C0007129|T191|PM|D015266|MSH|Tumor, Merkel Cell|8247/3
C0007129|T191|PM|D015266|MSH|Tumors, Merkle|8247/3
C0007129|T191|PN|NOCODE|MTH|Merkel cell carcinoma|8247/3
C0007129|T191|ET|209.36|MTHICD9|Merkel cell carcinoma NOS|8247/3
C0007129|T191|SY|C9231|NCI|Cutaneous Apudoma|8247/3
C0007129|T191|SY|C9231|NCI|Cutaneous Neuroendocrine Carcinoma|8247/3
C0007129|T191|PT|C9231|NCI|Merkel Cell Carcinoma|8247/3
C0007129|T191|SY|C9231|NCI|Neuroendocrine Carcinoma of Skin|8247/3
C0007129|T191|SY|C9231|NCI|Neuroendocrine Carcinoma of the Skin|8247/3
C0007129|T191|SY|C9231|NCI|Neuroendocrine Skin Carcinoma|8247/3
C0007129|T191|SY|C9231|NCI|Trabecular Skin Carcinoma|8247/3
C0007129|T191|PT|C9231|NCI_CPTAC|Merkel Cell Carcinoma|8247/3
C0007129|T191|PT|10029266|NCI_CTEP-SDC|Merkel cell tumor|8247/3
C0007129|T191|DN|C9231|NCI_CTRP|Merkel Cell Cancer|8247/3
C0007129|T191|PT|CDR0000046106|NCI_NCI-GLOSS|Merkel cell cancer|8247/3
C0007129|T191|PT|CDR0000658511|NCI_NCI-GLOSS|Merkel cell carcinoma|8247/3
C0007129|T191|PT|CDR0000579914|NCI_NCI-GLOSS|neuroendocrine carcinoma of the skin|8247/3
C0007129|T191|PT|CDR0000386222|NCI_NCI-GLOSS|trabecular cancer|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|adult neuroblastoma of the skin|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|carcinoma, Merkel cell|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|cutaneous APUDoma|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|cutaneous neuroendocrine tumor|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|endocrine carcinoma of the skin|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|MCC|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|Merkel cell cancer|8247/3
C0007129|T191|PSC|CDR0000038240|PDQ|Merkel cell carcinoma|8247/3
C0007129|T191|ET|CDR0000038240|PDQ|Merkel cell carcinoma|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|neuroendocrine carcinoma of the skin|8247/3
C0007129|T191|OP|CDR0000041900|PDQ|neuroendocrine carcinoma of the skin|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|primary small cell carcinoma of the skin|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|small cell neuroepithelial tumor of the skin|8247/3
C0007129|T191|SY|CDR0000038240|PDQ|trabecular carcinoma of the skin|8247/3
C0007129|T191|OP|X78T9|RCD|Apudoma of skin|8247/3
C0007129|T191|PT|X77nR|RCD|Merkel cell carcinoma|8247/3
C0007129|T191|SY|X77nR|RCD|Merkel cell tumour|8247/3
C0007129|T191|AB|X77nR|RCD|Trabecular cell carcinoma|8247/3
C0007129|T191|SY|X77nR|RCD|Trabecular cell carcinoma of skin|8247/3
C0007129|T191|SY|X77nR|RCDAE|Merkel cell tumor|8247/3
C0007129|T191|OP|BB5RA|RCDSY|Merkel cell carcinoma|8247/3
C0007129|T191|PT|254729005|SNOMEDCT_US|Apudoma of skin|8247/3
C0007129|T191|PT|253001006|SNOMEDCT_US|Merkel cell carcinoma|8247/3
C0007129|T191|PT|5052009|SNOMEDCT_US|Merkel cell carcinoma|8247/3
C0007129|T191|SY|5052009|SNOMEDCT_US|Merkel cell tumor|8247/3
C0007129|T191|SY|253001006|SNOMEDCT_US|Merkel cell tumor|8247/3
C0007129|T191|SYGB|253001006|SNOMEDCT_US|Merkel cell tumour|8247/3
C0007129|T191|SYGB|5052009|SNOMEDCT_US|Merkel cell tumour|8247/3
C0007129|T191|SY|5052009|SNOMEDCT_US|Primary cutaneous neuroendocrine carcinoma|8247/3
C0007129|T191|SY|253001006|SNOMEDCT_US|Trabecular cell carcinoma of skin|8247/3
C0003650|T191|PT|0000001404|CHV|apudoma|8248/1
C0003650|T191|SY|0000001404|CHV|apudomas|8248/1
C0003650|T191|SY|HP:0040192|HPO|amine precursor uptake and decarboxylation tumours|8248/1
C0003650|T191|PT|HP:0040192|HPO|APUdoma|8248/1
C0003650|T191|LLT|10003069|MDR|APUDoma|8248/1
C0003650|T191|PT|10003069|MDR|APUDoma|8248/1
C0003650|T191|LLT|10003070|MDR|APUDoma NOS|8248/1
C0003650|T191|PT|355431|MEDCIN|Apudoma|8248/1
C0003650|T191|SY|355431|MEDCIN|neuroendocrine tumor apudoma|8248/1
C0003650|T191|MH|D001079|MSH|Apudoma|8248/1
C0003650|T191|PM|D001079|MSH|Apudomas|8248/1
C0003650|T191|OP|C2879|NCI|Apudoma|8248/1
C0003650|T191|SY|C2879|NCI|Neoplasm of Diffuse Neuroendocrine System|8248/1
C0003650|T191|PT|C2879|NCI|Neoplasm of the Diffuse Neuroendocrine System|8248/1
C0003650|T191|PT|X77nZ|RCD|Apudoma|8248/1
C0003650|T191|OP|BB5y3|RCDSY|Apudoma|8248/1
C0003650|T191|PT|253008000|SNOMEDCT_US|Apudoma|8248/1
C0003650|T191|PT|74926005|SNOMEDCT_US|Apudoma|8248/1
C1266032|T191|PT|271487|MEDCIN|atypical carcinoid tumor|8249/3
C1708766|T191|PT|219650|MEDCIN|atypical carcinoid tumor of lung|8249/3
C1708766|T191|PT|219644|MEDCIN|malignant carcinoid tumor of lung|8249/3
C1266032|T191|PN|NOCODE|MTH|Atypical carcinoid tumor|8249/3
C1266032|T191|SY|TCGA|NCI|Atypical Carcinoid Tumor|8249/3
C1266032|T191|PT|C72074|NCI|Atypical Carcinoid Tumor|8249/3
C3272617|T191|PT|C96166|NCI|Digestive System Neuroendocrine Tumor G2|8249/3
C3272617|T191|SY|C96166|NCI|Gastrointestinal NET G2|8249/3
C3272617|T191|SY|C96166|NCI|Gastrointestinal Neuroendocrine Tumor G2|8249/3
C1333862|T191|OP|C35725|NCI|Grade II Neuroendocrine Carcinoma|8249/3
C1333862|T191|PT|C35725|NCI|Grade II Neuroendocrine Carcinoma|8249/3
C1708766|T191|PT|C45551|NCI|Lung Atypical Carcinoid Tumor|8249/3
C1708766|T191|SY|C45551|NCI|Lung Malignant Carcinoid Tumor|8249/3
C1266032|T191|SY|C72074|NCI|Malignant Carcinoid Tumor|8249/3
C1708766|T191|PT|C45551|NCI_CPTAC|Lung Atypical Carcinoid Tumor|8249/3
C1266032|T191|PT|128658008|SNOMEDCT_US|Atypical carcinoid tumor|8249/3
C1266032|T191|PTGB|128658008|SNOMEDCT_US|Atypical carcinoid tumour|8249/3
C1266148|T191|SY|127573000|SNOMEDCT_US|Grade 2 neuroendocrine carcinoma|8249/3
C1708766|T191|PT|123661000119106|SNOMEDCT_US|Malignant carcinoid tumor of lung|8249/3
C1708766|T191|IS|123661000119106|SNOMEDCT_US|Malignant carcinoid tumour of lung|8249/3
C1266148|T191|SY|127573000|SNOMEDCT_US|Moderately differentiated neuroendocrine carcinoma|8249/3
C1266148|T191|SY|127573000|SNOMEDCT_US|Neuroendocrine carcinoma, grade 2|8249/3
C1266148|T191|PT|127573000|SNOMEDCT_US|Neuroendocrine tumor grade 2|8249/3
C1266148|T191|PTGB|127573000|SNOMEDCT_US|Neuroendocrine tumour grade 2|8249/3
C0206676|T191|PT|MTHU003465|ICPC2ICD10ENG|adenomatosis; pulmonary|8250/1
C0206676|T191|PT|MTHU062956|ICPC2ICD10ENG|pulmonary; adenomatosis|8250/1
C0206676|T191|PT|sh85108994|LCH_NW|Pulmonary adenomatosis|8250/1
C0206676|T191|LLT|10037311|MDR|Pulmonary adenomatosis|8250/1
C0206676|T191|PM|D018255|MSH|Adenomatoses, Pulmonary|8250/1
C0206676|T191|DEV|D018255|MSH|ADENOMATOSIS PULM|8250/1
C0206676|T191|MH|D018255|MSH|Adenomatosis, Pulmonary|8250/1
C0206676|T191|DEV|D018255|MSH|PULM ADENOMATOSIS|8250/1
C0206676|T191|PM|D018255|MSH|Pulmonary Adenomatoses|8250/1
C0206676|T191|ET|D018255|MSH|Pulmonary Adenomatosis|8250/1
C0206676|T191|OP|C3763|NCI|Pulmonary Adenomatosis|8250/1
C0206676|T191|PT|C3763|NCI|Pulmonary Adenomatosis|8250/1
C0206676|T191|PT|BB5S0|RCD|Pulmonary adenomatosis|8250/1
C0206676|T191|PT|32434004|SNOMEDCT_US|Pulmonary adenomatosis|8250/1
C0007120|T191|NP|0000023036|AOD|alveolar cell carcinoma|8250/3
C0007120|T191|SY|0000002427|CHV|alveolar carcinoma|8250/3
C0007120|T191|SY|0000002427|CHV|alveolar cell carcinoma|8250/3
C0007120|T191|PT|0000050168|CHV|bronchioalveolar carcinoma|8250/3
C0007120|T191|SY|0000002427|CHV|bronchiolar carcinoma|8250/3
C0007120|T191|SY|0000002427|CHV|bronchiolo-alveolar carcinoma|8250/3
C0007120|T191|PT|0000002427|CHV|bronchioloalveolar carcinoma|8250/3
C0007120|T191|SY|NOCODE|DXP|CARCINOMA, ALVEOLAR|8250/3
C0007120|T191|SY|NOCODE|DXP|CARCINOMA, ALVEOLAR CELL|8250/3
C0007120|T191|SY|NOCODE|DXP|CARCINOMA, BRONCHIOLOALVEOLAR|8250/3
C0007120|T191|PT|HP:0006519|HPO|Alveolar cell carcinoma|8250/3
C0007120|T191|LLT|10049876|MDR|Alveolar cell carcinoma|8250/3
C0007120|T191|LLT|10006447|MDR|Bronchioalveolar carcinoma|8250/3
C0007120|T191|LLT|10058354|MDR|Bronchioloalveolar carcinoma|8250/3
C0007120|T191|PT|10058354|MDR|Bronchioloalveolar carcinoma|8250/3
C0007120|T191|PT|271477|MEDCIN|alveolar adenocarcinoma|8250/3
C0007120|T191|PT|31594|MEDCIN|bronchiolo-alveolar adenocarcinoma of lung|8250/3
C0007120|T191|ET|D002282|MSH|Adenocarcinoma, Alveolar|8250/3
C0007120|T191|PM|D002282|MSH|Adenocarcinoma, Bronchiolo Alveolar|8250/3
C0007120|T191|MH|D002282|MSH|Adenocarcinoma, Bronchiolo-Alveolar|8250/3
C0007120|T191|PM|D002282|MSH|Adenocarcinomas, Alveolar|8250/3
C0007120|T191|PM|D002282|MSH|Adenocarcinomas, Bronchiolo-Alveolar|8250/3
C0007120|T191|PM|D002282|MSH|Alveolar Adenocarcinoma|8250/3
C0007120|T191|PM|D002282|MSH|Alveolar Adenocarcinomas|8250/3
C0007120|T191|PM|D002282|MSH|Alveolar Carcinoma|8250/3
C0007120|T191|PM|D002282|MSH|Alveolar Carcinomas|8250/3
C0007120|T191|ET|D002282|MSH|Alveolar Cell Carcinoma|8250/3
C0007120|T191|PM|D002282|MSH|Alveolar Cell Carcinomas|8250/3
C0007120|T191|PM|D002282|MSH|Bronchiolar Carcinoma|8250/3
C0007120|T191|PM|D002282|MSH|Bronchiolar Carcinomas|8250/3
C0007120|T191|PM|D002282|MSH|Bronchiolo-Alveolar Adenocarcinoma|8250/3
C0007120|T191|PM|D002282|MSH|Bronchiolo-Alveolar Adenocarcinomas|8250/3
C0007120|T191|PM|D002282|MSH|Bronchiolo-Alveolar Carcinoma|8250/3
C0007120|T191|PM|D002282|MSH|Bronchiolo-Alveolar Carcinomas|8250/3
C0007120|T191|PM|D002282|MSH|Bronchioloalveolar Carcinoma|8250/3
C0007120|T191|PM|D002282|MSH|Bronchioloalveolar Carcinomas|8250/3
C0007120|T191|ET|D002282|MSH|Carcinoma, Alveolar|8250/3
C0007120|T191|PM|D002282|MSH|Carcinoma, Alveolar Cell|8250/3
C0007120|T191|ET|D002282|MSH|Carcinoma, Bronchiolar|8250/3
C0007120|T191|PM|D002282|MSH|Carcinoma, Bronchiolo Alveolar|8250/3
C0007120|T191|ET|D002282|MSH|Carcinoma, Bronchiolo-Alveolar|8250/3
C0007120|T191|ET|D002282|MSH|Carcinoma, Bronchioloalveolar|8250/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Alveolar|8250/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Alveolar Cell|8250/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Bronchiolar|8250/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Bronchiolo-Alveolar|8250/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Bronchioloalveolar|8250/3
C0007120|T191|PN|NOCODE|MTH|Bronchioloalveolar Adenocarcinoma|8250/3
C0007120|T191|AB|C2923|NCI|BAC|8250/3
C0007120|T191|OP|C2923|NCI|Bronchioalveolar Adenocarcinoma of Lung|8250/3
C0007120|T191|OP|C2923|NCI|Bronchioalveolar Adenocarcinoma of the Lung|8250/3
C0007120|T191|OP|C2923|NCI|Bronchioalveolar Lung Carcinoma|8250/3
C0007120|T191|OP|C2923|NCI|Bronchiolo-Alveolar Carcinoma of Lung|8250/3
C0007120|T191|OP|C2923|NCI|Bronchiolo-Alveolar Carcinoma of the Lung|8250/3
C0007120|T191|OP|C2923|NCI|Bronchiolo-Alveolar Lung Carcinoma|8250/3
C0007120|T191|OP|C2923|NCI|Bronchioloalveolar Adenocarcinoma of Lung|8250/3
C0007120|T191|OP|C2923|NCI|Bronchioloalveolar Adenocarcinoma of the Lung|8250/3
C0007120|T191|OP|C2923|NCI|Bronchioloalveolar Carcinoma|8250/3
C0007120|T191|OP|C2923|NCI|Bronchioloalveolar Lung Adenocarcinoma|8250/3
C0007120|T191|PT|C2923|NCI|Minimally Invasive Lung Adenocarcinoma|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|BAC|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioalveolar Adenocarcinoma of Lung|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioalveolar Adenocarcinoma of the Lung|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioalveolar Lung Carcinoma|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchiolo-Alveolar Carcinoma of Lung|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchiolo-Alveolar Carcinoma of the Lung|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchiolo-Alveolar Lung Carcinoma|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioloalveolar Adenocarcinoma of Lung|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioloalveolar Adenocarcinoma of the Lung|8250/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioloalveolar Lung Adenocarcinoma|8250/3
C0007120|T191|PT|C2923|NCI_CDISC|CARCINOMA, BRONCHIOLOALVEOLAR, MALIGNANT|8250/3
C0007120|T191|PT|10058354|NCI_CTEP-SDC|Bronchioloalveolar carcinoma|8250/3
C0007120|T191|DN|C2923|NCI_CTRP|Bronchioloalveolar Carcinoma|8250/3
C0007120|T191|AB|CDR0000043303|PDQ|BAC|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioalveolar Adenocarcinoma of Lung|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioalveolar Adenocarcinoma of the Lung|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioalveolar Lung Carcinoma|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchiolo-Alveolar Carcinoma of Lung|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchiolo-Alveolar Carcinoma of the Lung|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchiolo-Alveolar Lung Carcinoma|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioloalveolar Adenocarcinoma of Lung|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioloalveolar Adenocarcinoma of the Lung|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|bronchioloalveolar carcinoma|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioloalveolar Lung Adenocarcinoma|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|bronchoalveolar carcinoma|8250/3
C0007120|T191|PT|CDR0000043303|PDQ|bronchoalveolar cell lung cancer|8250/3
C0007120|T191|SY|CDR0000043303|PDQ|lung cancer, bronchoalveolar cell|8250/3
C0007120|T191|PT|R0121358|QMR|BRONCHIOLAR-ALVEOLAR CELL CARCINOMA|8250/3
C0007120|T191|PT|BB5S4|RCD|Alveolar adenocarcinoma|8250/3
C0007120|T191|SY|BB5S4|RCD|Alveolar carcinoma|8250/3
C0007120|T191|SY|XaBAp|RCD|Alveolar cell carcinoma|8250/3
C0007120|T191|AB|XaBAp|RCD|Bronchio-alveol adenocarc lung|8250/3
C0007120|T191|SY|XaBAp|RCD|Bronchiolar adenocarcinoma|8250/3
C0007120|T191|SY|XaBAp|RCD|Bronchiolar carcinoma|8250/3
C0007120|T191|AB|XaBAp|RCD|Bronchiolo-alveolar adenoca|8250/3
C0007120|T191|SY|XaBAp|RCD|Bronchiolo-alveolar adenocarcinoma|8250/3
C0007120|T191|PT|XaBAp|RCD|Bronchiolo-alveolar adenocarcinoma of lung|8250/3
C0007120|T191|SY|XaBAp|RCD|Bronchiolo-alveolar carcinoma|8250/3
C0007120|T191|SY|XaBAp|RCD|Bronchioloalveolar carcinoma|8250/3
C0007120|T191|AB|BB5S2|RCDSY|Bronchiolo-alveolar adenoca|8250/3
C0007120|T191|PT|BB5S2|RCDSY|Bronchiolo-alveolar adenocarcinoma|8250/3
C0007120|T191|PT|36310008|SNOMEDCT_US|Alveolar adenocarcinoma|8250/3
C0007120|T191|SY|36310008|SNOMEDCT_US|Alveolar carcinoma|8250/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Alveolar cell carcinoma|8250/3
C0007120|T191|SY|112677002|SNOMEDCT_US|Alveolar cell carcinoma|8250/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Bronchiolar adenocarcinoma|8250/3
C0007120|T191|SY|112677002|SNOMEDCT_US|Bronchiolar adenocarcinoma|8250/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Bronchiolar carcinoma|8250/3
C0007120|T191|SY|112677002|SNOMEDCT_US|Bronchiolar carcinoma|8250/3
C0007120|T191|PT|112677002|SNOMEDCT_US|Bronchiolo-alveolar adenocarcinoma|8250/3
C0007120|T191|SY|112677002|SNOMEDCT_US|Bronchiolo-alveolar carcinoma|8250/3
C0007120|T191|OAS|307595008|SNOMEDCT_US|Bronchioloalveolar adenocarcinoma|8250/3
C0007120|T191|OAP|307595008|SNOMEDCT_US|Bronchioloalveolar adenocarcinoma of lung|8250/3
C0007120|T191|OF|307595008|SNOMEDCT_US|Bronchioloalveolar adenocarcinoma of lung|8250/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Bronchioloalveolar carcinoma|8250/3
C0007120|T191|OAP|373627005|SNOMEDCT_US|Bronchioloalveolar carcinoma - disorder|8250/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Bronchoalveolar cancer|8250/3
C0334303|T191|PT|MTHU003472|ICPC2ICD10ENG|adenoma; alveolar|8251/0
C0334303|T191|PT|MTHU005099|ICPC2ICD10ENG|alveolar; adenoma|8251/0
C0334303|T191|SY|C4140|NCI|Adenoma of Alveoli|8251/0
C0334303|T191|SY|C4140|NCI|Adenoma of the Alveoli|8251/0
C0334303|T191|PT|C4140|NCI|Alveolar Adenoma|8251/0
C0334303|T191|SY|C4140|NCI_CDISC|Adenoma of Alveoli|8251/0
C0334303|T191|SY|C4140|NCI_CDISC|Adenoma of the Alveoli|8251/0
C0334303|T191|PT|C4140|NCI_CDISC|ADENOMA, BRONCHIOLOALVEOLAR, BENIGN|8251/0
C0334303|T191|PT|BB5S3|RCD|Alveolar adenoma|8251/0
C0334303|T191|PT|8097004|SNOMEDCT_US|Alveolar adenoma|8251/0
C4518389|T191|PT|734094002|SNOMEDCT_US|Atypical alveolar adenomatous hyperplasia|8251/0
C0007120|T191|NP|0000023036|AOD|alveolar cell carcinoma|8251/3
C0007120|T191|SY|0000002427|CHV|alveolar carcinoma|8251/3
C0007120|T191|SY|0000002427|CHV|alveolar cell carcinoma|8251/3
C0007120|T191|PT|0000050168|CHV|bronchioalveolar carcinoma|8251/3
C0007120|T191|SY|0000002427|CHV|bronchiolar carcinoma|8251/3
C0007120|T191|SY|0000002427|CHV|bronchiolo-alveolar carcinoma|8251/3
C0007120|T191|PT|0000002427|CHV|bronchioloalveolar carcinoma|8251/3
C0007120|T191|SY|NOCODE|DXP|CARCINOMA, ALVEOLAR|8251/3
C0007120|T191|SY|NOCODE|DXP|CARCINOMA, ALVEOLAR CELL|8251/3
C0007120|T191|SY|NOCODE|DXP|CARCINOMA, BRONCHIOLOALVEOLAR|8251/3
C0007120|T191|PT|HP:0006519|HPO|Alveolar cell carcinoma|8251/3
C0007120|T191|LLT|10049876|MDR|Alveolar cell carcinoma|8251/3
C0007120|T191|LLT|10006447|MDR|Bronchioalveolar carcinoma|8251/3
C0007120|T191|PT|10058354|MDR|Bronchioloalveolar carcinoma|8251/3
C0007120|T191|LLT|10058354|MDR|Bronchioloalveolar carcinoma|8251/3
C0007120|T191|PT|271477|MEDCIN|alveolar adenocarcinoma|8251/3
C0007120|T191|PT|31594|MEDCIN|bronchiolo-alveolar adenocarcinoma of lung|8251/3
C0007120|T191|ET|D002282|MSH|Adenocarcinoma, Alveolar|8251/3
C0007120|T191|PM|D002282|MSH|Adenocarcinoma, Bronchiolo Alveolar|8251/3
C0007120|T191|MH|D002282|MSH|Adenocarcinoma, Bronchiolo-Alveolar|8251/3
C0007120|T191|PM|D002282|MSH|Adenocarcinomas, Alveolar|8251/3
C0007120|T191|PM|D002282|MSH|Adenocarcinomas, Bronchiolo-Alveolar|8251/3
C0007120|T191|PM|D002282|MSH|Alveolar Adenocarcinoma|8251/3
C0007120|T191|PM|D002282|MSH|Alveolar Adenocarcinomas|8251/3
C0007120|T191|PM|D002282|MSH|Alveolar Carcinoma|8251/3
C0007120|T191|PM|D002282|MSH|Alveolar Carcinomas|8251/3
C0007120|T191|ET|D002282|MSH|Alveolar Cell Carcinoma|8251/3
C0007120|T191|PM|D002282|MSH|Alveolar Cell Carcinomas|8251/3
C0007120|T191|PM|D002282|MSH|Bronchiolar Carcinoma|8251/3
C0007120|T191|PM|D002282|MSH|Bronchiolar Carcinomas|8251/3
C0007120|T191|PM|D002282|MSH|Bronchiolo-Alveolar Adenocarcinoma|8251/3
C0007120|T191|PM|D002282|MSH|Bronchiolo-Alveolar Adenocarcinomas|8251/3
C0007120|T191|PM|D002282|MSH|Bronchiolo-Alveolar Carcinoma|8251/3
C0007120|T191|PM|D002282|MSH|Bronchiolo-Alveolar Carcinomas|8251/3
C0007120|T191|PM|D002282|MSH|Bronchioloalveolar Carcinoma|8251/3
C0007120|T191|PM|D002282|MSH|Bronchioloalveolar Carcinomas|8251/3
C0007120|T191|ET|D002282|MSH|Carcinoma, Alveolar|8251/3
C0007120|T191|PM|D002282|MSH|Carcinoma, Alveolar Cell|8251/3
C0007120|T191|ET|D002282|MSH|Carcinoma, Bronchiolar|8251/3
C0007120|T191|PM|D002282|MSH|Carcinoma, Bronchiolo Alveolar|8251/3
C0007120|T191|ET|D002282|MSH|Carcinoma, Bronchiolo-Alveolar|8251/3
C0007120|T191|ET|D002282|MSH|Carcinoma, Bronchioloalveolar|8251/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Alveolar|8251/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Alveolar Cell|8251/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Bronchiolar|8251/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Bronchiolo-Alveolar|8251/3
C0007120|T191|PM|D002282|MSH|Carcinomas, Bronchioloalveolar|8251/3
C0007120|T191|PN|NOCODE|MTH|Bronchioloalveolar Adenocarcinoma|8251/3
C0007120|T191|AB|C2923|NCI|BAC|8251/3
C0007120|T191|OP|C2923|NCI|Bronchioalveolar Adenocarcinoma of Lung|8251/3
C0007120|T191|OP|C2923|NCI|Bronchioalveolar Adenocarcinoma of the Lung|8251/3
C0007120|T191|OP|C2923|NCI|Bronchioalveolar Lung Carcinoma|8251/3
C0007120|T191|OP|C2923|NCI|Bronchiolo-Alveolar Carcinoma of Lung|8251/3
C0007120|T191|OP|C2923|NCI|Bronchiolo-Alveolar Carcinoma of the Lung|8251/3
C0007120|T191|OP|C2923|NCI|Bronchiolo-Alveolar Lung Carcinoma|8251/3
C0007120|T191|OP|C2923|NCI|Bronchioloalveolar Adenocarcinoma of Lung|8251/3
C0007120|T191|OP|C2923|NCI|Bronchioloalveolar Adenocarcinoma of the Lung|8251/3
C0007120|T191|OP|C2923|NCI|Bronchioloalveolar Carcinoma|8251/3
C0007120|T191|OP|C2923|NCI|Bronchioloalveolar Lung Adenocarcinoma|8251/3
C0007120|T191|PT|C2923|NCI|Minimally Invasive Lung Adenocarcinoma|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|BAC|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioalveolar Adenocarcinoma of Lung|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioalveolar Adenocarcinoma of the Lung|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioalveolar Lung Carcinoma|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchiolo-Alveolar Carcinoma of Lung|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchiolo-Alveolar Carcinoma of the Lung|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchiolo-Alveolar Lung Carcinoma|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioloalveolar Adenocarcinoma of Lung|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioloalveolar Adenocarcinoma of the Lung|8251/3
C0007120|T191|SY|C2923|NCI_CDISC|Bronchioloalveolar Lung Adenocarcinoma|8251/3
C0007120|T191|PT|C2923|NCI_CDISC|CARCINOMA, BRONCHIOLOALVEOLAR, MALIGNANT|8251/3
C0007120|T191|PT|10058354|NCI_CTEP-SDC|Bronchioloalveolar carcinoma|8251/3
C0007120|T191|DN|C2923|NCI_CTRP|Bronchioloalveolar Carcinoma|8251/3
C0007120|T191|AB|CDR0000043303|PDQ|BAC|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioalveolar Adenocarcinoma of Lung|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioalveolar Adenocarcinoma of the Lung|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioalveolar Lung Carcinoma|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchiolo-Alveolar Carcinoma of Lung|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchiolo-Alveolar Carcinoma of the Lung|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchiolo-Alveolar Lung Carcinoma|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioloalveolar Adenocarcinoma of Lung|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioloalveolar Adenocarcinoma of the Lung|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|bronchioloalveolar carcinoma|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|Bronchioloalveolar Lung Adenocarcinoma|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|bronchoalveolar carcinoma|8251/3
C0007120|T191|PT|CDR0000043303|PDQ|bronchoalveolar cell lung cancer|8251/3
C0007120|T191|SY|CDR0000043303|PDQ|lung cancer, bronchoalveolar cell|8251/3
C0007120|T191|PT|R0121358|QMR|BRONCHIOLAR-ALVEOLAR CELL CARCINOMA|8251/3
C0007120|T191|PT|BB5S4|RCD|Alveolar adenocarcinoma|8251/3
C0007120|T191|SY|BB5S4|RCD|Alveolar carcinoma|8251/3
C0007120|T191|SY|XaBAp|RCD|Alveolar cell carcinoma|8251/3
C0007120|T191|AB|XaBAp|RCD|Bronchio-alveol adenocarc lung|8251/3
C0007120|T191|SY|XaBAp|RCD|Bronchiolar adenocarcinoma|8251/3
C0007120|T191|SY|XaBAp|RCD|Bronchiolar carcinoma|8251/3
C0007120|T191|AB|XaBAp|RCD|Bronchiolo-alveolar adenoca|8251/3
C0007120|T191|SY|XaBAp|RCD|Bronchiolo-alveolar adenocarcinoma|8251/3
C0007120|T191|PT|XaBAp|RCD|Bronchiolo-alveolar adenocarcinoma of lung|8251/3
C0007120|T191|SY|XaBAp|RCD|Bronchiolo-alveolar carcinoma|8251/3
C0007120|T191|SY|XaBAp|RCD|Bronchioloalveolar carcinoma|8251/3
C0007120|T191|AB|BB5S2|RCDSY|Bronchiolo-alveolar adenoca|8251/3
C0007120|T191|PT|BB5S2|RCDSY|Bronchiolo-alveolar adenocarcinoma|8251/3
C0007120|T191|PT|36310008|SNOMEDCT_US|Alveolar adenocarcinoma|8251/3
C0007120|T191|SY|36310008|SNOMEDCT_US|Alveolar carcinoma|8251/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Alveolar cell carcinoma|8251/3
C0007120|T191|SY|112677002|SNOMEDCT_US|Alveolar cell carcinoma|8251/3
C0007120|T191|SY|112677002|SNOMEDCT_US|Bronchiolar adenocarcinoma|8251/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Bronchiolar adenocarcinoma|8251/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Bronchiolar carcinoma|8251/3
C0007120|T191|SY|112677002|SNOMEDCT_US|Bronchiolar carcinoma|8251/3
C0007120|T191|PT|112677002|SNOMEDCT_US|Bronchiolo-alveolar adenocarcinoma|8251/3
C0007120|T191|SY|112677002|SNOMEDCT_US|Bronchiolo-alveolar carcinoma|8251/3
C0007120|T191|OAS|307595008|SNOMEDCT_US|Bronchioloalveolar adenocarcinoma|8251/3
C0007120|T191|OAP|307595008|SNOMEDCT_US|Bronchioloalveolar adenocarcinoma of lung|8251/3
C0007120|T191|OF|307595008|SNOMEDCT_US|Bronchioloalveolar adenocarcinoma of lung|8251/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Bronchioloalveolar carcinoma|8251/3
C0007120|T191|OAP|373627005|SNOMEDCT_US|Bronchioloalveolar carcinoma - disorder|8251/3
C0007120|T191|OAS|373627005|SNOMEDCT_US|Bronchoalveolar cancer|8251/3
C1266034|T191|PT|C7269|NCI|Minimally Invasive Lung Non-Mucinous Adenocarcinoma|8252/3
C1266034|T191|OP|C7269|NCI|Non-Mucinous Bronchioloalveolar Carcinoma|8252/3
C1266034|T191|OP|C7269|NCI|Non-Mucinous Bronchioloalveolar Lung Carcinoma|8252/3
C1266034|T191|OP|C7269|NCI|Non-Mucinous Bronchoalveolar Lung Carcinoma|8252/3
C1266034|T191|SY|C7269|NCI|Non-Mucinous Minimally Invasive Lung Adenocarcinoma|8252/3
C1266034|T191|SY|128659000|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, Clara cell|8252/3
C1266034|T191|PT|128659000|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, non-mucinous|8252/3
C1266034|T191|SY|128659000|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, type II pneumocyte|8252/3
C2200125|T191|PT|219696|MEDCIN|mucinous bronchiolo-alveolar carcinoma of lung|8253/3
C1266035|T191|PN|NOCODE|MTH|Minimally Invasive Mucinous Lung Adenocarcinoma|8253/3
C2200125|T191|PN|NOCODE|MTH|mucinous bronchiolo-alveolar carcinoma of lung|8253/3
C1266035|T191|PT|C7268|NCI|Minimally Invasive Lung Mucinous Adenocarcinoma|8253/3
C1266035|T191|OP|C7268|NCI|Mucinous Bronchioloalveolar Carcinoma|8253/3
C1266035|T191|OP|C7268|NCI|Mucinous Bronchioloalveolar Lung Carcinoma|8253/3
C1266035|T191|OP|C7268|NCI|Mucinous Bronchoalveolar Lung Carcinoma|8253/3
C1266035|T191|SY|C7268|NCI|Mucinous Minimally Invasive Lung Adenocarcinoma|8253/3
C2200125|T191|SY|128660005|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, goblet cell type|8253/3
C2200125|T191|PT|128660005|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, mucinous|8253/3
C1266036|T191|OP|C7270|NCI|Indeterminate Bronchioloalveolar Carcinoma|8254/3
C1266036|T191|OP|C7270|NCI|Mixed Mucinous and Non-Mucinous Bronchioloalveolar Carcinoma|8254/3
C1266036|T191|PT|C7270|NCI|Mixed Mucinous and Non-Mucinous Bronchioloalveolar Carcinoma|8254/3
C1266036|T191|OP|C7270|NCI|Mixed Mucinous and Non-Mucinous Bronchioloalveolar Lung Carcinoma|8254/3
C1266036|T191|OP|C7270|NCI|Mixed Mucinous and Non-Mucinous Bronchoalveolar Lung Carcinoma|8254/3
C1266036|T191|SY|128661009|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, Clara cell and goblet cell type|8254/3
C1266036|T191|SY|128661009|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, indeterminate type|8254/3
C1266036|T191|PT|128661009|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, mixed mucinous and non-mucinous|8254/3
C1266036|T191|SY|128661009|SNOMEDCT_US|Bronchiolo-alveolar carcinoma, type II pneumocyte and goblet cell type|8254/3
C1879591|T191|OP|C65197|NCI|Lung Adenocarcinoma with Mixed Bronchioloalveolar and Invasive Components|8255/3
C1879591|T191|PT|C65197|NCI|Lung Adenocarcinoma with Mixed Bronchioloalveolar and Invasive Components|8255/3
C1879591|T191|SY|90600324|NCI_CTEP-SDC|Lung adenocar. w/ bronch. feat.|8255/3
C1879591|T191|PT|90600324|NCI_CTEP-SDC|Lung adenocarcinoma with bronchioloalveolar features|8255/3
C1266037|T191|SY|128662002|SNOMEDCT_US|Adenocarcinoma combined with other types of carcinoma|8255/3
C1266037|T191|PT|128662002|SNOMEDCT_US|Adenocarcinoma with mixed subtypes|8255/3
C0149845|T191|PT|0060740|CCPSS|BRONCHIAL ADENOMA NOS|8260/0
C0149845|T191|PT|0000016713|CHV|bronchial adenoma|8260/0
C0205650|T191|PT|0000020668|CHV|papillary adenoma|8260/0
C0149845|T191|SY|NOCODE|DXP|BRONCHUS, ADENOMA|8260/0
C0149845|T191|PT|MTHU003485|ICPC2ICD10ENG|adenoma; bronchus|8260/0
C0149845|T191|PT|MTHU012919|ICPC2ICD10ENG|bronchus; adenoma|8260/0
C0205650|T191|PEP|D000236|MSH|Adenoma, Papillary|8260/0
C0205650|T191|PM|D000236|MSH|Adenomas, Papillary|8260/0
C0205650|T191|PM|D000236|MSH|Papillary Adenoma|8260/0
C0205650|T191|PM|D000236|MSH|Papillary Adenomas|8260/0
C0205650|T191|PN|NOCODE|MTH|Papillary adenoma|8260/0
C0149845|T191|SY|C3494|NCI|Adenoma of Bronchus|8260/0
C0149845|T191|SY|C3494|NCI|Adenoma of the Bronchus|8260/0
C0149845|T191|SY|C3494|NCI|Bronchial Adenoma|8260/0
C0149845|T191|PT|C3494|NCI|Lung Papillary Adenoma|8260/0
C0205650|T191|PT|C79951|NCI|Papillary Adenoma|8260/0
C0149845|T191|SY|C3494|NCI|Papillary Adenoma of Type II Pneumocytes|8260/0
C0149845|T191|SY|C3494|NCI|Peripheral Papillary Tumor of Type II Pneumocytes|8260/0
C0149845|T191|SY|C3494|NCI|Type II Pneumocyte Adenoma|8260/0
C0149845|T191|PT|C3494|NCI_CDISC|ADENOMA, BRONCHIAL, BENIGN|8260/0
C0205650|T191|PT|C79951|NCI_CDISC|ADENOMA, PAPILLARY, BENIGN|8260/0
C0149845|T191|PT|CDR0000446531|NCI_NCI-GLOSS|bronchial adenoma|8260/0
C0149845|T191|PT|Xa98a|RCD|Bronchial adenoma|8260/0
C0205650|T191|PT|Xa98b|RCD|Papillary adenoma|8260/0
C0149845|T191|OP|BB5S1|RCDSY|Bronchial adenoma NOS|8260/0
C0205650|T191|OP|BB5T0|RCDSY|Papillary adenoma NOS|8260/0
C0149845|T191|SY|24482001|SNOMEDCT_US|Bronchial adenoma|8260/0
C0149845|T191|IS|24482001|SNOMEDCT_US|Bronchial adenoma, NOS|8260/0
C0205650|T191|PT|86143001|SNOMEDCT_US|Papillary adenoma|8260/0
C0205650|T191|IS|86143001|SNOMEDCT_US|Papillary adenoma, NOS|8260/0
C2348239|T191|SY|HP:0030393|HPO|Aggressive papillary middle ear tumor|8260/1
C2348239|T191|PT|HP:0030393|HPO|Endolymphatic sac tumor|8260/1
C2348239|T191|SY|HP:0030393|HPO|Heffner tumor|8260/1
C2348239|T191|SY|HP:0030393|HPO|Low-grade adenocarcinoma of endolymphatic sac origin|8260/1
C2348239|T191|SY|C67560|NCI|Aggressive Papillary Tumor of the Temporal Bone|8260/1
C2348239|T191|AB|C67560|NCI|ELST|8260/1
C2348239|T191|PT|C67560|NCI|Endolymphatic Sac Tumor|8260/1
C2348239|T191|DN|C67560|NCI_CTRP|Endolymphatic Sac Tumor|8260/1
C2348239|T191|SY|CDR0000729549|PDQ|aggressive papillary tumor of the temporal bone|8260/1
C2348239|T191|AB|CDR0000729549|PDQ|ELST|8260/1
C2348239|T191|PT|CDR0000729549|PDQ|endolymphatic sac tumor|8260/1
C2348239|T191|PT|699817008|SNOMEDCT_US|Endolymphatic sac tumor|8260/1
C2348239|T191|PTGB|699817008|SNOMEDCT_US|Endolymphatic sac tumour|8260/1
C2348239|T191|SY|699817008|SNOMEDCT_US|Neoplasm of endolymphatic sac|8260/1
C0001420|T191|SY|0000000710|CHV|adenocarcinoma papillary|8260/3
C0001420|T191|PT|0000000710|CHV|papillary adenocarcinoma|8260/3
C1306837|T191|PT|0000057924|CHV|papillary renal cell carcinoma|8260/3
C1306837|T191|PT|HP:0006766|HPO|Papillary renal cell carcinoma|8260/3
C0001420|T191|LA|LA26093-7|LNC|Papillary adenocarcinoma|8260/3
C1306837|T191|PT|10078493|MDR|Papillary renal cell carcinoma|8260/3
C1306837|T191|LLT|10078493|MDR|Papillary renal cell carcinoma|8260/3
C0001420|T191|PT|271459|MEDCIN|papillary adenocarcinoma|8260/3
C0001420|T191|MH|D000231|MSH|Adenocarcinoma, Papillary|8260/3
C0001420|T191|PM|D000231|MSH|Adenocarcinomas, Papillary|8260/3
C1306837|T191|ET|D002292|MSH|Chromophil Renal Cell Carcinoma|8260/3
C0001420|T191|PM|D000231|MSH|Papillary Adenocarcinoma|8260/3
C0001420|T191|PM|D000231|MSH|Papillary Adenocarcinomas|8260/3
C1306837|T191|PEP|D002292|MSH|Papillary Renal Cell Carcinoma|8260/3
C1306837|T191|ET|D002292|MSH|Renal Cell Carcinoma, Papillary|8260/3
C0001420|T191|PN|NOCODE|MTH|Papillary adenocarcinoma|8260/3
C1306837|T191|PN|NOCODE|MTH|Papillary Renal Cell Carcinoma|8260/3
C1306837|T191|OP|C6975|NCI|Chromophil Carcinoma of Kidney|8260/3
C1306837|T191|OP|C6975|NCI|Chromophil Carcinoma of the Kidney|8260/3
C1306837|T191|OP|C6975|NCI|Chromophil Renal Cell Carcinoma|8260/3
C0001420|T191|PT|C2853|NCI|Papillary Adenocarcinoma|8260/3
C1306837|T191|PT|C6975|NCI|Papillary Renal Cell Carcinoma|8260/3
C1306837|T191|SY|TCGA|NCI|Papillary Renal Cell Carcinoma|8260/3
C1306837|T191|AB|C6975|NCI|PRCC|8260/3
C0001420|T191|PT|C2853|NCI_CDISC|ADENOCARCINOMA, PAPILLARY, MALIGNANT|8260/3
C1306837|T191|PT|10033702|NCI_CTEP-SDC|Papillary renal cell carcinoma|8260/3
C1306837|T191|DN|C6975|NCI_CTRP|Papillary Renal Cell Cancer|8260/3
C1306837|T191|SY|CDR0000544836|PDQ|Chromophil Carcinoma of Kidney|8260/3
C1306837|T191|SY|CDR0000544836|PDQ|Chromophil Carcinoma of the Kidney|8260/3
C1306837|T191|SY|CDR0000544836|PDQ|Chromophil Renal Cell Carcinoma|8260/3
C1306837|T191|PT|CDR0000544836|PDQ|papillary renal cell carcinoma|8260/3
C0001420|T191|PT|Xa98c|RCD|Papillary adenocarcinoma|8260/3
C0001420|T191|OA|BB5T1|RCDSY|Papillary adenoca. NOS|8260/3
C0001420|T191|OP|BB5T1|RCDSY|Papillary adenocarcinoma NOS|8260/3
C0001420|T191|PT|4797003|SNOMEDCT_US|Papillary adenocarcinoma|8260/3
C0001420|T191|IS|4797003|SNOMEDCT_US|Papillary adenocarcinoma, NOS|8260/3
C1306837|T191|PT|733608000|SNOMEDCT_US|Papillary renal cell carcinoma|8260/3
C1306837|T191|PT|733607005|SNOMEDCT_US|Papillary renal cell carcinoma|8260/3
C1306837|T191|IS|4797003|SNOMEDCT_US|Papillary renal cell carcinoma|8260/3
C0206674|T191|PT|BI00286|BI|villous adenoma|8261/0
C0206674|T191|PT|0018527|CCPSS|ADENOMA VILLOUS|8261/0
C0206674|T191|SY|0000021012|CHV|adenoma villous|8261/0
C0206674|T191|PT|0000021012|CHV|villous adenoma|8261/0
C0206674|T191|SY|0000021012|CHV|villous adenomas|8261/0
C0206674|T191|PT|U000064|COSTAR|VILLOUS ADENOMA|8261/0
C0206674|T191|LA|LA15389-2|LNC|Villous adenoma|8261/0
C0206674|T191|LA|LA26486-3|LNC|Villous adenoma, NOS|8261/0
C0206674|T191|MH|D018253|MSH|Adenoma, Villous|8261/0
C0206674|T191|PM|D018253|MSH|Adenomas, Villous|8261/0
C0206674|T191|PM|D018253|MSH|Villous Adenoma|8261/0
C0206674|T191|PM|D018253|MSH|Villous Adenomas|8261/0
C0206674|T191|PN|NOCODE|MTH|Adenoma, Villous|8261/0
C0206674|T191|PT|C7399|NCI|Villous Adenoma|8261/0
C0206674|T191|PT|CDR0000044809|NCI_NCI-GLOSS|villous adenoma|8261/0
C0206674|T191|PT|Xa98d|RCD|Villous adenoma|8261/0
C0206674|T191|SY|Xa98d|RCD|Villous papilloma|8261/0
C0206674|T191|OP|BB5U0|RCDSY|Villous adenoma NOS|8261/0
C0206674|T191|OAP|67662001|SNOMEDCT_US|Villous adenoma|8261/0
C0206674|T191|PT|128859003|SNOMEDCT_US|Villous adenoma|8261/0
C0206674|T191|IS|67662001|SNOMEDCT_US|Villous adenoma -RETIRED-|8261/0
C0206674|T191|OF|67662001|SNOMEDCT_US|Villous adenoma -RETIRED-|8261/0
C0206674|T191|IS|67662001|SNOMEDCT_US|Villous adenoma, NOS|8261/0
C0206674|T191|IS|67662001|SNOMEDCT_US|Villous papilloma|8261/0
C0206674|T191|SY|128859003|SNOMEDCT_US|Villous papilloma|8261/0
C0334304|T191|PT|271388|MEDCIN|adenocarcinoma in situ in villous adenoma|8261/2
C0334304|T191|PT|C8376|NCI|Adenocarcinoma In Situ in Villous Adenoma|8261/2
C0334304|T191|OA|BB510|RCD|Adenoca situ in villous adenom|8261/2
C0334304|T191|OP|BB510|RCD|Adenocarcinoma in situ in villous adenoma|8261/2
C0334304|T191|OA|BB510|RCDSY|Adenocarc in situ vill aden|8261/2
C0334304|T191|PT|99741000119100|SNOMEDCT_US|Adenocarcinoma in situ in villous adenoma|8261/2
C0334304|T191|PT|4935000|SNOMEDCT_US|Adenocarcinoma in situ in villous adenoma|8261/2
C0334305|T191|PT|271461|MEDCIN|adenocarcinoma in villous adenoma|8261/3
C0334305|T191|PT|C4141|NCI|Adenocarcinoma in Villous Adenoma|8261/3
C0334305|T191|AB|X77nL|RCD|Adenoca in villous adenoma|8261/3
C0334305|T191|PT|X77nL|RCD|Adenocarcinoma in villous adenoma|8261/3
C0334305|T191|OA|BB5U1|RCDSY|Adenoca.in villous adenoma|8261/3
C0334305|T191|OP|BB5U1|RCDSY|Adenocarcinoma in villous adenoma|8261/3
C0334305|T191|OP|BB5Uz|RCDSY|Villous adenoma or adenocarcinoma NOS|8261/3
C0334305|T191|OA|BB5U.|RCDSY|Villous adenoma/ca|8261/3
C0334305|T191|OA|BB5Uz|RCDSY|Villous adenoma/ca NOS|8261/3
C0334305|T191|OP|BB5U.|RCDSY|Villous adenomas and adenocarcinomas|8261/3
C0334305|T191|PT|36087009|SNOMEDCT_US|Adenocarcinoma in villous adenoma|8261/3
C0334305|T191|PT|29431000119108|SNOMEDCT_US|Adenocarcinoma in villous adenoma|8261/3
C0334306|T191|PT|271460|MEDCIN|villous adenocarcinoma|8262/3
C0334306|T191|PT|C4142|NCI|Villous Adenocarcinoma|8262/3
C0334306|T191|PT|BB5U2|RCD|Villous adenocarcinoma|8262/3
C0334306|T191|PT|28558000|SNOMEDCT_US|Villous adenocarcinoma|8262/3
C0334307|T191|PT|0035663|CCPSS|ADENOMA TUBULOVILLOUS|8263/0
C0334307|T191|SY|0000029956|CHV|adenomas tubulovillous|8263/0
C0334307|T191|PT|0000029956|CHV|tubulovillous adenoma|8263/0
C0334307|T191|LA|LA26487-1|LNC|Tubulovillous adenoma, NOS|8263/0
C1708181|T191|PT|39454|MEDCIN|tubulopapillary adenoma of gallbladder|8263/0
C1708181|T191|PT|C43603|NCI|Gallbladder Tubulopapillary Adenoma|8263/0
C0334307|T191|PT|C4143|NCI|Tubulovillous Adenoma|8263/0
C0334307|T191|PT|CDR0000044808|NCI_NCI-GLOSS|tubulovillous adenoma|8263/0
C0334307|T191|SY|BB5U3|RCD|Papillotubular adenoma|8263/0
C0334307|T191|PT|BB5U3|RCD|Tubulovillous adenoma|8263/0
C0334307|T191|SY|BB5U3|RCD|Villoglandular adenoma|8263/0
C0334307|T191|SY|61722000|SNOMEDCT_US|Papillotubular adenoma|8263/0
C0334307|T191|SY|61722000|SNOMEDCT_US|Tubulo-papillary adenoma|8263/0
C0334307|T191|OAP|154632002|SNOMEDCT_US|Tubulovillous adenoma|8263/0
C0334307|T191|OF|154632002|SNOMEDCT_US|Tubulovillous adenoma|8263/0
C0334307|T191|PT|61722000|SNOMEDCT_US|Tubulovillous adenoma|8263/0
C0334307|T191|IS|61722000|SNOMEDCT_US|Tubulovillous adenoma, NOS|8263/0
C0334307|T191|SY|61722000|SNOMEDCT_US|Villoglandular adenoma|8263/0
C0334308|T191|PT|271389|MEDCIN|adenocarcinoma in situ in tubulovillous adenoma|8263/2
C0334308|T191|PT|C4144|NCI|Adenocarcinoma In Situ in Tubulovillous Adenoma|8263/2
C0334308|T191|AB|X77nJ|RCD|Adenoca situ tubulovil adenoma|8263/2
C0334308|T191|PT|X77nJ|RCD|Adenocarcinoma in situ in tubulovillous adenoma|8263/2
C0334308|T191|AB|X77nJ|RCDSY|Adencar in situ tubvil adnm|8263/2
C0334308|T191|OAP|189581002|SNOMEDCT_US|Adenocarcinoma in situ in tubulovillous adenoma|8263/2
C0334308|T191|OF|189581002|SNOMEDCT_US|Adenocarcinoma in situ in tubulovillous adenoma|8263/2
C0334308|T191|PT|51617009|SNOMEDCT_US|Adenocarcinoma in situ in tubulovillous adenoma|8263/2
C0334309|T191|PT|271462|MEDCIN|adenocarcinoma in tubulovillous adenoma|8263/3
C0334309|T191|PT|C4145|NCI|Adenocarcinoma in Tubulovillous Adenoma|8263/3
C0334309|T191|AB|X77nM|RCD|Adenoca in tubulovill adenoma|8263/3
C0334309|T191|PT|X77nM|RCD|Adenocarcinoma in tubulovillous adenoma|8263/3
C0334309|T191|AB|X77nM|RCDSY|Adenocar tubulovil adenoma|8263/3
C0334309|T191|OF|189583004|SNOMEDCT_US|Adenocarcinoma in tubulovillous adenoma|8263/3
C0334309|T191|PT|5658009|SNOMEDCT_US|Adenocarcinoma in tubulovillous adenoma|8263/3
C0334309|T191|OAP|189583004|SNOMEDCT_US|Adenocarcinoma in tubulovillous adenoma|8263/3
C0334309|T191|SY|5658009|SNOMEDCT_US|Papillotubular adenocarcinoma|8263/3
C0334309|T191|SY|5658009|SNOMEDCT_US|Tubulopapillary adenocarcinoma|8263/3
C3839292|T191|PT|703551008|SNOMEDCT_US|Villoglandular carcinoma|8263/3
C1266038|T191|PT|C65198|NCI|Glandular Papillomatosis|8264/0
C1266038|T191|PT|128663007|SNOMEDCT_US|Papillomatosis, glandular|8264/0
C3472608|T191|LA|LA26496-2|LNC|Micropapillary carcinoma|8265/3
C3272815|T191|PT|C96491|NCI|Colorectal Micropapillary Adenocarcinoma|8265/3
C3838947|T191|SY|C36084|NCI|Infiltrating Micropapillary Breast Carcinoma|8265/3
C3838947|T191|PT|C36084|NCI|Invasive Micropapillary Breast Carcinoma|8265/3
C3838947|T191|PT|703578005|SNOMEDCT_US|Invasive micropapillary carcinoma of breast|8265/3
C4518217|T191|PT|733878002|SNOMEDCT_US|Micropapillary adenocarcinoma|8265/3
C3472608|T191|PT|450895005|SNOMEDCT_US|Micropapillary carcinoma|8265/3
C0001432|T191|SY|0000000717|CHV|adenoma chromophobe|8270/0
C0001432|T191|SY|0000000717|CHV|adenoma chromophobe pituitary|8270/0
C0001432|T191|PT|0000000717|CHV|chromophobe adenoma|8270/0
C0001432|T191|MH|D000238|MSH|Adenoma, Chromophobe|8270/0
C0001432|T191|PM|D000238|MSH|Adenomas, Chromophobe|8270/0
C0001432|T191|PM|D000238|MSH|Chromophobe Adenoma|8270/0
C0001432|T191|PM|D000238|MSH|Chromophobe Adenomas|8270/0
C0001432|T191|OP|C2857|NCI|Chromophobe Adenoma|8270/0
C0001432|T191|OP|C2857|NCI|Chromophobe Adenoma of Pituitary Gland|8270/0
C0001432|T191|OP|C2857|NCI|Chromophobe Adenoma of the Pituitary Gland|8270/0
C0001432|T191|OP|C2857|NCI|Pituitary Chromophobe Adenoma|8270/0
C0001432|T191|PT|C2857|NCI|Pituitary Gland Chromophobe Adenoma|8270/0
C0001432|T191|OP|C2857|NCI|Pituitary Gland Chromophobe Adenoma|8270/0
C0001432|T191|DN|C2857|NCI_CTRP|Pituitary Gland Chromophobe Adenoma|8270/0
C0001432|T191|SY|CDR0000040036|PDQ|adenoma, chromophobe, pituitary|8270/0
C0001432|T191|SY|CDR0000040036|PDQ|Chromophobe Adenoma|8270/0
C0001432|T191|SY|CDR0000040036|PDQ|Chromophobe Adenoma of Pituitary Gland|8270/0
C0001432|T191|SY|CDR0000040036|PDQ|Chromophobe Adenoma of the Pituitary Gland|8270/0
C0001432|T191|SY|CDR0000040036|PDQ|chromophobe adenoma, pituitary|8270/0
C0001432|T191|PT|CDR0000040036|PDQ|pituitary chromophobe adenoma|8270/0
C0001432|T191|IS|CDR0000040036|PDQ|Pituitary Gland Chromophobe Adenoma|8270/0
C0001432|T191|PT|BB5V0|RCD|Chromophobe adenoma|8270/0
C0001432|T191|PT|37039006|SNOMEDCT_US|Chromophobe adenoma|8270/0
C1266042|T191|LLT|10080544|MDR|Chromophobe renal cell carcinoma|8270/3
C1266042|T191|PT|10080544|MDR|Chromophobe renal cell carcinoma|8270/3
C1266042|T191|PT|234162|MEDCIN|chromophobe type renal cell carcinoma|8270/3
C1266042|T191|PEP|D002292|MSH|Chromophobe Renal Cell Carcinoma|8270/3
C3887514|T191|PN|NOCODE|MTH|Chromophobe carcinoma|8270/3
C1266042|T191|PN|NOCODE|MTH|Chromophobe Renal Cell Carcinoma|8270/3
C1266042|T191|SY|C4146|NCI|Chromophobe Adenocarcinoma|8270/3
C1266042|T191|SY|C4146|NCI|Chromophobe Carcinoma|8270/3
C1266042|T191|SY|C4146|NCI|Chromophobe Carcinoma of Kidney|8270/3
C1266042|T191|SY|C4146|NCI|Chromophobe Carcinoma of the Kidney|8270/3
C1266042|T191|SY|C4146|NCI|Chromophobe Cell Carcinoma of Kidney|8270/3
C1266042|T191|SY|C4146|NCI|Chromophobe Cell Carcinoma of the Kidney|8270/3
C1266042|T191|PT|C4146|NCI|Chromophobe Renal Cell Carcinoma|8270/3
C1266042|T191|SY|TCGA|NCI|Chromophobe Renal Cell Carcinoma|8270/3
C1266042|T191|SY|C4146|NCI|Renal Cell Carcinoma, Chromophobe Type|8270/3
C1266042|T191|DN|C4146|NCI_CTRP|Chromophobe Renal Cell Cancer|8270/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe adenocarcinoma|8270/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe carcinoma|8270/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe carcinoma of kidney|8270/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe carcinoma of the kidney|8270/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe cell carcinoma of kidney|8270/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe cell carcinoma of the kidney|8270/3
C1266042|T191|PT|CDR0000777276|PDQ|chromophobe renal cell carcinoma|8270/3
C1266042|T191|SY|CDR0000777276|PDQ|renal cell carcinoma, chromophobe type|8270/3
C3887514|T191|SY|BB5V1|RCD|Chromophobe adenocarcinoma|8270/3
C3887514|T191|PT|BB5V1|RCD|Chromophobe carcinoma|8270/3
C3887514|T191|SY|1443001|SNOMEDCT_US|Chromophobe adenocarcinoma|8270/3
C3887514|T191|PT|1443001|SNOMEDCT_US|Chromophobe carcinoma|8270/3
C1266042|T191|SY|128667008|SNOMEDCT_US|Chromophobe cell renal carcinoma|8270/3
C1266042|T191|PT|733471003|SNOMEDCT_US|Chromophobe renal cell carcinoma|8270/3
C1266042|T191|PT|128667008|SNOMEDCT_US|Renal cell carcinoma, chromophobe cell|8270/3
C0033375|T191|PT|1013462|CCPSS|PITUITARY PROLACTINOMA|8271/0
C0033375|T191|PT|0043313|CCPSS|PROLACTINOMA|8271/0
C0033375|T191|SY|0000010174|CHV|adenoma prolactin secreting|8271/0
C0033375|T191|PT|0000047991|CHV|pituitary prolactinoma|8271/0
C0033375|T191|SY|0000047991|CHV|pituitary prolactinomas|8271/0
C0033375|T191|PT|0000010174|CHV|prolactinoma|8271/0
C0033375|T191|SY|0000010174|CHV|prolactinomas|8271/0
C0033375|T191|ET|2006-7421|CSP|prolactinoma|8271/0
C0033375|T191|DI|U001506|DXP|PITUITARY ADENOMA, PROLACTIN SECRETING|8271/0
C0033375|T191|SY|NOCODE|DXP|PROLACTINOMA|8271/0
C0033375|T191|PT|HP:0006767|HPO|Pituitary prolactin cell adenoma|8271/0
C0033375|T191|SY|HP:0006767|HPO|Pituitary prolactinoma|8271/0
C0033375|T191|SY|HP:0006767|HPO|Prolactin-secreting pituitary adenoma|8271/0
C0033375|T191|PT|HP:0040278|HPO|Prolactinoma|8271/0
C0033375|T191|PT|MTHU061947|ICPC2ICD10ENG|prolactinoma; unspecified site|8271/0
C0033375|T191|PT|sh85107392|LCH_NW|Prolactinoma|8271/0
C0033375|T191|LLT|10036832|MDR|Prolactinoma|8271/0
C0033375|T191|SY|30506|MEDCIN|pituitary prolactinoma|8271/0
C0033375|T191|PT|30506|MEDCIN|prolactinoma of pituitary gland|8271/0
C0033375|T191|ET|5328|MEDLINEPLUS|Prolactinoma|8271/0
C0033375|T191|PM|D015175|MSH|Adenoma, Lactotroph|8271/0
C0033375|T191|ET|D015175|MSH|Adenoma, Prolactin-Secreting, Pituitary|8271/0
C0033375|T191|PM|D015175|MSH|Adenomas, Lactotroph|8271/0
C0033375|T191|ET|D015175|MSH|Lactotroph Adenoma|8271/0
C0033375|T191|PM|D015175|MSH|Lactotroph Adenomas|8271/0
C0033375|T191|PM|D015175|MSH|Pituitary Adenoma, PRL-Secreting|8271/0
C0033375|T191|PM|D015175|MSH|Pituitary Adenoma, Prolactin Secreting|8271/0
C0033375|T191|PM|D015175|MSH|Pituitary Adenoma, Prolactin-Producing|8271/0
C0033375|T191|ET|D015175|MSH|Pituitary Adenoma, Prolactin-Secreting|8271/0
C0033375|T191|PM|D015175|MSH|Pituitary Adenomas, PRL-Secreting|8271/0
C0033375|T191|PM|D015175|MSH|Pituitary Adenomas, Prolactin-Producing|8271/0
C0033375|T191|PM|D015175|MSH|Pituitary Adenomas, Prolactin-Secreting|8271/0
C0033375|T191|PM|D015175|MSH|PRL Secreting Pituitary Adenoma|8271/0
C0033375|T191|ET|D015175|MSH|PRL-Secreting Pituitary Adenoma|8271/0
C0033375|T191|PM|D015175|MSH|PRL-Secreting Pituitary Adenomas|8271/0
C0033375|T191|PM|D015175|MSH|Prolactin Producing Pituitary Adenoma|8271/0
C0033375|T191|PM|D015175|MSH|Prolactin Secreting Pituitary Adenoma|8271/0
C0033375|T191|ET|D015175|MSH|Prolactin-Producing Pituitary Adenoma|8271/0
C0033375|T191|PM|D015175|MSH|Prolactin-Producing Pituitary Adenomas|8271/0
C0033375|T191|ET|D015175|MSH|Prolactin-Secreting Pituitary Adenoma|8271/0
C0033375|T191|PM|D015175|MSH|Prolactin-Secreting Pituitary Adenomas|8271/0
C0033375|T191|MH|D015175|MSH|Prolactinoma|8271/0
C0033375|T191|ET|D015175|MSH|Prolactinoma, Familial|8271/0
C0033375|T191|PM|D015175|MSH|Prolactinomas|8271/0
C0033375|T191|PN|NOCODE|MTH|Prolactinoma|8271/0
C0033375|T191|SY|C3342|NCI|Lactotrope Adenoma|8271/0
C0033375|T191|PT|C3342|NCI|Lactotroph Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Lactotroph Cell Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Pituitary Gland Prolactinoma|8271/0
C0033375|T191|SY|C3342|NCI|Pituitary Prolactinoma|8271/0
C0033375|T191|SY|C3342|NCI|PRL Producing Pituitary Gland Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Producing Adenoma of Pituitary|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Producing Adenoma of Pituitary Gland|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Producing Adenoma of the Pituitary|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Producing Adenoma of the Pituitary Gland|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Producing Pituitary Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Producing Pituitary Gland Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Secreting Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Secreting Adenoma of Pituitary|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Secreting Adenoma of Pituitary Gland|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Secreting Adenoma of the Pituitary|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Secreting Adenoma of the Pituitary Gland|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Secreting Pituitary Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin Secreting Pituitary Gland Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Prolactin-Producing Pituitary Gland Adenoma|8271/0
C0033375|T191|SY|C3342|NCI|Prolactinoma|8271/0
C0033375|T191|SY|C3342|NCI|Prolactinoma of Pituitary|8271/0
C0033375|T191|SY|C3342|NCI|Prolactinoma of Pituitary Gland|8271/0
C0033375|T191|SY|C3342|NCI|Prolactinoma of the Pituitary|8271/0
C0033375|T191|SY|C3342|NCI|Prolactinoma of the Pituitary Gland|8271/0
C0033375|T191|DN|C3342|NCI_CTRP|Prolactin-Producing Pituitary Gland Adenoma|8271/0
C0033375|T191|PT|C3342|NCI_NICHD|Prolactinoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|adenoma, prolactin secreting|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Lactotroph Adenoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Pituitary Gland Prolactinoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Pituitary Prolactinoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|PRL Producing Pituitary Gland Adenoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Producing Adenoma of Pituitary|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Producing Adenoma of Pituitary Gland|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Producing Adenoma of the Pituitary|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Producing Adenoma of the Pituitary Gland|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Producing Pituitary Adenoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Producing Pituitary Gland Adenoma|8271/0
C0033375|T191|PT|CDR0000040033|PDQ|prolactin secreting adenoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Secreting Adenoma of Pituitary|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Secreting Adenoma of Pituitary Gland|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Secreting Adenoma of the Pituitary|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Secreting Adenoma of the Pituitary Gland|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Secreting Pituitary Adenoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactin Secreting Pituitary Gland Adenoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactinoma|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactinoma of Pituitary|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactinoma of Pituitary Gland|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactinoma of the Pituitary|8271/0
C0033375|T191|SY|CDR0000040033|PDQ|Prolactinoma of the Pituitary Gland|8271/0
C0033375|T191|PT|R0121734|QMR|PROLACTINOMA|8271/0
C0033375|T191|AB|X77nb|RCD|Prolactin-secret pit adenoma|8271/0
C0033375|T191|SY|X77nb|RCD|Prolactin-secreting pituitary adenoma|8271/0
C0033375|T191|PT|X77nb|RCD|Prolactinoma|8271/0
C0033375|T191|OP|BB5y4|RCDSY|Prolactinoma|8271/0
C0033375|T191|SY|134209002|SNOMEDCT_US|Prolactin-secreting pituitary adenoma|8271/0
C0033375|T191|PT|34337008|SNOMEDCT_US|Prolactinoma|8271/0
C0033375|T191|PT|134209002|SNOMEDCT_US|Prolactinoma|8271/0
C0033375|T191|OAP|367098005|SNOMEDCT_US|Prolactinoma|8271/0
C0033375|T191|OF|134209002|SNOMEDCT_US|Prolactinoma|8271/0
C0033375|T191|OF|367098005|SNOMEDCT_US|Prolactinoma|8271/0
C0032000|T191|PT|0039068|CCPSS|PITUITARY ADENOMA|8272/0
C0032000|T191|SY|0000009757|CHV|adenoma pituitary|8272/0
C0032000|T191|SY|0000009757|CHV|adenomas pituitary|8272/0
C0032000|T191|PT|0000009757|CHV|pituitary adenoma|8272/0
C0032000|T191|PT|584|COSTAR|PITUITARY ADENOMA|8272/0
C0032000|T191|SY|HP:0002893|HPO|Noncancerous tumor in pituitary gland|8272/0
C0032000|T191|PT|HP:0002893|HPO|Pituitary adenoma|8272/0
C0032000|T191|PT|T73010|ICPC2P|Adenoma;pituitary|8272/0
C0032000|T191|PTN|T73010|ICPC2P|pituitary adenoma|8272/0
C0032000|T191|LLT|10035079|MDR|Pituitary adenoma|8272/0
C0032000|T191|PT|354687|MEDCIN|Pituitary adenoma|8272/0
C0032000|T191|PM|D010911|MSH|Adenoma, Pituitary|8272/0
C0032000|T191|PM|D010911|MSH|Adenomas, Pituitary|8272/0
C0032000|T191|PEP|D010911|MSH|Pituitary Adenoma|8272/0
C0032000|T191|PM|D010911|MSH|Pituitary Adenomas|8272/0
C0032000|T191|PN|NOCODE|MTH|Pituitary Adenoma|8272/0
C0032000|T191|SY|C3329|NCI|Adenoma of Pituitary|8272/0
C0032000|T191|SY|C3329|NCI|Adenoma of Pituitary Gland|8272/0
C0032000|T191|SY|C3329|NCI|Adenoma of the Pituitary|8272/0
C0032000|T191|SY|C3329|NCI|Adenoma of the Pituitary Gland|8272/0
C0032000|T191|SY|C3329|NCI|Pituitary Adenoma|8272/0
C0032000|T191|PT|C3329|NCI|Pituitary Gland Adenoma|8272/0
C0032000|T191|SY|C3329|NCI_CDISC|Adenoma of Pituitary|8272/0
C0032000|T191|SY|C3329|NCI_CDISC|Adenoma of Pituitary Gland|8272/0
C0032000|T191|SY|C3329|NCI_CDISC|Adenoma of the Pituitary|8272/0
C0032000|T191|SY|C3329|NCI_CDISC|Adenoma of the Pituitary Gland|8272/0
C0032000|T191|PT|C3329|NCI_CDISC|ADENOMA, ANTERIOR LOBE PITUITARY GLAND, BENIGN|8272/0
C0032000|T191|SY|C3329|NCI_CDISC|Pituitary Adenoma|8272/0
C0032000|T191|PT|C3329|NCI_NICHD|Pituitary Gland Adenoma|8272/0
C0032000|T191|PT|X78aD|RCD|Pituitary adenoma|8272/0
C0032000|T191|OAS|154621002|SNOMEDCT_US|Adenoma - pituitary|8272/0
C0032000|T191|OAS|269643009|SNOMEDCT_US|Adenoma - pituitary|8272/0
C0032000|T191|SY|254956000|SNOMEDCT_US|Adenoma of pituitary|8272/0
C4518348|T191|PT|734037007|SNOMEDCT_US|Ectopic pituitary adenoma|8272/0
C0032000|T191|OAS|189178001|SNOMEDCT_US|Pituitary adenoma|8272/0
C0032000|T191|OAS|269643009|SNOMEDCT_US|Pituitary adenoma|8272/0
C0032000|T191|OAS|154621002|SNOMEDCT_US|Pituitary adenoma|8272/0
C0032000|T191|PT|254956000|SNOMEDCT_US|Pituitary adenoma|8272/0
C0032000|T191|PT|128664001|SNOMEDCT_US|Pituitary adenoma|8272/0
C0032000|T191|OAP|367095008|SNOMEDCT_US|Pituitary adenoma - disorder|8272/0
C0032000|T191|OF|367095008|SNOMEDCT_US|Pituitary adenoma - disorder|8272/0
C0032000|T191|SY|128664001|SNOMEDCT_US|Pituitary adenoma, no ICD-O subtype|8272/0
C0032000|T191|SY|128664001|SNOMEDCT_US|Pituitary adenoma, no International Classification of Diseases for Oncology subtype|8272/0
C0346300|T191|SY|0000031059|CHV|carcinoma pituitary|8272/3
C0346300|T191|PT|0000031059|CHV|pituitary carcinoma|8272/3
C0346300|T191|ET|2006-7421|CSP|pituitary cancer|8272/3
C0346300|T191|PT|HP:0011763|HPO|Pituitary carcinoma|8272/3
C0346300|T191|PT|sh2010009989|LCH_NW|Pituitary gland--Cancer|8272/3
C0346300|T191|PT|30508|MEDCIN|carcinoma of pituitary gland|8272/3
C0346300|T191|SY|30508|MEDCIN|pituitary carcinoma|8272/3
C0346300|T191|ET|D010911|MSH|Cancer of Pituitary|8272/3
C0346300|T191|ET|D010911|MSH|Cancer of the Pituitary|8272/3
C0346300|T191|PM|D010911|MSH|Cancer, Pituitary|8272/3
C0346300|T191|PM|D010911|MSH|Cancers, Pituitary|8272/3
C0346300|T191|PM|D010911|MSH|Carcinoma, Pituitary|8272/3
C0346300|T191|PM|D010911|MSH|Carcinomas, Pituitary|8272/3
C0346300|T191|ET|D010911|MSH|Pituitary Cancer|8272/3
C0346300|T191|PM|D010911|MSH|Pituitary Cancers|8272/3
C0346300|T191|PEP|D010911|MSH|Pituitary Carcinoma|8272/3
C0346300|T191|PM|D010911|MSH|Pituitary Carcinomas|8272/3
C0346300|T191|PN|NOCODE|MTH|Pituitary carcinoma|8272/3
C0346300|T191|SY|C4536|NCI|Cancer of Pituitary|8272/3
C0346300|T191|SY|C4536|NCI|Cancer of Pituitary Gland|8272/3
C0346300|T191|SY|C4536|NCI|Cancer of the Pituitary|8272/3
C0346300|T191|SY|C4536|NCI|Cancer of the Pituitary Gland|8272/3
C0346300|T191|SY|C4536|NCI|Carcinoma of Pituitary|8272/3
C0346300|T191|SY|C4536|NCI|Carcinoma of Pituitary Gland|8272/3
C0346300|T191|SY|C4536|NCI|Carcinoma of the Pituitary|8272/3
C0346300|T191|SY|C4536|NCI|Carcinoma of the Pituitary Gland|8272/3
C0346300|T191|SY|C4536|NCI|Pituitary Carcinoma|8272/3
C0346300|T191|SY|C4536|NCI|Pituitary Gland Adenocarcinoma|8272/3
C0346300|T191|SY|C4536|NCI|Pituitary Gland Cancer|8272/3
C0346300|T191|PT|C4536|NCI|Pituitary Gland Carcinoma|8272/3
C0346300|T191|PT|C4536|NCI_CPTAC|Pituitary Gland Carcinoma|8272/3
C0346300|T191|PT|10035106|NCI_CTEP-SDC|Pituitary gland cancer, NOS|8272/3
C0346300|T191|DN|C4536|NCI_CTRP|Pituitary Gland Cancer|8272/3
C0346300|T191|PT|C4536|NCI_CTRP|Pituitary Gland Carcinoma|8272/3
C0346300|T191|PT|X78aB|RCD|Pituitary carcinoma|8272/3
C0346300|T191|PT|128665000|SNOMEDCT_US|Pituitary carcinoma|8272/3
C0346300|T191|PT|254955001|SNOMEDCT_US|Pituitary carcinoma|8272/3
C0001433|T191|PM|D000239|MSH|Acidophil Adenoma|8280/0
C0001433|T191|PM|D000239|MSH|Acidophil Adenomas|8280/0
C0001433|T191|PM|D000239|MSH|Acidophilic Adenoma|8280/0
C0001433|T191|PM|D000239|MSH|Acidophilic Adenomas|8280/0
C0001433|T191|MH|D000239|MSH|Adenoma, Acidophil|8280/0
C0001433|T191|ET|D000239|MSH|Adenoma, Acidophilic|8280/0
C0001433|T191|ET|D000239|MSH|Adenoma, Eosinophil|8280/0
C0001433|T191|ET|D000239|MSH|Adenoma, Eosinophilic|8280/0
C0001433|T191|PM|D000239|MSH|Adenomas, Acidophil|8280/0
C0001433|T191|PM|D000239|MSH|Adenomas, Acidophilic|8280/0
C0001433|T191|PM|D000239|MSH|Adenomas, Eosinophil|8280/0
C0001433|T191|PM|D000239|MSH|Adenomas, Eosinophilic|8280/0
C0001433|T191|PM|D000239|MSH|Eosinophil Adenoma|8280/0
C0001433|T191|PM|D000239|MSH|Eosinophil Adenomas|8280/0
C0001433|T191|PM|D000239|MSH|Eosinophilic Adenoma|8280/0
C0001433|T191|PM|D000239|MSH|Eosinophilic Adenomas|8280/0
C0001433|T191|OP|C6780|NCI|Acidophil Adenoma|8280/0
C0001433|T191|OP|C6780|NCI|Eosinophil Adenoma|8280/0
C0001433|T191|OP|C6780|NCI|Pituitary Gland Acidophil Adenoma|8280/0
C0001433|T191|PT|C6780|NCI|Pituitary Gland Acidophil Adenoma|8280/0
C0001433|T191|DN|C6780|NCI_CTRP|Pituitary Gland Acidophil Adenoma|8280/0
C0001433|T191|SY|CDR0000040034|PDQ|Acidophil Adenoma|8280/0
C0001433|T191|SY|CDR0000040034|PDQ|adenoma, eosinophilic, pituitary|8280/0
C0001433|T191|SY|CDR0000040034|PDQ|adenoma, growth hormone secreting|8280/0
C0001433|T191|SY|CDR0000040034|PDQ|Eosinophil Adenoma|8280/0
C0001433|T191|SY|CDR0000040034|PDQ|eosinophilic adenoma, pituitary|8280/0
C0001433|T191|SY|CDR0000040034|PDQ|growth hormone secreting adenoma|8280/0
C0001433|T191|SY|CDR0000040034|PDQ|pituitary adenoma, eosinophilic|8280/0
C0001433|T191|PT|CDR0000040034|PDQ|pituitary eosinophilic adenoma|8280/0
C0001433|T191|IS|CDR0000040034|PDQ|Pituitary Gland Acidophil Adenoma|8280/0
C0001433|T191|PT|BB5V2|RCD|Acidophil adenoma|8280/0
C0001433|T191|SY|BB5V2|RCD|Eosinophil adenoma|8280/0
C0001433|T191|PT|21109002|SNOMEDCT_US|Acidophil adenoma|8280/0
C0001433|T191|SY|21109002|SNOMEDCT_US|Eosinophil adenoma|8280/0
C0334311|T191|PT|MTHU002952|ICPC2ICD10ENG|acidophil; carcinoma, unspecified site|8280/3
C0334311|T191|PT|MTHU014725|ICPC2ICD10ENG|carcinoma; acidophil, unspecified site|8280/3
C0334311|T191|PT|236422|MEDCIN|acidophil carcinoma of pituitary gland|8280/3
C0334311|T191|PN|NOCODE|MTH|Acidophil carcinoma|8280/3
C0334311|T191|OP|C4147|NCI|Acidophil Adenocarcinoma|8280/3
C0334311|T191|OP|C4147|NCI|Acidophil Carcinoma|8280/3
C0334311|T191|OP|C4147|NCI|Eosinophil Adenocarcinoma|8280/3
C0334311|T191|OP|C4147|NCI|Eosinophil Carcinoma|8280/3
C0334311|T191|OP|C4147|NCI|Pituitary Gland Acidophil Carcinoma|8280/3
C0334311|T191|PT|C4147|NCI|Pituitary Gland Acidophil Carcinoma|8280/3
C0334311|T191|SY|BB5V3|RCD|Acidophil adenocarcinoma|8280/3
C0334311|T191|PT|BB5V3|RCD|Acidophil carcinoma|8280/3
C0334311|T191|SY|BB5V3|RCD|Eosinophil adenocarcinoma|8280/3
C0334311|T191|SY|BB5V3|RCD|Eosinophil carcinoma|8280/3
C0334311|T191|SY|51217003|SNOMEDCT_US|Acidophil adenocarcinoma|8280/3
C0334311|T191|PT|51217003|SNOMEDCT_US|Acidophil carcinoma|8280/3
C0334311|T191|SY|51217003|SNOMEDCT_US|Eosinophil adenocarcinoma|8280/3
C0334311|T191|SY|51217003|SNOMEDCT_US|Eosinophil carcinoma|8280/3
C0334312|T191|OP|C4148|NCI|Mixed Acidophil-Basophil Adenoma|8281/0
C0334312|T191|OP|C4148|NCI|Mixed Eosinophil-Basophil Adenoma|8281/0
C0334312|T191|OP|C4148|NCI|Pituitary Gland Mixed Acidophil-Basophil Adenoma|8281/0
C0334312|T191|PT|C4148|NCI|Pituitary Gland Mixed Acidophil-Basophil Adenoma|8281/0
C0334312|T191|AB|BB5V4|RCD|Mixed acidoph-basophil adenoma|8281/0
C0334312|T191|PT|BB5V4|RCD|Mixed acidophil-basophil adenoma|8281/0
C0334312|T191|PT|48619006|SNOMEDCT_US|Mixed acidophil-basophil adenoma|8281/0
C0334313|T191|PT|MTHU002954|ICPC2ICD10ENG|acidophil-basophil; carcinoma, unspecified site|8281/3
C0334313|T191|PT|MTHU009798|ICPC2ICD10ENG|basophil-acidophil; carcinoma, unspecified site|8281/3
C0334313|T191|PT|MTHU014726|ICPC2ICD10ENG|carcinoma; acidophil-basophil, unspecified site|8281/3
C0334313|T191|PT|236467|MEDCIN|mixed acidophil-basophil carcinoma of pituitary gland|8281/3
C0334313|T191|OP|C4149|NCI|Mixed Acidophil-Basophil Adenocarcinoma|8281/3
C0334313|T191|OP|C4149|NCI|Mixed Acidophil-Basophil Carcinoma|8281/3
C0334313|T191|OP|C4149|NCI|Mixed Eosinophil-Basophil Carcinoma|8281/3
C0334313|T191|OP|C4149|NCI|Pituitary Gland Mixed Acidophil-Basophil Carcinoma|8281/3
C0334313|T191|PT|C4149|NCI|Pituitary Gland Mixed Acidophil-Basophil Carcinoma|8281/3
C0334313|T191|AB|BB5V5|RCD|Mixed acidophil-basophil ca|8281/3
C0334313|T191|PT|BB5V5|RCD|Mixed acidophil-basophil carcinoma|8281/3
C0334313|T191|PT|23444003|SNOMEDCT_US|Mixed acidophil-basophil carcinoma|8281/3
C1510502|T191|LLT|10048757|MDR|Oncocytoma|8290/0
C1510502|T191|PT|10048757|MDR|Oncocytoma|8290/0
C1510502|T191|LLT|10048760|MDR|Oxyphil adenoma|8290/0
C1510502|T191|MH|D018249|MSH|Adenoma, Oxyphilic|8290/0
C1510502|T191|ET|D018249|MSH|Oncocytoma|8290/0
C1510502|T191|PM|D018249|MSH|Oxyphilic Adenoma|8290/0
C1510502|T191|PN|NOCODE|MTH|Oxyphilic Adenoma|8290/0
C2986561|T191|PN|NOCODE|MTH|Spindle Cell Oncocytoma of the Adenohypophysis|8290/0
C2986561|T191|OP|C94537|NCI|Folliculo-Stellate Cell Tumor of the Pituitary|8290/0
C1510502|T191|PT|C3759|NCI|Oncocytic Adenoma|8290/0
C1510502|T191|SY|C3759|NCI|Oxyphilic Adenoma|8290/0
C2986561|T191|AB|C94537|NCI|SCO|8290/0
C2986561|T191|PT|C94537|NCI|Spindle Cell Oncocytoma|8290/0
C2986561|T191|OP|C94537|NCI|Spindle Cell Oncocytoma of the Adenohypophysis|8290/0
C1510502|T191|SY|BB5W0|RCD|Oncocytic adenoma|8290/0
C1510502|T191|SY|BB5W0|RCD|Oncocytoma|8290/0
C1510502|T191|PT|BB5W0|RCD|Oxyphilic adenoma|8290/0
C1510502|T191|SY|89439007|SNOMEDCT_US|Follicular adenoma, oxyphilic cell|8290/0
C1510502|T191|SY|89439007|SNOMEDCT_US|Oncocytic adenoma|8290/0
C4518222|T191|PT|733886002|SNOMEDCT_US|Oncocytic papillary cystadenoma|8290/0
C1510502|T191|SY|89439007|SNOMEDCT_US|Oncocytoma|8290/0
C1510502|T191|PT|89439007|SNOMEDCT_US|Oxyphilic adenoma|8290/0
C2986561|T191|PT|703844007|SNOMEDCT_US|Spindle cell oncocytoma|8290/0
C0205642|T191|SY|0000020663|CHV|carcinoma oncocytic|8290/3
C0205642|T191|PT|0000020663|CHV|hurthle cell carcinoma|8290/3
C0205642|T191|PT|MTHU003391|ICPC2ICD10ENG|adenocarcinoma; Hurthle cell|8290/3
C0205642|T191|PT|MTHU014767|ICPC2ICD10ENG|carcinoma; Hurthle cell|8290/3
C0205642|T191|PT|MTHU035792|ICPC2ICD10ENG|Hurthle cell; adenocarcinoma|8290/3
C0205642|T191|PT|MTHU035794|ICPC2ICD10ENG|Hurthle cell; carcinoma|8290/3
C0205642|T191|PT|10066136|MDR|Huerthle cell carcinoma|8290/3
C0205642|T191|LLT|10066136|MDR|Huerthle cell carcinoma|8290/3
C0205642|T191|LLT|10080260|MDR|Hurthle cell carcinoma|8290/3
C0205642|T191|LLT|10075558|MDR|Oxyphilic adenocarcinoma|8290/3
C0205642|T191|PT|271478|MEDCIN|oxyphilic adenocarcinoma|8290/3
C0205642|T191|PEP|D000230|MSH|Adenocarcinoma, Oxyphilic|8290/3
C0205642|T191|PM|D000230|MSH|Adenocarcinomas, Oxyphilic|8290/3
C0205642|T191|PM|D000230|MSH|Oxyphilic Adenocarcinoma|8290/3
C0205642|T191|PM|D000230|MSH|Oxyphilic Adenocarcinomas|8290/3
C0205642|T191|SY|C3679|NCI|Hurthle Cell Adenocarcinoma|8290/3
C0205642|T191|SY|C3679|NCI|Hurthle Cell Carcinoma|8290/3
C0205642|T191|SY|C3679|NCI|Oncocytic Adenocarcinoma|8290/3
C0205642|T191|SY|C3679|NCI|Oncocytic Carcinoma|8290/3
C0205642|T191|PT|C3679|NCI|Oxyphilic Adenocarcinoma|8290/3
C0205642|T191|SY|C3679|NCI_CDISC|Hurthle Cell Adenocarcinoma|8290/3
C0205642|T191|SY|C3679|NCI_CDISC|Hurthle Cell Carcinoma|8290/3
C0205642|T191|SY|C3679|NCI_CDISC|Oncocytic Adenocarcinoma|8290/3
C0205642|T191|SY|C3679|NCI_CDISC|Oncocytic Carcinoma|8290/3
C0205642|T191|PT|C3679|NCI_CDISC|ONCOCYTOMA, MALIGNANT|8290/3
C0205642|T191|SY|BB5W1|RCD|Hurthle cell adenocarcinoma|8290/3
C0205642|T191|SY|BB5W1|RCD|Hurthle cell carcinoma|8290/3
C0205642|T191|SY|BB5W1|RCD|Oncocytic adenocarcinoma|8290/3
C0205642|T191|SY|BB5W1|RCD|Oncocytic carcinoma|8290/3
C0205642|T191|PT|BB5W1|RCD|Oxyphilic adenocarcinoma|8290/3
C0205642|T191|SY|57596004|SNOMEDCT_US|Follicular carcinoma, oxyphilic cell|8290/3
C0205642|T191|SY|57596004|SNOMEDCT_US|Hurthle cell adenocarcinoma|8290/3
C0205642|T191|SY|57596004|SNOMEDCT_US|Hurthle cell carcinoma|8290/3
C0205642|T191|SY|57596004|SNOMEDCT_US|Oncocytic adenocarcinoma|8290/3
C0205642|T191|SY|57596004|SNOMEDCT_US|Oncocytic carcinoma|8290/3
C0205642|T191|PT|443261008|SNOMEDCT_US|Oxyphilic adenocarcinoma|8290/3
C0205642|T191|PT|57596004|SNOMEDCT_US|Oxyphilic adenocarcinoma|8290/3
C0001431|T191|MH|D000237|MSH|Adenoma, Basophil|8300/0
C0001431|T191|ET|D000237|MSH|Adenoma, Basophilic|8300/0
C0001431|T191|PM|D000237|MSH|Adenomas, Basophil|8300/0
C0001431|T191|PM|D000237|MSH|Adenomas, Basophilic|8300/0
C0001431|T191|PM|D000237|MSH|Basophil Adenoma|8300/0
C0001431|T191|PM|D000237|MSH|Basophil Adenomas|8300/0
C0001431|T191|PM|D000237|MSH|Basophilic Adenoma|8300/0
C0001431|T191|PM|D000237|MSH|Basophilic Adenomas|8300/0
C0001431|T191|OP|C2856|NCI|Basophilic Adenoma|8300/0
C0001431|T191|OP|C2856|NCI|Basophilic Pituitary Gland Adenoma|8300/0
C0001431|T191|OP|C2856|NCI|Mucoid Cell Adenoma|8300/0
C0001431|T191|OP|C2856|NCI|Pituitary Basophilic Adenoma|8300/0
C0001431|T191|PT|C2856|NCI|Pituitary Gland Basophil Adenoma|8300/0
C0001431|T191|OP|C2856|NCI|Pituitary Gland Basophil Adenoma|8300/0
C0001431|T191|DN|C2856|NCI_CTRP|Pituitary Gland Basophil Adenoma|8300/0
C0001431|T191|SY|CDR0000040031|PDQ|adenoma, basophilic, pituitary|8300/0
C0001431|T191|SY|CDR0000040031|PDQ|Basophilic Adenoma|8300/0
C0001431|T191|SY|CDR0000040031|PDQ|basophilic adenoma, pituitary|8300/0
C0001431|T191|SY|CDR0000040031|PDQ|Basophilic Pituitary Gland Adenoma|8300/0
C0001431|T191|SY|CDR0000040031|PDQ|Mucoid Cell Adenoma|8300/0
C0001431|T191|PT|CDR0000040031|PDQ|pituitary basophilic adenoma|8300/0
C0001431|T191|IS|CDR0000040031|PDQ|Pituitary Gland Basophil Adenoma|8300/0
C0001431|T191|PT|BB5V6|RCD|Basophil adenoma|8300/0
C0001431|T191|SY|BB5V6|RCD|Mucoid cell adenoma|8300/0
C0001431|T191|PT|9436005|SNOMEDCT_US|Basophil adenoma|8300/0
C0001431|T191|SY|9436005|SNOMEDCT_US|Mucoid cell adenoma|8300/0
C0334314|T191|PN|NOCODE|MTH|Basophilic Adenocarcinoma|8300/3
C0334314|T191|PT|C4150|NCI|Basophilic Adenocarcinoma|8300/3
C0334314|T191|SY|C4150|NCI|Basophilic Carcinoma|8300/3
C0334314|T191|SY|BB5V7|RCD|Basophil adenocarcinoma|8300/3
C0334314|T191|PT|BB5V7|RCD|Basophil carcinoma|8300/3
C0334314|T191|SY|BB5V7|RCD|Mucoid cell adenocarcinoma|8300/3
C0334314|T191|SY|47107000|SNOMEDCT_US|Basophil adenocarcinoma|8300/3
C0334314|T191|PT|47107000|SNOMEDCT_US|Basophil carcinoma|8300/3
C0334314|T191|SY|47107000|SNOMEDCT_US|Mucoid cell adenocarcinoma|8300/3
C0334315|T191|PT|C4151|NCI|Clear Cell Adenoma|8310/0
C0334315|T191|PT|C4151|NCI_CDISC|ADENOMA, CLEAR CELL, BENIGN|8310/0
C0334315|T191|PT|BB5X0|RCD|Clear cell adenoma|8310/0
C0334315|T191|PT|1752006|SNOMEDCT_US|Clear cell adenoma|8310/0
C0206681|T191|SY|0000021016|CHV|adenocarcinoma cell clear|8310/3
C0206681|T191|SY|0000021016|CHV|carcinoma cell clear|8310/3
C0206681|T191|SY|0000021016|CHV|carcinoma clear cell|8310/3
C0206681|T191|SY|0000021016|CHV|carcinomas cell clear|8310/3
C0206681|T191|SY|0000021016|CHV|clear cell adenocarcinoma|8310/3
C0206681|T191|PT|0000021016|CHV|clear cell carcinoma|8310/3
C0206681|T191|PT|271475|MEDCIN|clear cell adenocarcinoma|8310/3
C0206681|T191|MH|D018262|MSH|Adenocarcinoma, Clear Cell|8310/3
C0206681|T191|PM|D018262|MSH|Adenocarcinomas, Clear Cell|8310/3
C0206681|T191|PM|D018262|MSH|Clear Cell Adenocarcinoma|8310/3
C0206681|T191|PM|D018262|MSH|Clear Cell Adenocarcinomas|8310/3
C0206681|T191|PT|C36815|NCI|Adenocarcinoma Clear Cell|8310/3
C0206681|T191|PT|C3766|NCI|Clear Cell Adenocarcinoma|8310/3
C0206681|T191|SY|TCGA|NCI|Clear Cell Adenocarcinoma|8310/3
C0206681|T191|SY|C3766|NCI|Clear Cell Carcinoma|8310/3
C0206681|T191|SY|C36815|NCI|Malignant Glandular Clear Cell|8310/3
C0206681|T191|SY|C3766|NCI|Mesonephroid Clear Cell Adenocarcinoma|8310/3
C0206681|T191|SY|C3766|NCI|Mesonephroid Clear Cell Carcinoma|8310/3
C0206681|T191|PT|C3766|NCI_CDISC|ADENOCARCINOMA, CLEAR CELL, MALIGNANT|8310/3
C0206681|T191|SY|C3766|NCI_CDISC|Clear Cell Carcinoma|8310/3
C0206681|T191|SY|C3766|NCI_CDISC|Mesonephroid Clear Cell Adenocarcinoma|8310/3
C0206681|T191|SY|C3766|NCI_CDISC|Mesonephroid Clear Cell Carcinoma|8310/3
C0206681|T191|PT|CDR0000335091|NCI_NCI-GLOSS|clear cell adenocarcinoma|8310/3
C0206681|T191|PT|CDR0000045063|NCI_NCI-GLOSS|clear cell carcinoma|8310/3
C0206681|T191|PT|Xa98e|RCD|Clear cell adenocarcinoma|8310/3
C0206681|T191|SY|Xa98e|RCD|Clear cell carcinoma|8310/3
C0206681|T191|AB|Xa98e|RCD|Mesonephr clear cell adenoca|8310/3
C0206681|T191|SY|Xa98e|RCD|Mesonephroid clear cell adenocarcinoma|8310/3
C0206681|T191|OA|BB5X1|RCDSY|Clear cell adenocarcin NOS|8310/3
C0206681|T191|OP|BB5X1|RCDSY|Clear cell adenocarcinoma NOS|8310/3
C0206681|T191|PT|30546008|SNOMEDCT_US|Clear cell adenocarcinoma|8310/3
C0206681|T191|SY|30546008|SNOMEDCT_US|Clear cell adenocarcinoma, mesonephroid|8310/3
C0206681|T191|IS|30546008|SNOMEDCT_US|Clear cell adenocarcinoma, NOS|8310/3
C0206681|T191|SY|30546008|SNOMEDCT_US|Clear cell carcinoma|8310/3
C0206681|T191|SY|30546008|SNOMEDCT_US|Mesonephroid clear cell adenocarcinoma|8310/3
C0007134|T191|PT|1007858|CCPSS|RENAL CELL CARCINOMA|8311/1
C0007134|T191|SY|0000002435|CHV|adenocarcinoma cells renal|8311/1
C0007134|T191|SY|0000002435|CHV|adenocarcinoma kidneys|8311/1
C0007134|T191|SY|0000002435|CHV|adenocarcinoma of kidney|8311/1
C0007134|T191|SY|0000002435|CHV|adenocarcinoma of the kidney|8311/1
C0007134|T191|SY|0000002435|CHV|adenocarcinoma renal|8311/1
C0007134|T191|SY|0000002435|CHV|cancer cell renal|8311/1
C0007134|T191|SY|0000002435|CHV|cancer cells renal|8311/1
C0007134|T191|SY|0000002435|CHV|carcinoma cell renal|8311/1
C0007134|T191|SY|0000002435|CHV|carcinoma cells renal|8311/1
C0007134|T191|SY|0000002435|CHV|carcinoma kidney|8311/1
C0007134|T191|SY|0000002435|CHV|carcinoma of kidney|8311/1
C0007134|T191|SY|0000002435|CHV|carcinoma renal|8311/1
C0007134|T191|SY|0000002435|CHV|carcinomas renal|8311/1
C0007134|T191|SY|0000002435|CHV|cell renal cancer|8311/1
C0007134|T191|SY|0000002435|CHV|grawitz tumor|8311/1
C0007134|T191|SY|0000002435|CHV|hypernephroid carcinomas|8311/1
C0007134|T191|SY|0000002435|CHV|hypernephroma|8311/1
C0007134|T191|SY|0000002435|CHV|kidney adenocarcinoma|8311/1
C0007134|T191|SY|0000002435|CHV|kidney carcinoma|8311/1
C0007134|T191|SY|0000002435|CHV|of kidney carcinoma|8311/1
C0007134|T191|SY|0000002435|CHV|rcc|8311/1
C0007134|T191|SY|0000002435|CHV|rccs|8311/1
C0007134|T191|SY|0000002435|CHV|renal adenocarcinoma|8311/1
C0007134|T191|SY|0000002435|CHV|renal carcinoma|8311/1
C0007134|T191|SY|0000002435|CHV|renal cell cancer|8311/1
C0007134|T191|PT|0000002435|CHV|renal cell carcinoma|8311/1
C0007134|T191|ET|4003-0049|CSP|adenocarcinoma of kidney|8311/1
C0007134|T191|ET|4003-0049|CSP|RCC|8311/1
C0007134|T191|PT|4003-0049|CSP|renal cell carcinoma|8311/1
C0007134|T191|GT|CARCINOMA|CST|RENAL CARCINOMA|8311/1
C0007134|T191|SY|NOCODE|DXP|RENAL CANCER, ADENOCARCINOMA|8311/1
C0007134|T191|DI|U001659|DXP|RENAL CELL CARCINOMA|8311/1
C0007134|T191|SY|HP:0005584|HPO|Cancer starting in small tubes in kidneys|8311/1
C0007134|T191|SY|HP:0005584|HPO|Hypernephroma|8311/1
C0007134|T191|SY|HP:0005584|HPO|Renal carcinoma|8311/1
C0007134|T191|PT|HP:0005584|HPO|Renal cell carcinoma|8311/1
C0007134|T191|PT|MTHU003411|ICPC2ICD10ENG|adenocarcinoma; renal cell|8311/1
C0007134|T191|PT|MTHU014796|ICPC2ICD10ENG|carcinoma; renal cell|8311/1
C0007134|T191|PT|MTHU053171|ICPC2ICD10ENG|renal cell; adenocarcinoma|8311/1
C0007134|T191|PT|MTHU053172|ICPC2ICD10ENG|renal cell; carcinoma|8311/1
C0007134|T191|PT|U75003|ICPC2P|Carcinoma;kidney|8311/1
C0007134|T191|PTN|U75003|ICPC2P|renal carcinoma|8311/1
C0007134|T191|PT|sh93001433|LCH_NW|Renal cell carcinoma|8311/1
C0007134|T191|LLT|10001174|MDR|Adenocarcinoma of kidney|8311/1
C0007134|T191|LLT|10072444|MDR|Grawitz tumor|8311/1
C0007134|T191|LLT|10072445|MDR|Grawitz tumour|8311/1
C0334316|T191|LLT|10067945|MDR|Hypernephroid tumor|8311/1
C0334316|T191|LLT|10067968|MDR|Hypernephroid tumour|8311/1
C0007134|T191|LLT|10038401|MDR|Renal cell adenocarcinoma|8311/1
C0007134|T191|LLT|10038407|MDR|Renal cell cancer|8311/1
C0007134|T191|PT|10067946|MDR|Renal cell carcinoma|8311/1
C0007134|T191|LLT|10067946|MDR|Renal cell carcinoma|8311/1
C0007134|T191|LLT|10038409|MDR|Renal cell carcinoma NOS|8311/1
C0007134|T191|LLT|10038415|MDR|Renal cell carcinoma stage unspecified|8311/1
C0007134|T191|PT|234168|MEDCIN|adenocarcinoma of kidney|8311/1
C0007134|T191|SY|234168|MEDCIN|renal adenocarcinoma|8311/1
C0007134|T191|PT|31535|MEDCIN|renal cell carcinoma|8311/1
C0007134|T191|ET|D002292|MSH|Adenocarcinoma Of Kidney|8311/1
C0007134|T191|PM|D002292|MSH|Adenocarcinoma Of Kidneys|8311/1
C0007134|T191|ET|D002292|MSH|Adenocarcinoma, Renal|8311/1
C0007134|T191|ET|D002292|MSH|Adenocarcinoma, Renal Cell|8311/1
C0007134|T191|PM|D002292|MSH|Adenocarcinomas, Renal|8311/1
C0007134|T191|PM|D002292|MSH|Adenocarcinomas, Renal Cell|8311/1
C0007134|T191|PM|D002292|MSH|Cancer, Renal Cell|8311/1
C0007134|T191|PM|D002292|MSH|Cancers, Renal Cell|8311/1
C0007134|T191|PM|D002292|MSH|Carcinoma, Nephroid|8311/1
C0007134|T191|MH|D002292|MSH|Carcinoma, Renal Cell|8311/1
C0007134|T191|PM|D002292|MSH|Carcinomas, Nephroid|8311/1
C0007134|T191|PM|D002292|MSH|Carcinomas, Renal Cell|8311/1
C0007134|T191|PM|D002292|MSH|Kidney, Adenocarcinoma Of|8311/1
C0007134|T191|PM|D002292|MSH|Kidneys, Adenocarcinoma Of|8311/1
C0007134|T191|ET|D002292|MSH|Nephroid Carcinoma|8311/1
C0007134|T191|PM|D002292|MSH|Nephroid Carcinomas|8311/1
C0007134|T191|PM|D002292|MSH|Renal Adenocarcinoma|8311/1
C0007134|T191|PM|D002292|MSH|Renal Adenocarcinomas|8311/1
C0007134|T191|PM|D002292|MSH|Renal Cell Adenocarcinoma|8311/1
C0007134|T191|PM|D002292|MSH|Renal Cell Adenocarcinomas|8311/1
C0007134|T191|ET|D002292|MSH|Renal Cell Cancer|8311/1
C0007134|T191|PM|D002292|MSH|Renal Cell Cancers|8311/1
C0007134|T191|ET|D002292|MSH|Renal Cell Carcinoma|8311/1
C0007134|T191|PM|D002292|MSH|Renal Cell Carcinomas|8311/1
C0007134|T191|PN|NOCODE|MTH|Renal Cell Carcinoma|8311/1
C0007134|T191|SY|C9385|NCI|Adenocarcinoma of Kidney|8311/1
C0007134|T191|SY|C9385|NCI|Adenocarcinoma of the Kidney|8311/1
C0007134|T191|SY|C9385|NCI|Kidney Adenocarcinoma|8311/1
C0007134|T191|AB|C9385|NCI|RCC|8311/1
C0007134|T191|SY|C9385|NCI|Renal Cell Adenocarcinoma|8311/1
C0007134|T191|SY|C9385|NCI|Renal Cell Cancer|8311/1
C0007134|T191|PT|C9385|NCI|Renal Cell Carcinoma|8311/1
C0007134|T191|SY|TCGA|NCI|Renal Cell Carcinoma|8311/1
C0007134|T191|SY|C9385|NCI|Renal Cell Carcinoma, Stage Unspecified|8311/1
C0007134|T191|SY|C9385|NCI_CDISC|Adenocarcinoma of Kidney|8311/1
C0007134|T191|SY|C9385|NCI_CDISC|Adenocarcinoma of the Kidney|8311/1
C0007134|T191|PT|C9385|NCI_CDISC|CARCINOMA, RENAL CELL, MALIGNANT|8311/1
C0007134|T191|SY|C9385|NCI_CDISC|Kidney Adenocarcinoma|8311/1
C0007134|T191|SY|C9385|NCI_CDISC|RCC|8311/1
C0007134|T191|SY|C9385|NCI_CDISC|Renal Cell Adenocarcinoma|8311/1
C0007134|T191|SY|C9385|NCI_CDISC|Renal Cell Cancer|8311/1
C0007134|T191|SY|C9385|NCI_CDISC|Renal Cell Carcinoma, Stage Unspecified|8311/1
C0007134|T191|PT|10038415|NCI_CTEP-SDC|Renal cell carcinoma, NOS|8311/1
C0007134|T191|DN|C9385|NCI_CTRP|Renal Cell Cancer|8311/1
C0007134|T191|PT|C9385|NCI_CTRP|Renal Cell Cancer|8311/1
C0007134|T191|SY|C9385|NCI_CTRP|Renal Cell Carcinoma|8311/1
C0007134|T191|PT|CDR0000661353|NCI_NCI-GLOSS|renal cell adenocarcinoma|8311/1
C0007134|T191|PT|CDR0000044988|NCI_NCI-GLOSS|renal cell cancer|8311/1
C0007134|T191|PT|CDR0000661352|NCI_NCI-GLOSS|renal cell carcinoma|8311/1
C0007134|T191|PT|C9385|NCI_NICHD|Renal Cell Carcinoma|8311/1
C0007134|T191|SY|CDR0000039996|PDQ|adenocarcinoma of kidney|8311/1
C0007134|T191|SY|CDR0000039996|PDQ|adenocarcinoma of the kidney|8311/1
C0007134|T191|SY|CDR0000039996|PDQ|kidney adenocarcinoma|8311/1
C0007134|T191|AB|CDR0000039996|PDQ|RCC|8311/1
C0007134|T191|OP|CDR0000039996|PDQ|renal cell adenocarcinoma|8311/1
C0007134|T191|SY|CDR0000039996|PDQ|renal cell carcinoma|8311/1
C0007134|T191|SY|CDR0000039996|PDQ|renal cell carcinoma, stage unspecified|8311/1
C0007134|T191|PT|R0121764|QMR|RENAL CELL CARCINOMA|8311/1
C0007134|T191|SY|X78Yx|RCD|Adenocarcinoma of kidney|8311/1
C0334316|T191|PT|BB5Y.|RCD|Hypernephroid tumour|8311/1
C0007134|T191|SY|X78Yx|RCD|Renal cell adenocarcinoma|8311/1
C0007134|T191|SY|X78Yx|RCD|Renal cell carcinoma|8311/1
C0007134|T191|PT|BB5a0|RCD|Renal cell carcinoma - morphology|8311/1
C0007134|T191|AB|BB5a0|RCD|Renal cell carcinoma-morpholog|8311/1
C0334316|T191|PT|BB5Y.|RCDAE|Hypernephroid tumor|8311/1
C0007134|T191|IS|254915003|SNOMEDCT_US|Adenocarcinoma of kidney|8311/1
C0334316|T191|PT|30713000|SNOMEDCT_US|Hypernephroid tumor|8311/1
C0334316|T191|PTGB|30713000|SNOMEDCT_US|Hypernephroid tumour|8311/1
C0007134|T191|SY|702391001|SNOMEDCT_US|Hypernephroma|8311/1
C0007134|T191|IS|254915003|SNOMEDCT_US|Renal cell adenocarcinoma|8311/1
C0007134|T191|SY|41607009|SNOMEDCT_US|Renal cell adenocarcinoma|8311/1
C0007134|T191|PT|702391001|SNOMEDCT_US|Renal cell carcinoma|8311/1
C0007134|T191|IS|254915003|SNOMEDCT_US|Renal cell carcinoma|8311/1
C0007134|T191|PT|41607009|SNOMEDCT_US|Renal cell carcinoma|8311/1
C0007134|T191|SY|41607009|SNOMEDCT_US|Renal cell carcinoma - morphology|8311/1
C0007134|T191|PT|1007858|CCPSS|RENAL CELL CARCINOMA|8312/3
C0007134|T191|SY|0000002435|CHV|adenocarcinoma cells renal|8312/3
C0007134|T191|SY|0000002435|CHV|adenocarcinoma kidneys|8312/3
C0007134|T191|SY|0000002435|CHV|adenocarcinoma of kidney|8312/3
C0007134|T191|SY|0000002435|CHV|adenocarcinoma of the kidney|8312/3
C0007134|T191|SY|0000002435|CHV|adenocarcinoma renal|8312/3
C0007134|T191|SY|0000002435|CHV|cancer cell renal|8312/3
C0007134|T191|SY|0000002435|CHV|cancer cells renal|8312/3
C0007134|T191|SY|0000002435|CHV|carcinoma cell renal|8312/3
C0007134|T191|SY|0000002435|CHV|carcinoma cells renal|8312/3
C0007134|T191|SY|0000002435|CHV|carcinoma kidney|8312/3
C0007134|T191|SY|0000002435|CHV|carcinoma of kidney|8312/3
C0007134|T191|SY|0000002435|CHV|carcinoma renal|8312/3
C0007134|T191|SY|0000002435|CHV|carcinomas renal|8312/3
C0007134|T191|SY|0000002435|CHV|cell renal cancer|8312/3
C0007134|T191|SY|0000002435|CHV|grawitz tumor|8312/3
C0007134|T191|SY|0000002435|CHV|hypernephroid carcinomas|8312/3
C0007134|T191|SY|0000002435|CHV|hypernephroma|8312/3
C0007134|T191|SY|0000002435|CHV|kidney adenocarcinoma|8312/3
C0007134|T191|SY|0000002435|CHV|kidney carcinoma|8312/3
C0007134|T191|SY|0000002435|CHV|of kidney carcinoma|8312/3
C0007134|T191|SY|0000002435|CHV|rcc|8312/3
C0007134|T191|SY|0000002435|CHV|rccs|8312/3
C0007134|T191|SY|0000002435|CHV|renal adenocarcinoma|8312/3
C0007134|T191|SY|0000002435|CHV|renal carcinoma|8312/3
C0007134|T191|SY|0000002435|CHV|renal cell cancer|8312/3
C0007134|T191|PT|0000002435|CHV|renal cell carcinoma|8312/3
C0007134|T191|ET|4003-0049|CSP|adenocarcinoma of kidney|8312/3
C0007134|T191|ET|4003-0049|CSP|RCC|8312/3
C0007134|T191|PT|4003-0049|CSP|renal cell carcinoma|8312/3
C0007134|T191|GT|CARCINOMA|CST|RENAL CARCINOMA|8312/3
C0007134|T191|SY|NOCODE|DXP|RENAL CANCER, ADENOCARCINOMA|8312/3
C0007134|T191|DI|U001659|DXP|RENAL CELL CARCINOMA|8312/3
C0007134|T191|SY|HP:0005584|HPO|Cancer starting in small tubes in kidneys|8312/3
C0007134|T191|SY|HP:0005584|HPO|Hypernephroma|8312/3
C0007134|T191|SY|HP:0005584|HPO|Renal carcinoma|8312/3
C0007134|T191|PT|HP:0005584|HPO|Renal cell carcinoma|8312/3
C0007134|T191|PT|MTHU003411|ICPC2ICD10ENG|adenocarcinoma; renal cell|8312/3
C0007134|T191|PT|MTHU014796|ICPC2ICD10ENG|carcinoma; renal cell|8312/3
C0007134|T191|PT|MTHU053171|ICPC2ICD10ENG|renal cell; adenocarcinoma|8312/3
C0007134|T191|PT|MTHU053172|ICPC2ICD10ENG|renal cell; carcinoma|8312/3
C0007134|T191|PT|U75003|ICPC2P|Carcinoma;kidney|8312/3
C0007134|T191|PTN|U75003|ICPC2P|renal carcinoma|8312/3
C0007134|T191|PT|sh93001433|LCH_NW|Renal cell carcinoma|8312/3
C0007134|T191|LLT|10001174|MDR|Adenocarcinoma of kidney|8312/3
C0007134|T191|LLT|10072444|MDR|Grawitz tumor|8312/3
C0007134|T191|LLT|10072445|MDR|Grawitz tumour|8312/3
C0007134|T191|LLT|10038401|MDR|Renal cell adenocarcinoma|8312/3
C0007134|T191|LLT|10038407|MDR|Renal cell cancer|8312/3
C0007134|T191|LLT|10067946|MDR|Renal cell carcinoma|8312/3
C0007134|T191|PT|10067946|MDR|Renal cell carcinoma|8312/3
C0007134|T191|LLT|10038409|MDR|Renal cell carcinoma NOS|8312/3
C0007134|T191|LLT|10038415|MDR|Renal cell carcinoma stage unspecified|8312/3
C4049328|T191|LLT|10064886|MDR|Renal medullary carcinoma|8312/3
C0007134|T191|PT|234168|MEDCIN|adenocarcinoma of kidney|8312/3
C4518356|T191|PT|368156|MEDCIN|MiT family translocation renal cell carcinoma|8312/3
C0007134|T191|SY|234168|MEDCIN|renal adenocarcinoma|8312/3
C0007134|T191|PT|31535|MEDCIN|renal cell carcinoma|8312/3
C4518356|T191|SY|368156|MEDCIN|renal malignant carcinoma renal cell, MiT family translocation|8312/3
C0007134|T191|ET|D002292|MSH|Adenocarcinoma Of Kidney|8312/3
C0007134|T191|PM|D002292|MSH|Adenocarcinoma Of Kidneys|8312/3
C0007134|T191|ET|D002292|MSH|Adenocarcinoma, Renal|8312/3
C0007134|T191|ET|D002292|MSH|Adenocarcinoma, Renal Cell|8312/3
C0007134|T191|PM|D002292|MSH|Adenocarcinomas, Renal|8312/3
C0007134|T191|PM|D002292|MSH|Adenocarcinomas, Renal Cell|8312/3
C0007134|T191|PM|D002292|MSH|Cancer, Renal Cell|8312/3
C0007134|T191|PM|D002292|MSH|Cancers, Renal Cell|8312/3
C0007134|T191|PM|D002292|MSH|Carcinoma, Nephroid|8312/3
C0007134|T191|MH|D002292|MSH|Carcinoma, Renal Cell|8312/3
C0007134|T191|PM|D002292|MSH|Carcinomas, Nephroid|8312/3
C0007134|T191|PM|D002292|MSH|Carcinomas, Renal Cell|8312/3
C0007134|T191|PM|D002292|MSH|Kidney, Adenocarcinoma Of|8312/3
C0007134|T191|PM|D002292|MSH|Kidneys, Adenocarcinoma Of|8312/3
C0007134|T191|ET|D002292|MSH|Nephroid Carcinoma|8312/3
C0007134|T191|PM|D002292|MSH|Nephroid Carcinomas|8312/3
C0007134|T191|PM|D002292|MSH|Renal Adenocarcinoma|8312/3
C0007134|T191|PM|D002292|MSH|Renal Adenocarcinomas|8312/3
C0007134|T191|PM|D002292|MSH|Renal Cell Adenocarcinoma|8312/3
C0007134|T191|PM|D002292|MSH|Renal Cell Adenocarcinomas|8312/3
C0007134|T191|ET|D002292|MSH|Renal Cell Cancer|8312/3
C0007134|T191|PM|D002292|MSH|Renal Cell Cancers|8312/3
C0007134|T191|ET|D002292|MSH|Renal Cell Carcinoma|8312/3
C0007134|T191|PM|D002292|MSH|Renal Cell Carcinomas|8312/3
C0007134|T191|PN|NOCODE|MTH|Renal Cell Carcinoma|8312/3
C0007134|T191|SY|C9385|NCI|Adenocarcinoma of Kidney|8312/3
C0007134|T191|SY|C9385|NCI|Adenocarcinoma of the Kidney|8312/3
C0007134|T191|SY|C9385|NCI|Kidney Adenocarcinoma|8312/3
C4049328|T191|PT|C7572|NCI|Kidney Medullary Carcinoma|8312/3
C0007134|T191|AB|C9385|NCI|RCC|8312/3
C0007134|T191|SY|C9385|NCI|Renal Cell Adenocarcinoma|8312/3
C0007134|T191|SY|C9385|NCI|Renal Cell Cancer|8312/3
C0007134|T191|PT|C9385|NCI|Renal Cell Carcinoma|8312/3
C0007134|T191|SY|TCGA|NCI|Renal Cell Carcinoma|8312/3
C0007134|T191|SY|C9385|NCI|Renal Cell Carcinoma, Stage Unspecified|8312/3
C4049328|T191|SY|C7572|NCI|Renal Medullary Carcinoma|8312/3
C0007134|T191|SY|C9385|NCI_CDISC|Adenocarcinoma of Kidney|8312/3
C0007134|T191|SY|C9385|NCI_CDISC|Adenocarcinoma of the Kidney|8312/3
C0007134|T191|PT|C9385|NCI_CDISC|CARCINOMA, RENAL CELL, MALIGNANT|8312/3
C0007134|T191|SY|C9385|NCI_CDISC|Kidney Adenocarcinoma|8312/3
C0007134|T191|SY|C9385|NCI_CDISC|RCC|8312/3
C0007134|T191|SY|C9385|NCI_CDISC|Renal Cell Adenocarcinoma|8312/3
C0007134|T191|SY|C9385|NCI_CDISC|Renal Cell Cancer|8312/3
C0007134|T191|SY|C9385|NCI_CDISC|Renal Cell Carcinoma, Stage Unspecified|8312/3
C0007134|T191|PT|10038415|NCI_CTEP-SDC|Renal cell carcinoma, NOS|8312/3
C0007134|T191|PT|C9385|NCI_CTRP|Renal Cell Cancer|8312/3
C0007134|T191|DN|C9385|NCI_CTRP|Renal Cell Cancer|8312/3
C0007134|T191|SY|C9385|NCI_CTRP|Renal Cell Carcinoma|8312/3
C0007134|T191|PT|CDR0000661353|NCI_NCI-GLOSS|renal cell adenocarcinoma|8312/3
C0007134|T191|PT|CDR0000044988|NCI_NCI-GLOSS|renal cell cancer|8312/3
C0007134|T191|PT|CDR0000661352|NCI_NCI-GLOSS|renal cell carcinoma|8312/3
C0007134|T191|PT|C9385|NCI_NICHD|Renal Cell Carcinoma|8312/3
C0007134|T191|SY|CDR0000039996|PDQ|adenocarcinoma of kidney|8312/3
C0007134|T191|SY|CDR0000039996|PDQ|adenocarcinoma of the kidney|8312/3
C0007134|T191|SY|CDR0000039996|PDQ|kidney adenocarcinoma|8312/3
C0007134|T191|AB|CDR0000039996|PDQ|RCC|8312/3
C0007134|T191|OP|CDR0000039996|PDQ|renal cell adenocarcinoma|8312/3
C0007134|T191|SY|CDR0000039996|PDQ|renal cell carcinoma|8312/3
C0007134|T191|SY|CDR0000039996|PDQ|renal cell carcinoma, stage unspecified|8312/3
C0007134|T191|PT|R0121764|QMR|RENAL CELL CARCINOMA|8312/3
C0007134|T191|SY|X78Yx|RCD|Adenocarcinoma of kidney|8312/3
C0007134|T191|SY|X78Yx|RCD|Renal cell adenocarcinoma|8312/3
C0007134|T191|SY|X78Yx|RCD|Renal cell carcinoma|8312/3
C0007134|T191|PT|BB5a0|RCD|Renal cell carcinoma - morphology|8312/3
C0007134|T191|AB|BB5a0|RCD|Renal cell carcinoma-morpholog|8312/3
C0007134|T191|IS|254915003|SNOMEDCT_US|Adenocarcinoma of kidney|8312/3
C0007134|T191|SY|702391001|SNOMEDCT_US|Hypernephroma|8312/3
C4518356|T191|PT|764694005|SNOMEDCT_US|MiT family translocation renal cell carcinoma|8312/3
C4518356|T191|PT|733881007|SNOMEDCT_US|MiT family translocation renal cell carcinoma|8312/3
C4707257|T191|PT|764990003|SNOMEDCT_US|Mucinous tubular and spindle cell renal carcinoma|8312/3
C0007134|T191|SY|41607009|SNOMEDCT_US|Renal cell adenocarcinoma|8312/3
C0007134|T191|IS|254915003|SNOMEDCT_US|Renal cell adenocarcinoma|8312/3
C0007134|T191|PT|702391001|SNOMEDCT_US|Renal cell carcinoma|8312/3
C0007134|T191|IS|254915003|SNOMEDCT_US|Renal cell carcinoma|8312/3
C0007134|T191|PT|41607009|SNOMEDCT_US|Renal cell carcinoma|8312/3
C0007134|T191|SY|41607009|SNOMEDCT_US|Renal cell carcinoma - morphology|8312/3
C4049328|T191|PT|765094003|SNOMEDCT_US|Renal medullary carcinoma|8312/3
C4049328|T191|PT|765095002|SNOMEDCT_US|Renal medullary carcinoma|8312/3
C4707257|T191|PT|764991004|SNOMEDCT_US|Renal mucinous tubular and spindle cell carcinoma|8312/3
C4707257|T191|SY|764990003|SNOMEDCT_US|Renal mucinous tubular and spindle cell carcinoma|8312/3
C4518356|T191|SY|764694005|SNOMEDCT_US|Translocation renal cell carcinoma|8312/3
C0334317|T191|SY|0000000711|CHV|cystadenofibroma|8313/0
C0334317|T191|SY|0000000711|CHV|cystadenofibromas|8313/0
C0334317|T191|PT|MTHU020306|ICPC2ICD10ENG|cystadenofibroma; unspecified site|8313/0
C0334317|T191|PM|D062625|MSH|Adenofibroma, Clear Cell|8313/0
C0334317|T191|PM|D062625|MSH|Adenofibromas, Clear Cell|8313/0
C0334317|T191|ET|D062625|MSH|Clear Cell Adenofibroma|8313/0
C0334317|T191|PM|D062625|MSH|Clear Cell Adenofibromas|8313/0
C0334317|T191|MH|D062625|MSH|Cystadenofibroma|8313/0
C0334317|T191|PM|D062625|MSH|Cystadenofibromas|8313/0
C0334317|T191|PT|C8987|NCI|Clear Cell Adenofibroma|8313/0
C0334317|T191|PT|C8985|NCI|Cystadenofibroma|8313/0
C0334317|T191|PT|BB5Z.|RCD|Clear cell adenofibroma|8313/0
C0334317|T191|SY|Xa9A5|RCD|Cystadenofibroma|8313/0
C0334317|T191|PT|58161009|SNOMEDCT_US|Clear cell adenofibroma|8313/0
C0334317|T191|SY|2962009|SNOMEDCT_US|Cystadenofibroma|8313/0
C0334317|T191|IS|2962009|SNOMEDCT_US|Cystadenofibroma, NOS|8313/0
C1511258|T191|PT|C40081|NCI|Borderline Ovarian Clear Cell Adenofibroma|8313/1
C1266039|T191|PT|128890001|SNOMEDCT_US|Clear cell adenofibroma of borderline malignancy|8313/1
C1266039|T191|SY|128890001|SNOMEDCT_US|Clear cell borderline tumor|8313/1
C1266039|T191|SYGB|128890001|SNOMEDCT_US|Clear cell borderline tumour|8313/1
C1266039|T191|SY|128890001|SNOMEDCT_US|Clear cell cystadenofibroma of borderline malignancy|8313/1
C1266039|T191|SY|128890001|SNOMEDCT_US|Clear cell tumor, atypical proliferative|8313/1
C1266039|T191|SYGB|128890001|SNOMEDCT_US|Clear cell tumour, atypical proliferative|8313/1
C2075522|T191|PT|233240|MEDCIN|clear cell adenocarcinofibroma of ovary|8313/3
C2075522|T191|PT|C40079|NCI|Ovarian Clear Cell Adenocarcinofibroma|8313/3
C2075522|T191|SY|C40079|NCI|Ovarian Clear Cell Malignant Adenofibroma|8313/3
C1266040|T191|PT|128891002|SNOMEDCT_US|Clear cell adenocarcinofibroma|8313/3
C1266040|T191|SY|128891002|SNOMEDCT_US|Clear cell cystadenocarcinofibroma|8313/3
C0334318|T191|PT|MTHU014788|ICPC2ICD10ENG|carcinoma; lipid-rich|8314/3
C0334318|T191|PT|MTHU045551|ICPC2ICD10ENG|lipid-rich; carcinoma|8314/3
C0334318|T191|PT|C4152|NCI|Lipid-Rich Carcinoma|8314/3
C0334318|T191|PT|C4152|NCI_CPTAC|Lipid-Rich Carcinoma|8314/3
C0334318|T191|PT|X77nG|RCD|Lipid-rich carcinoma|8314/3
C0334318|T191|OF|189655006|SNOMEDCT_US|Lipid-rich carcinoma|8314/3
C0334318|T191|PT|3839000|SNOMEDCT_US|Lipid-rich carcinoma|8314/3
C0334318|T191|OAP|189655006|SNOMEDCT_US|Lipid-rich carcinoma|8314/3
C0334319|T191|PT|C4153|NCI|Glycogen-Rich Carcinoma|8315/3
C0334319|T191|PT|C4153|NCI_CPTAC|Glycogen-Rich Carcinoma|8315/3
C0334319|T191|PT|X77nH|RCD|Glycogen-rich carcinoma|8315/3
C0334319|T191|OAP|189656007|SNOMEDCT_US|Glycogen-rich carcinoma|8315/3
C0334319|T191|OF|189656007|SNOMEDCT_US|Glycogen-rich carcinoma|8315/3
C0334319|T191|PT|74280008|SNOMEDCT_US|Glycogen-rich carcinoma|8315/3
C0334319|T191|SY|74280008|SNOMEDCT_US|Glycogen-rich clear cell carcinoma|8315/3
C1266041|T191|PT|234161|MEDCIN|cyst-associated renal cell carcinoma|8316/3
C0346249|T191|PT|234178|MEDCIN|cystadenocarcinoma of kidney|8316/3
C0346249|T191|OP|C4524|NCI|Multilocular Clear Cell Renal Cell Carcinoma|8316/3
C0346249|T191|PT|C4524|NCI|Multilocular Cystic Renal Neoplasm of Low Malignant Potential|8316/3
C0346249|T191|OP|C4524|NCI|Renal Cystadenocarcinoma|8316/3
C4288091|T191|PT|C126303|NCI|Tubulocystic Renal Cell Carcinoma|8316/3
C0346249|T191|DN|C4524|NCI_CTRP|Multilocular Cystic Renal Cell Cancer|8316/3
C4288091|T191|DN|C126303|NCI_CTRP|Tubulocystic Renal Cell Cancer|8316/3
C0346249|T191|PT|X78Yy|RCD|Cystadenocarcinoma of kidney|8316/3
C1266041|T191|PT|128666004|SNOMEDCT_US|Cyst-associated renal cell carcinoma|8316/3
C0346249|T191|PT|254916002|SNOMEDCT_US|Cystadenocarcinoma of kidney|8316/3
C4518347|T191|PT|734036003|SNOMEDCT_US|Multilocular cystic renal cell neoplasm of low malignant potential|8316/3
C4288091|T191|PT|733602004|SNOMEDCT_US|Tubulocystic renal cell carcinoma|8316/3
C4288091|T191|PT|733603009|SNOMEDCT_US|Tubulocystic renal cell carcinoma|8316/3
C1266042|T191|LLT|10080544|MDR|Chromophobe renal cell carcinoma|8317/3
C1266042|T191|PT|10080544|MDR|Chromophobe renal cell carcinoma|8317/3
C1266042|T191|PT|234162|MEDCIN|chromophobe type renal cell carcinoma|8317/3
C1266042|T191|PEP|D002292|MSH|Chromophobe Renal Cell Carcinoma|8317/3
C1266042|T191|PN|NOCODE|MTH|Chromophobe Renal Cell Carcinoma|8317/3
C1266042|T191|SY|C4146|NCI|Chromophobe Adenocarcinoma|8317/3
C1266042|T191|SY|C4146|NCI|Chromophobe Carcinoma|8317/3
C1266042|T191|SY|C4146|NCI|Chromophobe Carcinoma of Kidney|8317/3
C1266042|T191|SY|C4146|NCI|Chromophobe Carcinoma of the Kidney|8317/3
C1266042|T191|SY|C4146|NCI|Chromophobe Cell Carcinoma of Kidney|8317/3
C1266042|T191|SY|C4146|NCI|Chromophobe Cell Carcinoma of the Kidney|8317/3
C1266042|T191|PT|C4146|NCI|Chromophobe Renal Cell Carcinoma|8317/3
C1266042|T191|SY|TCGA|NCI|Chromophobe Renal Cell Carcinoma|8317/3
C1266042|T191|SY|C4146|NCI|Renal Cell Carcinoma, Chromophobe Type|8317/3
C1266042|T191|DN|C4146|NCI_CTRP|Chromophobe Renal Cell Cancer|8317/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe adenocarcinoma|8317/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe carcinoma|8317/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe carcinoma of kidney|8317/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe carcinoma of the kidney|8317/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe cell carcinoma of kidney|8317/3
C1266042|T191|SY|CDR0000777276|PDQ|chromophobe cell carcinoma of the kidney|8317/3
C1266042|T191|PT|CDR0000777276|PDQ|chromophobe renal cell carcinoma|8317/3
C1266042|T191|SY|CDR0000777276|PDQ|renal cell carcinoma, chromophobe type|8317/3
C1266042|T191|SY|128667008|SNOMEDCT_US|Chromophobe cell renal carcinoma|8317/3
C1266042|T191|PT|733471003|SNOMEDCT_US|Chromophobe renal cell carcinoma|8317/3
C1266042|T191|PT|128667008|SNOMEDCT_US|Renal cell carcinoma, chromophobe cell|8317/3
C1266043|T191|LLT|10066352|MDR|Renal cell carcinoma with sarcomatoid features|8318/3
C1266043|T191|PT|234163|MEDCIN|sarcomatoid renal cell carcinoma|8318/3
C1266043|T191|PEP|D002292|MSH|Sarcomatoid Renal Cell Carcinoma|8318/3
C1266043|T191|PT|C27893|NCI|Sarcomatoid Renal Cell Carcinoma|8318/3
C1266043|T191|SY|10066352|NCI_CTEP-SDC|RCC w/ sarcomatoid features|8318/3
C1266043|T191|PT|10066352|NCI_CTEP-SDC|Renal cell carcinoma with sarcomatoid features|8318/3
C1266043|T191|DN|C27893|NCI_CTRP|Sarcomatoid Renal Cell Cancer|8318/3
C1266043|T191|PT|128668003|SNOMEDCT_US|Renal cell carcinoma, sarcomatoid|8318/3
C1266043|T191|SY|128668003|SNOMEDCT_US|Renal cell carcinoma, spindle cell|8318/3
C1266044|T191|SY|0000056679|CHV|bellini duct carcinoma|8319/3
C1266044|T191|PT|0000056679|CHV|collecting duct carcinoma|8319/3
C1266044|T191|LLT|10073252|MDR|Carcinoma of the collecting ducts of Bellini|8319/3
C1266044|T191|LLT|10066351|MDR|Collecting duct renal cancer|8319/3
C1266044|T191|PT|234164|MEDCIN|collecting duct carcinoma of kidney|8319/3
C1266044|T191|PM|D002292|MSH|Carcinoma, Collecting Duct|8319/3
C1266044|T191|PM|D002292|MSH|Carcinomas, Collecting Duct|8319/3
C1266044|T191|ET|D002292|MSH|Collecting Duct Carcinoma|8319/3
C1266044|T191|ET|D002292|MSH|Collecting Duct Carcinoma of the Kidney|8319/3
C1266044|T191|PM|D002292|MSH|Collecting Duct Carcinomas|8319/3
C1266044|T191|ET|D002292|MSH|Renal Collecting Duct Carcinoma|8319/3
C1266044|T191|PN|NOCODE|MTH|Collecting Duct Carcinoma of the Kidney|8319/3
C1266044|T191|OP|C6194|NCI|Bellini Duct Carcinoma|8319/3
C1266044|T191|SY|C6194|NCI|Carcinoma of Collecting Ducts of Bellini|8319/3
C1266044|T191|SY|C6194|NCI|Carcinoma of Kidney Collecting Duct|8319/3
C1266044|T191|SY|C6194|NCI|Carcinoma of Renal Collecting Duct|8319/3
C1266044|T191|SY|C6194|NCI|Carcinoma of the Collecting Ducts of Bellini|8319/3
C1266044|T191|SY|C6194|NCI|Carcinoma of the Kidney Collecting Duct|8319/3
C1266044|T191|SY|C6194|NCI|Carcinoma of the Renal Collecting Duct|8319/3
C1266044|T191|PT|C6194|NCI|Collecting Duct Carcinoma|8319/3
C1266044|T191|SY|C6194|NCI|Collecting Duct Renal Cell Carcinoma|8319/3
C1266044|T191|SY|C6194|NCI|Kidney Collecting Duct Carcinoma|8319/3
C1266044|T191|SY|C6194|NCI|Renal Collecting Duct Carcinoma|8319/3
C1266044|T191|PT|10066351|NCI_CTEP-SDC|Collecting duct renal cancer|8319/3
C1266044|T191|PT|CDR0000584378|NCI_NCI-GLOSS|BDC|8319/3
C1266044|T191|PT|CDR0000044754|NCI_NCI-GLOSS|Bellini duct carcinoma|8319/3
C1266044|T191|SY|733470002|SNOMEDCT_US|Bellini carcinoma|8319/3
C1266044|T191|SY|733470002|SNOMEDCT_US|Bellini duct carcinoma|8319/3
C1266044|T191|SY|128669006|SNOMEDCT_US|Bellini duct carcinoma|8319/3
C1266044|T191|PT|128669006|SNOMEDCT_US|Collecting duct carcinoma|8319/3
C1266044|T191|PT|733470002|SNOMEDCT_US|Collecting duct carcinoma of kidney|8319/3
C1266044|T191|SY|128669006|SNOMEDCT_US|Renal carcinoma, collecting duct type|8319/3
C1266044|T191|SY|733470002|SNOMEDCT_US|Renal collecting duct carcinoma|8319/3
C0205644|T191|PT|271449|MEDCIN|granular cell carcinoma|8320/3
C0205644|T191|ET|D000230|MSH|Adenocarcinoma, Granular Cell|8320/3
C0205644|T191|PM|D000230|MSH|Adenocarcinomas, Granular Cell|8320/3
C0205644|T191|PEP|D000230|MSH|Carcinoma, Granular Cell|8320/3
C0205644|T191|PM|D000230|MSH|Carcinomas, Granular Cell|8320/3
C0205644|T191|PM|D000230|MSH|Granular Cell Adenocarcinoma|8320/3
C0205644|T191|PM|D000230|MSH|Granular Cell Adenocarcinomas|8320/3
C0205644|T191|PM|D000230|MSH|Granular Cell Carcinoma|8320/3
C0205644|T191|PM|D000230|MSH|Granular Cell Carcinomas|8320/3
C0205644|T191|SY|C3681|NCI|Granular Cell Adenocarcinoma|8320/3
C0205644|T191|PT|C3681|NCI|Granular Cell Carcinoma|8320/3
C0205644|T191|SY|BB5b.|RCD|Granular cell adenocarcinoma|8320/3
C0205644|T191|PT|BB5b.|RCD|Granular cell carcinoma|8320/3
C0205644|T191|SY|69028005|SNOMEDCT_US|Granular cell adenocarcinoma|8320/3
C0205644|T191|PT|69028005|SNOMEDCT_US|Granular cell carcinoma|8320/3
C0334320|T191|PT|0052939|CCPSS|PARATHYROID ADENOMA CHIEF CELL|8321/0
C0334320|T191|PT|MTHU003487|ICPC2ICD10ENG|adenoma; chief cell|8321/0
C0334320|T191|PT|MTHU016136|ICPC2ICD10ENG|chief cell; adenoma|8321/0
C0334320|T191|LLT|10033941|MDR|Parathyroid chief cell adenoma|8321/0
C0334320|T191|SY|C4154|NCI|Chief Cell Adenoma|8321/0
C0334320|T191|SY|C4154|NCI|Chief Cell Adenoma of Parathyroid|8321/0
C0334320|T191|SY|C4154|NCI|Chief Cell Adenoma of Parathyroid Gland|8321/0
C0334320|T191|SY|C4154|NCI|Chief Cell Adenoma of the Parathyroid|8321/0
C0334320|T191|SY|C4154|NCI|Chief Cell Adenoma of the Parathyroid Gland|8321/0
C0334320|T191|SY|C4154|NCI|Parathyroid Chief Cell Adenoma|8321/0
C0334320|T191|PT|C4154|NCI|Parathyroid Gland Chief Cell Adenoma|8321/0
C0334320|T191|DN|C4154|NCI_CTRP|Parathyroid Gland Chief Cell Adenoma|8321/0
C0334320|T191|SY|CDR0000039992|PDQ|Chief Cell Adenoma|8321/0
C0334320|T191|SY|CDR0000039992|PDQ|Chief Cell Adenoma of Parathyroid|8321/0
C0334320|T191|SY|CDR0000039992|PDQ|Chief Cell Adenoma of Parathyroid Gland|8321/0
C0334320|T191|SY|CDR0000039992|PDQ|chief cell adenoma of the parathyroid|8321/0
C0334320|T191|SY|CDR0000039992|PDQ|Chief Cell Adenoma of the Parathyroid Gland|8321/0
C0334320|T191|PT|CDR0000039992|PDQ|parathyroid chief cell adenoma|8321/0
C0334320|T191|SY|CDR0000039992|PDQ|Parathyroid Gland Chief Cell Adenoma|8321/0
C0334320|T191|PT|BB5c0|RCD|Chief cell adenoma|8321/0
C0334320|T191|PT|12205003|SNOMEDCT_US|Chief cell adenoma|8321/0
C0334321|T191|PT|MTHU003530|ICPC2ICD10ENG|adenoma; water-clear cell|8322/0
C0334321|T191|PT|MTHU082134|ICPC2ICD10ENG|water-clear cell; adenoma|8322/0
C0334321|T191|PT|C4155|NCI|Parathyroid Gland Water-Clear Cell Adenoma|8322/0
C0334321|T191|SY|C4155|NCI|Water-Clear Cell Adenoma|8322/0
C0334321|T191|PT|BB5c1|RCD|Water-clear cell adenoma|8322/0
C0334321|T191|PT|26638004|SNOMEDCT_US|Water-clear cell adenoma|8322/0
C0334322|T191|PT|MTHU003423|ICPC2ICD10ENG|adenocarcinoma; water-clear cell|8322/3
C0334322|T191|PT|MTHU014828|ICPC2ICD10ENG|carcinoma; water-clear cell|8322/3
C0334322|T191|PT|MTHU082133|ICPC2ICD10ENG|water-clear cell; adenocarcinoma|8322/3
C0334322|T191|PT|MTHU082135|ICPC2ICD10ENG|water-clear cell; carcinoma|8322/3
C0334322|T191|OP|C4156|NCI|Water-Clear Cell Adenocarcinoma|8322/3
C0334322|T191|PT|C4156|NCI|Water-Clear Cell Adenocarcinoma|8322/3
C0334322|T191|AB|BB5c2|RCD|Water-clear cell adenoca|8322/3
C0334322|T191|PT|BB5c2|RCD|Water-clear cell adenocarcinoma|8322/3
C0334322|T191|SY|BB5c2|RCD|Water-clear cell carcinoma|8322/3
C0334322|T191|PT|80727009|SNOMEDCT_US|Water-clear cell adenocarcinoma|8322/3
C0334322|T191|SY|80727009|SNOMEDCT_US|Water-clear cell carcinoma|8322/3
C0334323|T191|PT|C4157|NCI|Mixed Cell Adenoma|8323/0
C0334323|T191|PT|BB5d0|RCD|Mixed cell adenoma|8323/0
C0334323|T191|PT|89773001|SNOMEDCT_US|Mixed cell adenoma|8323/0
C1332596|T191|PT|C7281|NCI|Borderline Ovarian Seromucinous Tumor/Atypical Proliferative Ovarian Seromucinous Tumor|8323/1
C1302387|T191|PT|399417005|SNOMEDCT_US|Mixed epithelial tumor of borderline malignancy|8323/1
C1302387|T191|PTGB|399417005|SNOMEDCT_US|Mixed epithelial tumour of borderline malignancy|8323/1
C0334324|T191|PT|271479|MEDCIN|mixed cell adenocarcinoma|8323/3
C0334324|T191|OP|C4158|NCI|Mixed Cell Adenocarcinoma|8323/3
C0334324|T191|PT|C4158|NCI|Mixed Cell Adenocarcinoma|8323/3
C0334324|T191|PT|BB5d1|RCD|Mixed cell adenocarcinoma|8323/3
C0334324|T191|PT|38958001|SNOMEDCT_US|Mixed cell adenocarcinoma|8323/3
C0334325|T191|PT|0000029957|CHV|adenolipoma|8324/0
C0334325|T191|SY|0000029957|CHV|lipoadenoma|8324/0
C0334325|T191|LLT|10057341|MDR|Adenolipoma|8324/0
C0334325|T191|PT|10057341|MDR|Adenolipoma|8324/0
C0334325|T191|PT|C4159|NCI|Lipoadenoma|8324/0
C0334325|T191|PT|C4159|NCI_CDISC|ADENOLIPOMA, BENIGN|8324/0
C0334325|T191|SY|BB5e.|RCD|Adenolipoma|8324/0
C0334325|T191|PT|BB5e.|RCD|Lipoadenoma|8324/0
C0334325|T191|SY|22024005|SNOMEDCT_US|Adenolipoma|8324/0
C0334325|T191|PT|22024005|SNOMEDCT_US|Lipoadenoma|8324/0
C1266045|T191|SY|C27253|NCI|Kidney Embryonal Adenoma|8325/0
C1266045|T191|PT|C27253|NCI|Metanephric Adenoma|8325/0
C1266045|T191|PT|128670007|SNOMEDCT_US|Metanephric adenoma|8325/0
C0205647|T191|PT|0056333|CCPSS|ADENOMA FOLLICULAR|8330/0
C0151468|T191|PT|1008962|CCPSS|THYROID ADENOMA|8330/0
C0151468|T191|PT|0050841|CCPSS|THYROID ADENOMA FOLLICULAR|8330/0
C0205647|T191|SY|0000020666|CHV|adenoma follicular|8330/0
C0151468|T191|SY|0000031068|CHV|adenoma follicular thyroid|8330/0
C0151468|T191|SY|0000016975|CHV|adenoma thyroid|8330/0
C0151468|T191|SY|0000016975|CHV|adenomas thyroid|8330/0
C0205647|T191|PT|0000020666|CHV|follicular adenoma|8330/0
C0151468|T191|SY|0000031068|CHV|follicular adenoma thyroid|8330/0
C0151468|T191|PT|0000016975|CHV|thyroid adenoma|8330/0
C0151468|T191|PT|0000031068|CHV|thyroid follicular adenoma|8330/0
C0151468|T191|PT|U000672|COSTAR|THYROID ADENOMA|8330/0
C0151468|T191|GT|ADENOMA THYR|CST|ADENOMA THYROID|8330/0
C0151468|T191|PT|ADENOMA THYR|CST|THYROID ADENOMA|8330/0
C0151468|T191|DI|U001862|DXP|THYROID ADENOMA|8330/0
C0151468|T191|PT|HP:0000854|HPO|Thyroid adenoma|8330/0
C0151468|T191|PT|HP:0011774|HPO|Thyroid follicular adenoma|8330/0
C0151468|T191|PT|T72001|ICPC2P|Adenoma;thyroid|8330/0
C0151468|T191|PTN|T72001|ICPC2P|thyroid adenoma|8330/0
C0151468|T191|LLT|10001237|MDR|Adenoma thyroid|8330/0
C0151468|T191|LLT|10043688|MDR|Thyroid adenoma|8330/0
C0151468|T191|PT|10043688|MDR|Thyroid adenoma|8330/0
C0151468|T191|LLT|10043690|MDR|Thyroid adenoma NOS|8330/0
C0151468|T191|PT|31674|MEDCIN|adenoma of thyroid gland|8330/0
C0151468|T191|PT|38683|MEDCIN|follicular adenoma of thyroid gland|8330/0
C0151468|T191|SY|38683|MEDCIN|follicular thyroid adenoma|8330/0
C0151468|T191|SY|31674|MEDCIN|thyroid adenoma|8330/0
C0205647|T191|PEP|D000236|MSH|Adenoma, Follicular|8330/0
C0151468|T191|PM|D013964|MSH|Adenoma, Thyroid|8330/0
C0205647|T191|PM|D000236|MSH|Adenomas, Follicular|8330/0
C0151468|T191|PM|D013964|MSH|Adenomas, Thyroid|8330/0
C0205647|T191|PM|D000236|MSH|Follicular Adenoma|8330/0
C0205647|T191|PM|D000236|MSH|Follicular Adenomas|8330/0
C0151468|T191|PEP|D013964|MSH|Thyroid Adenoma|8330/0
C0151468|T191|PM|D013964|MSH|Thyroid Adenomas|8330/0
C0205647|T191|PN|NOCODE|MTH|Follicular adenoma|8330/0
C0151468|T191|PN|NOCODE|MTH|Thyroid Gland Follicular Adenoma|8330/0
C0151468|T191|SY|C3502|NCI|Adenoma of the Thyroid|8330/0
C0151468|T191|SY|C3502|NCI|Adenoma of the Thyroid Gland|8330/0
C0151468|T191|SY|C3502|NCI|Adenoma of Thyroid|8330/0
C0151468|T191|SY|C3502|NCI|Adenoma of Thyroid Gland|8330/0
C0151468|T191|SY|C3502|NCI|Follicular Adenoma|8330/0
C0151468|T191|SY|C3502|NCI|Follicular Adenoma of the Thyroid|8330/0
C0151468|T191|SY|C3502|NCI|Follicular Adenoma of the Thyroid Gland|8330/0
C0151468|T191|SY|C3502|NCI|Follicular Adenoma of Thyroid|8330/0
C0151468|T191|SY|C3502|NCI|Follicular Adenoma of Thyroid Gland|8330/0
C0151468|T191|SY|C3502|NCI|Thyroid Adenoma|8330/0
C0151468|T191|SY|C3502|NCI|Thyroid Follicular Adenoma|8330/0
C0151468|T191|SY|C3502|NCI|Thyroid Gland Adenoma|8330/0
C0151468|T191|PT|C3502|NCI|Thyroid Gland Follicular Adenoma|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Adenoma of the Thyroid|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Adenoma of the Thyroid Gland|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Adenoma of Thyroid|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Adenoma of Thyroid Gland|8330/0
C0151468|T191|PT|C3502|NCI_CDISC|ADENOMA, FOLLICULAR CELL, BENIGN|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Follicular Adenoma|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Follicular Adenoma of the Thyroid|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Follicular Adenoma of the Thyroid Gland|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Follicular Adenoma of Thyroid|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Follicular Adenoma of Thyroid Gland|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Thyroid Adenoma|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Thyroid Follicular Adenoma|8330/0
C0151468|T191|SY|C3502|NCI_CDISC|Thyroid Gland Adenoma|8330/0
C0151468|T191|PT|C3502|NCI_NICHD|Thyroid Adenoma|8330/0
C0205647|T191|PT|BB5f0|RCD|Follicular adenoma|8330/0
C0151468|T191|PT|X78cV|RCD|Thyroid adenoma|8330/0
C0151468|T191|PT|X78cW|RCD|Thyroid follicular adenoma|8330/0
C0151468|T191|OAS|189174004|SNOMEDCT_US|Adenoma of thyroid gland|8330/0
C0151468|T191|OAS|154623004|SNOMEDCT_US|Adenoma thyroid gland|8330/0
C0151468|T191|OAS|269644003|SNOMEDCT_US|Adenoma thyroid gland|8330/0
C0205647|T191|PT|55021007|SNOMEDCT_US|Follicular adenoma|8330/0
C0151468|T191|OAS|189174004|SNOMEDCT_US|Thyroid adenoma|8330/0
C0151468|T191|OAS|154623004|SNOMEDCT_US|Thyroid adenoma|8330/0
C0151468|T191|OAS|269644003|SNOMEDCT_US|Thyroid adenoma|8330/0
C0151468|T191|PT|255033000|SNOMEDCT_US|Thyroid adenoma|8330/0
C0151468|T191|PT|255034006|SNOMEDCT_US|Thyroid follicular adenoma|8330/0
C0151468|T191|PT|1100|WHO|THYROID ADENOMA|8330/0
C1266046|T191|SY|C27729|NCI|Atypical Follicular Adenoma|8330/1
C1266046|T191|SY|C27729|NCI|Thyroid Gland Atypical Follicular Adenoma|8330/1
C1266046|T191|SY|C27729|NCI|Thyroid Gland Well-Differentiated Neoplasm of Uncertain Malignant Potential|8330/1
C1266046|T191|PT|C27729|NCI|Thyroid Gland Well-Differentiated Tumor of Uncertain Malignant Potential|8330/1
C1266046|T191|AB|C27729|NCI|WDT-UMP|8330/1
C1266046|T191|PT|128892009|SNOMEDCT_US|Atypical follicular adenoma|8330/1
C0206682|T191|PT|0030530|CCPSS|FOLLICULAR CARCINOMA|8330/3
C0206682|T191|SY|0000016755|CHV|adenocarcinoma thyroid|8330/3
C0206682|T191|SY|0000027295|CHV|cancer follicular thyroid|8330/3
C0206682|T191|SY|0000021017|CHV|carcinoma follicular|8330/3
C0206682|T191|SY|0000016755|CHV|carcinoma follicular thyroid|8330/3
C0206682|T191|SY|0000021017|CHV|carcinomas follicular|8330/3
C0206682|T191|PT|0000021017|CHV|follicular carcinoma|8330/3
C0206682|T191|SY|0000016755|CHV|follicular carcinoma thyroid|8330/3
C0206682|T191|PT|0000027295|CHV|follicular thyroid cancer|8330/3
C0206682|T191|PT|0000016755|CHV|follicular thyroid carcinoma|8330/3
C0206682|T191|SY|0000027295|CHV|thyroid follicular cancer|8330/3
C0206682|T191|SY|0000016755|CHV|thyroid follicular carcinoma|8330/3
C0206682|T191|SY|NOCODE|DXP|THYROID CANCER, FOLLICULAR CARCINOMA|8330/3
C0206682|T191|DI|U001866|DXP|THYROID, CARCINOMA, FOLLICULAR|8330/3
C0206682|T191|PT|HP:0006731|HPO|Follicular thyroid carcinoma|8330/3
C0206682|T191|PT|MTHU003385|ICPC2ICD10ENG|adenocarcinoma; follicular, well differentiated|8330/3
C0206682|T191|PT|MTHU014757|ICPC2ICD10ENG|carcinoma; follicular, pure|8330/3
C0206682|T191|PT|MTHU014753|ICPC2ICD10ENG|carcinoma; follicular, well differentiated|8330/3
C0206682|T191|PT|MTHU029186|ICPC2ICD10ENG|follicular; adenocarcinoma, well differentiated|8330/3
C0206682|T191|PT|MTHU029191|ICPC2ICD10ENG|follicular; carcinoma, well differentiated|8330/3
C0206682|T191|PT|31676|MEDCIN|follicular adenocarcinoma of thyroid gland|8330/3
C0206682|T191|PT|351571|MEDCIN|follicular thyroid carcinoma|8330/3
C0206682|T191|SY|351571|MEDCIN|thyroid malignant carcinoma follicualr|8330/3
C0206682|T191|MH|D018263|MSH|Adenocarcinoma, Follicular|8330/3
C0206682|T191|PM|D018263|MSH|Adenocarcinomas, Follicular|8330/3
C0206682|T191|PM|D018263|MSH|Carcinoma, Follicular Thyroid|8330/3
C0206682|T191|PM|D018263|MSH|Carcinomas, Follicular Thyroid|8330/3
C0206682|T191|PM|D018263|MSH|Follicular Adenocarcinoma|8330/3
C0206682|T191|PM|D018263|MSH|Follicular Adenocarcinomas|8330/3
C0206682|T191|ET|D018263|MSH|Follicular Thyroid Carcinoma|8330/3
C0206682|T191|PM|D018263|MSH|Follicular Thyroid Carcinomas|8330/3
C0206682|T191|ET|D018263|MSH|Thyroid Carcinoma, Follicular|8330/3
C0206682|T191|PM|D018263|MSH|Thyroid Carcinomas, Follicular|8330/3
C0206682|T191|PN|NOCODE|MTH|Follicular thyroid carcinoma|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Adenocarcinoma|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Cancer of the Thyroid|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Cancer of the Thyroid Gland|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Cancer of Thyroid|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Cancer of Thyroid Gland|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma of the Thyroid|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma of the Thyroid Gland|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma of Thyroid|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma of Thyroid Gland|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Thyroid Cancer|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Thyroid Carcinoma|8330/3
C0206682|T191|SY|C8054|NCI|Follicular Thyroid Gland Carcinoma|8330/3
C0206682|T191|AB|C8054|NCI|FTC|8330/3
C0206682|T191|SY|C8054|NCI|Thyroid Follicular Carcinoma|8330/3
C0206682|T191|PT|C8054|NCI|Thyroid Gland Follicular Carcinoma|8330/3
C0206682|T191|SY|C8054|NCI|Well-Differentiated Follicular Adenocarcinoma|8330/3
C0206682|T191|SY|C8054|NCI|Well-Differentiated Follicular Carcinoma|8330/3
C0206682|T191|PT|C8054|NCI_CDISC|CARCINOMA, FOLLICULAR CELL, MALIGNANT|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Adenocarcinoma|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Cancer of the Thyroid|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Cancer of the Thyroid Gland|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Cancer of Thyroid|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Cancer of Thyroid Gland|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma of the Thyroid|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma of the Thyroid Gland|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma of Thyroid|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma of Thyroid Gland|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Thyroid Cancer|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Thyroid Carcinoma|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Thyroid Gland Carcinoma|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Thyroid Follicular Carcinoma|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Well-differentiated Follicular Adenocarcinoma|8330/3
C0206682|T191|SY|C8054|NCI_CDISC|Well-differentiated Follicular Carcinoma|8330/3
C0206682|T191|PT|10016935|NCI_CTEP-SDC|Follicular thyroid carcinoma|8330/3
C0206682|T191|DN|C8054|NCI_CTRP|Thyroid Gland Follicular Cancer|8330/3
C0206682|T191|PT|CDR0000044544|NCI_NCI-GLOSS|follicular thyroid cancer|8330/3
C0206682|T191|PT|C8054|NCI_NICHD|Follicular Thyroid Carcinoma|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Adenocarcinoma|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma of the Thyroid|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma of the Thyroid Gland|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma of Thyroid|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma of Thyroid Gland|8330/3
C0206682|T191|PT|CDR0000040218|PDQ|follicular thyroid cancer|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Thyroid Carcinoma|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Thyroid Gland Carcinoma|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Thyroid Follicular Carcinoma|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Thyroid Gland Follicular Carcinoma|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Well-Differentiated Follicular Adenocarcinoma|8330/3
C0206682|T191|SY|CDR0000040218|PDQ|Well-Differentiated Follicular Carcinoma|8330/3
C0206682|T191|PT|R0121929|QMR|THYROID FOLLICULAR CARCINOMA|8330/3
C0206682|T191|AB|BB5f2|RCD|Follicular adenoca - well diff|8330/3
C0206682|T191|PT|Xa98P|RCD|Follicular adenocarcinoma|8330/3
C0206682|T191|PT|BB5f2|RCD|Follicular adenocarcinoma - well differentiated|8330/3
C0206682|T191|AB|BB5f2|RCD|Follicular ca - well diff|8330/3
C0206682|T191|SY|Xa98P|RCD|Follicular carcinoma|8330/3
C0206682|T191|SY|BB5f2|RCD|Follicular carcinoma - well differentiated|8330/3
C0206682|T191|PT|X78cP|RCD|Follicular thyroid carcinoma|8330/3
C0206682|T191|AB|X78cP|RCD|FTC - Follicular thyroid carc|8330/3
C0206682|T191|SY|X78cP|RCD|FTC - Follicular thyroid carcinoma|8330/3
C0206682|T191|OA|BB5f1|RCDSY|Follicular adenocarc.NOS|8330/3
C0206682|T191|OP|BB5f1|RCDSY|Follicular adenocarcinoma NOS|8330/3
C0206682|T191|PT|5257006|SNOMEDCT_US|Follicular adenocarcinoma|8330/3
C0206682|T191|SY|28173006|SNOMEDCT_US|Follicular adenocarcinoma - well differentiated|8330/3
C0206682|T191|IS|5257006|SNOMEDCT_US|Follicular adenocarcinoma, NOS|8330/3
C0206682|T191|PT|28173006|SNOMEDCT_US|Follicular adenocarcinoma, well differentiated|8330/3
C0206682|T191|SY|5257006|SNOMEDCT_US|Follicular carcinoma|8330/3
C0206682|T191|SY|28173006|SNOMEDCT_US|Follicular carcinoma - well differentiated|8330/3
C1720506|T191|PT|421686008|SNOMEDCT_US|Follicular carcinoma, clear cell|8330/3
C0206682|T191|IS|5257006|SNOMEDCT_US|Follicular carcinoma, NOS|8330/3
C0206682|T191|SY|28173006|SNOMEDCT_US|Follicular carcinoma, well differentiated|8330/3
C1720470|T191|PT|420301000|SNOMEDCT_US|Follicular carcinoma, widely invasive|8330/3
C0206682|T191|PT|255028004|SNOMEDCT_US|Follicular thyroid carcinoma|8330/3
C0206682|T191|IS|255028004|SNOMEDCT_US|FTC - Follicular thyroid carcinoma|8330/3
C0206682|T191|SY|255028004|SNOMEDCT_US|FTC - follicular thyroid carcinoma|8330/3
C0206682|T191|PT|0030530|CCPSS|FOLLICULAR CARCINOMA|8331/3
C0206682|T191|SY|0000016755|CHV|adenocarcinoma thyroid|8331/3
C0206682|T191|SY|0000027295|CHV|cancer follicular thyroid|8331/3
C0206682|T191|SY|0000021017|CHV|carcinoma follicular|8331/3
C0206682|T191|SY|0000016755|CHV|carcinoma follicular thyroid|8331/3
C0206682|T191|SY|0000021017|CHV|carcinomas follicular|8331/3
C0206682|T191|PT|0000021017|CHV|follicular carcinoma|8331/3
C0206682|T191|SY|0000016755|CHV|follicular carcinoma thyroid|8331/3
C0206682|T191|PT|0000027295|CHV|follicular thyroid cancer|8331/3
C0206682|T191|PT|0000016755|CHV|follicular thyroid carcinoma|8331/3
C0206682|T191|SY|0000027295|CHV|thyroid follicular cancer|8331/3
C0206682|T191|SY|0000016755|CHV|thyroid follicular carcinoma|8331/3
C0206682|T191|SY|NOCODE|DXP|THYROID CANCER, FOLLICULAR CARCINOMA|8331/3
C0206682|T191|DI|U001866|DXP|THYROID, CARCINOMA, FOLLICULAR|8331/3
C0206682|T191|PT|HP:0006731|HPO|Follicular thyroid carcinoma|8331/3
C0206682|T191|PT|MTHU003385|ICPC2ICD10ENG|adenocarcinoma; follicular, well differentiated|8331/3
C0206682|T191|PT|MTHU014757|ICPC2ICD10ENG|carcinoma; follicular, pure|8331/3
C0206682|T191|PT|MTHU014753|ICPC2ICD10ENG|carcinoma; follicular, well differentiated|8331/3
C0206682|T191|PT|MTHU029186|ICPC2ICD10ENG|follicular; adenocarcinoma, well differentiated|8331/3
C0206682|T191|PT|MTHU029191|ICPC2ICD10ENG|follicular; carcinoma, well differentiated|8331/3
C0206682|T191|PT|31676|MEDCIN|follicular adenocarcinoma of thyroid gland|8331/3
C0206682|T191|PT|351571|MEDCIN|follicular thyroid carcinoma|8331/3
C0206682|T191|SY|351571|MEDCIN|thyroid malignant carcinoma follicualr|8331/3
C0206682|T191|MH|D018263|MSH|Adenocarcinoma, Follicular|8331/3
C0206682|T191|PM|D018263|MSH|Adenocarcinomas, Follicular|8331/3
C0206682|T191|PM|D018263|MSH|Carcinoma, Follicular Thyroid|8331/3
C0206682|T191|PM|D018263|MSH|Carcinomas, Follicular Thyroid|8331/3
C0206682|T191|PM|D018263|MSH|Follicular Adenocarcinoma|8331/3
C0206682|T191|PM|D018263|MSH|Follicular Adenocarcinomas|8331/3
C0206682|T191|ET|D018263|MSH|Follicular Thyroid Carcinoma|8331/3
C0206682|T191|PM|D018263|MSH|Follicular Thyroid Carcinomas|8331/3
C0206682|T191|ET|D018263|MSH|Thyroid Carcinoma, Follicular|8331/3
C0206682|T191|PM|D018263|MSH|Thyroid Carcinomas, Follicular|8331/3
C0206682|T191|PN|NOCODE|MTH|Follicular thyroid carcinoma|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Adenocarcinoma|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Cancer of the Thyroid|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Cancer of the Thyroid Gland|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Cancer of Thyroid|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Cancer of Thyroid Gland|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma of the Thyroid|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma of the Thyroid Gland|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma of Thyroid|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Carcinoma of Thyroid Gland|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Thyroid Cancer|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Thyroid Carcinoma|8331/3
C0206682|T191|SY|C8054|NCI|Follicular Thyroid Gland Carcinoma|8331/3
C0206682|T191|AB|C8054|NCI|FTC|8331/3
C0206682|T191|SY|C8054|NCI|Thyroid Follicular Carcinoma|8331/3
C0206682|T191|PT|C8054|NCI|Thyroid Gland Follicular Carcinoma|8331/3
C0206682|T191|SY|C8054|NCI|Well-Differentiated Follicular Adenocarcinoma|8331/3
C0206682|T191|SY|C8054|NCI|Well-Differentiated Follicular Carcinoma|8331/3
C0206682|T191|PT|C8054|NCI_CDISC|CARCINOMA, FOLLICULAR CELL, MALIGNANT|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Adenocarcinoma|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Cancer of the Thyroid|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Cancer of the Thyroid Gland|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Cancer of Thyroid|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Cancer of Thyroid Gland|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma of the Thyroid|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma of the Thyroid Gland|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma of Thyroid|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Carcinoma of Thyroid Gland|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Thyroid Cancer|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Thyroid Carcinoma|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Follicular Thyroid Gland Carcinoma|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Thyroid Follicular Carcinoma|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Well-differentiated Follicular Adenocarcinoma|8331/3
C0206682|T191|SY|C8054|NCI_CDISC|Well-differentiated Follicular Carcinoma|8331/3
C0206682|T191|PT|10016935|NCI_CTEP-SDC|Follicular thyroid carcinoma|8331/3
C0206682|T191|DN|C8054|NCI_CTRP|Thyroid Gland Follicular Cancer|8331/3
C0206682|T191|PT|CDR0000044544|NCI_NCI-GLOSS|follicular thyroid cancer|8331/3
C0206682|T191|PT|C8054|NCI_NICHD|Follicular Thyroid Carcinoma|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Adenocarcinoma|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma of the Thyroid|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma of the Thyroid Gland|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma of Thyroid|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Carcinoma of Thyroid Gland|8331/3
C0206682|T191|PT|CDR0000040218|PDQ|follicular thyroid cancer|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Thyroid Carcinoma|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Follicular Thyroid Gland Carcinoma|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Thyroid Follicular Carcinoma|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Thyroid Gland Follicular Carcinoma|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Well-Differentiated Follicular Adenocarcinoma|8331/3
C0206682|T191|SY|CDR0000040218|PDQ|Well-Differentiated Follicular Carcinoma|8331/3
C0206682|T191|PT|R0121929|QMR|THYROID FOLLICULAR CARCINOMA|8331/3
C0206682|T191|AB|BB5f2|RCD|Follicular adenoca - well diff|8331/3
C0206682|T191|PT|Xa98P|RCD|Follicular adenocarcinoma|8331/3
C0206682|T191|PT|BB5f2|RCD|Follicular adenocarcinoma - well differentiated|8331/3
C0206682|T191|AB|BB5f2|RCD|Follicular ca - well diff|8331/3
C0206682|T191|SY|Xa98P|RCD|Follicular carcinoma|8331/3
C0206682|T191|SY|BB5f2|RCD|Follicular carcinoma - well differentiated|8331/3
C0206682|T191|PT|X78cP|RCD|Follicular thyroid carcinoma|8331/3
C0206682|T191|AB|X78cP|RCD|FTC - Follicular thyroid carc|8331/3
C0206682|T191|SY|X78cP|RCD|FTC - Follicular thyroid carcinoma|8331/3
C0206682|T191|OA|BB5f1|RCDSY|Follicular adenocarc.NOS|8331/3
C0206682|T191|OP|BB5f1|RCDSY|Follicular adenocarcinoma NOS|8331/3
C0206682|T191|PT|5257006|SNOMEDCT_US|Follicular adenocarcinoma|8331/3
C0206682|T191|SY|28173006|SNOMEDCT_US|Follicular adenocarcinoma - well differentiated|8331/3
C0206682|T191|IS|5257006|SNOMEDCT_US|Follicular adenocarcinoma, NOS|8331/3
C0206682|T191|PT|28173006|SNOMEDCT_US|Follicular adenocarcinoma, well differentiated|8331/3
C0206682|T191|SY|5257006|SNOMEDCT_US|Follicular carcinoma|8331/3
C0206682|T191|SY|28173006|SNOMEDCT_US|Follicular carcinoma - well differentiated|8331/3
C0206682|T191|IS|5257006|SNOMEDCT_US|Follicular carcinoma, NOS|8331/3
C0206682|T191|SY|28173006|SNOMEDCT_US|Follicular carcinoma, well differentiated|8331/3
C0206682|T191|PT|255028004|SNOMEDCT_US|Follicular thyroid carcinoma|8331/3
C0206682|T191|IS|255028004|SNOMEDCT_US|FTC - Follicular thyroid carcinoma|8331/3
C0206682|T191|SY|255028004|SNOMEDCT_US|FTC - follicular thyroid carcinoma|8331/3
C0334327|T191|PT|MTHU003388|ICPC2ICD10ENG|adenocarcinoma; follicular, trabecular|8332/3
C0334327|T191|PT|MTHU003422|ICPC2ICD10ENG|adenocarcinoma; trabecular follicular|8332/3
C0334327|T191|PT|MTHU014756|ICPC2ICD10ENG|carcinoma; follicular, trabecular|8332/3
C0334327|T191|PT|MTHU014827|ICPC2ICD10ENG|carcinoma; trabecular, follicular|8332/3
C0334327|T191|PT|MTHU029189|ICPC2ICD10ENG|follicular; adenocarcinoma, trabecular|8332/3
C0334327|T191|PT|MTHU029195|ICPC2ICD10ENG|follicular; carcinoma, trabecular|8332/3
C0334327|T191|PT|MTHU042863|ICPC2ICD10ENG|Langhans; wuchernde Struma|8332/3
C0334327|T191|PT|MTHU074798|ICPC2ICD10ENG|trabecular; follicular adenocarcinoma|8332/3
C0334327|T191|PT|MTHU082488|ICPC2ICD10ENG|wuchernde Struma Langhans|8332/3
C0302182|T191|PT|271476|MEDCIN|trabecular adenocarcinoma|8332/3
C0334327|T191|PN|NOCODE|MTH|Trabecular Follicular Adenocarcinoma|8332/3
C0302182|T191|PT|C4068|NCI|Trabecular Adenocarcinoma|8332/3
C0302182|T191|SY|C4068|NCI|Trabecular Carcinoma|8332/3
C0334327|T191|AB|BB5f3|RCD|Follicular adenoca - mod diff|8332/3
C0334327|T191|AB|BB5f3|RCD|Follicular adenoca- trabecular|8332/3
C0334327|T191|SY|BB5f3|RCD|Follicular adenocarcinoma - moderately differentiated|8332/3
C0334327|T191|PT|BB5f3|RCD|Follicular adenocarcinoma - trabecular|8332/3
C0334327|T191|AB|BB5f3|RCD|Follicular ca - trabecular|8332/3
C0334327|T191|SY|BB5f3|RCD|Follicular carcinoma - moderately differentiated|8332/3
C0334327|T191|SY|BB5f3|RCD|Follicular carcinoma - trabecular|8332/3
C0334327|T191|AB|BB5f3|RCD|Follicular carcinoma-mod diff|8332/3
C0302182|T191|PT|BB5F.|RCD|Trabecular adenocarcinoma|8332/3
C0302182|T191|SY|BB5F.|RCD|Trabecular carcinoma|8332/3
C0334327|T191|SY|BB5f3|RCD|Wuchernde Struma Langhans|8332/3
C0334327|T191|SY|72174007|SNOMEDCT_US|Follicular adenocarcinoma - moderately differentiated|8332/3
C0334327|T191|SY|72174007|SNOMEDCT_US|Follicular adenocarcinoma - trabecular|8332/3
C0334327|T191|SY|72174007|SNOMEDCT_US|Follicular adenocarcinoma, moderately differentiated|8332/3
C0334327|T191|PT|72174007|SNOMEDCT_US|Follicular adenocarcinoma, trabecular|8332/3
C0334327|T191|SY|72174007|SNOMEDCT_US|Follicular carcinoma - moderately differentiated|8332/3
C0334327|T191|SY|72174007|SNOMEDCT_US|Follicular carcinoma - trabecular|8332/3
C0334327|T191|SY|72174007|SNOMEDCT_US|Follicular carcinoma, moderately differentiated|8332/3
C0334327|T191|SY|72174007|SNOMEDCT_US|Follicular carcinoma, trabecular|8332/3
C0302182|T191|PT|29792007|SNOMEDCT_US|Trabecular adenocarcinoma|8332/3
C0302182|T191|SY|29792007|SNOMEDCT_US|Trabecular carcinoma|8332/3
C0334327|T191|IS|72174007|SNOMEDCT_US|Wuchernde Struma Langhans|8332/3
C0334328|T191|SY|0000029958|CHV|adenoma fetal|8333/0
C0334328|T191|PT|0000029958|CHV|microfollicular adenoma|8333/0
C0334328|T191|SY|C4160|NCI|Fetal Adenoma|8333/0
C0334328|T191|SY|C4160|NCI|Microfollicular Adenoma|8333/0
C0334328|T191|SY|C4160|NCI|Thyroid Gland Fetal Adenoma|8333/0
C0334328|T191|PT|C4160|NCI|Thyroid Gland Microfollicular Adenoma|8333/0
C0334328|T191|SY|BB5f4|RCD|Fetal adenoma|8333/0
C0334328|T191|PT|BB5f4|RCD|Microfollicular adenoma|8333/0
C0334328|T191|SY|30301008|SNOMEDCT_US|Fetal adenoma|8333/0
C0334328|T191|SY|30301008|SNOMEDCT_US|Foetal adenoma|8333/0
C0334328|T191|PT|30301008|SNOMEDCT_US|Microfollicular adenoma|8333/0
C1266047|T191|PN|NOCODE|MTH|Fetal adenocarcinoma|8333/3
C1708045|T191|PN|NOCODE|MTH|Fetal Lung Adenocarcinoma|8333/3
C1708045|T191|SY|C45509|NCI|Fetal Adenocarcinoma|8333/3
C1708045|T191|SY|TCGA|NCI|Fetal Lung Adenocarcinoma|8333/3
C1708045|T191|PT|C45509|NCI|Lung Fetal Adenocarcinoma|8333/3
C1708045|T191|SY|C45509|NCI|Pulmonary Adenocarcinoma of Fetal Type|8333/3
C1708045|T191|SY|C45509|NCI|Pulmonary Endodermal Tumor Resembling Fetal Lung|8333/3
C1708045|T191|SY|C45509|NCI|Well-Differentiated Fetal Lung Adenocarcinoma|8333/3
C1266047|T191|PT|128893004|SNOMEDCT_US|Fetal adenocarcinoma|8333/3
C1266047|T191|SY|128893004|SNOMEDCT_US|Foetal adenocarcinoma|8333/3
C0334329|T191|PT|MTHU017231|ICPC2ICD10ENG|colloid; adenoma, unspecified site|8334/0
C0334329|T191|SY|C4161|NCI|Colloid Adenoma|8334/0
C0334329|T191|SY|C4161|NCI|Macrofollicular Adenoma|8334/0
C0334329|T191|PT|C4161|NCI|Thyroid Gland Macrofollicular Adenoma|8334/0
C0334329|T191|SY|BB5f5|RCD|Colloid adenoma|8334/0
C0334329|T191|PT|BB5f5|RCD|Macrofollicular adenoma|8334/0
C0334329|T191|SY|26545006|SNOMEDCT_US|Colloid adenoma|8334/0
C0334329|T191|PT|26545006|SNOMEDCT_US|Macrofollicular adenoma|8334/0
C1883338|T191|PT|236230|MEDCIN|minimally invasive follicular carcinoma of the thyroid gland|8335/3
C1883338|T191|SY|236230|MEDCIN|minimally invasive follicular carcinoma of thyroid gland|8335/3
C1883338|T191|SY|C65200|NCI|FTC, Minimally Invasive|8335/3
C1883338|T191|PT|C65200|NCI|Thyroid Gland Follicular Carcinoma, Minimally Invasive|8335/3
C1266048|T191|PT|789444007|SNOMEDCT_US|Encapsulated follicular carcinoma|8335/3
C1266048|T191|IS|128671006|SNOMEDCT_US|Follicular carcinoma, encapsulated|8335/3
C1266048|T191|SY|789444007|SNOMEDCT_US|Follicular carcinoma, encapsulated|8335/3
C1720448|T191|PT|422350000|SNOMEDCT_US|Follicular carcinoma, grossly encapsulated with angioinvasion|8335/3
C1266048|T191|PT|128671006|SNOMEDCT_US|Follicular carcinoma, minimally invasive|8335/3
C1336751|T191|PN|NOCODE|MTH|Thyroid Hyalinizing Trabecular Adenoma|8336/0
C1336751|T191|SY|C6846|NCI|Hyalinizing Trabecular Adenoma of the Thyroid|8336/0
C1336751|T191|SY|C6846|NCI|Hyalinizing Trabecular Adenoma of Thyroid|8336/0
C1336751|T191|SY|C6846|NCI|Hyalinizing Trabecular Tumor|8336/0
C1336751|T191|SY|C6846|NCI|Paraganglioma-like Adenoma|8336/0
C1336751|T191|AB|C6846|NCI|PLAT|8336/0
C1336751|T191|PT|C6846|NCI|Thyroid Gland Hyalinizing Trabecular Tumor|8336/0
C1336751|T191|SY|C6846|NCI|Thyroid Hyalinizing Trabecular Adenoma|8336/0
C1336751|T191|DN|C6846|NCI_CTRP|Thyroid Gland Hyalinizing Trabecular Tumor|8336/0
C1266049|T191|PTGB|128672004|SNOMEDCT_US|Hyalinising trabecular adenoma|8336/0
C1336751|T191|PTGB|722214003|SNOMEDCT_US|Hyalinising trabecular tumour|8336/0
C1266049|T191|PT|128672004|SNOMEDCT_US|Hyalinizing trabecular adenoma|8336/0
C1336751|T191|PT|722214003|SNOMEDCT_US|Hyalinizing trabecular tumor|8336/0
C1266050|T191|PT|0000056680|CHV|insular carcinoma|8337/3
C1266050|T191|PT|10076603|MDR|Poorly differentiated thyroid carcinoma|8337/3
C1266050|T191|LLT|10076603|MDR|Poorly differentiated thyroid carcinoma|8337/3
C1266050|T191|PN|NOCODE|MTH|Poorly Differentiated Thyroid Carcinoma|8337/3
C1266050|T191|SY|C6040|NCI|Insular Carcinoma|8337/3
C1266050|T191|AB|C6040|NCI|PDTC|8337/3
C1266050|T191|SY|C6040|NCI|Poorly Differentiated Carcinoma of the Thyroid Gland|8337/3
C1266050|T191|SY|C6040|NCI|Poorly Differentiated Carcinoma of Thyroid Gland|8337/3
C1266050|T191|SY|C6040|NCI|Poorly Differentiated Thyroid Carcinoma|8337/3
C1266050|T191|PT|C6040|NCI|Poorly Differentiated Thyroid Gland Carcinoma|8337/3
C1266050|T191|SY|C6040|NCI|Thyroid Gland Poorly Differentiated Carcinoma|8337/3
C1266050|T191|DN|C6040|NCI_CTRP|Poorly Differentiated Thyroid Gland Cancer|8337/3
C1266050|T191|SY|CDR0000038462|PDQ|insular carcinoma|8337/3
C1266050|T191|PT|CDR0000038462|PDQ|insular thyroid cancer|8337/3
C1266050|T191|SY|CDR0000038462|PDQ|poorly differentiated carcinoma of the thyroid gland|8337/3
C1266050|T191|SY|CDR0000038462|PDQ|poorly differentiated carcinoma of thyroid gland|8337/3
C1266050|T191|SY|CDR0000038462|PDQ|poorly differentiated thyroid carcinoma|8337/3
C1266050|T191|SY|CDR0000038462|PDQ|poorly differentiated thyroid gland carcinoma|8337/3
C1266050|T191|SY|CDR0000038462|PDQ|thyroid gland poorly differentiated carcinoma|8337/3
C1266050|T191|PT|128673009|SNOMEDCT_US|Insular carcinoma|8337/3
C0206683|T191|PT|MTHU003384|ICPC2ICD10ENG|adenocarcinoma; follicular with papillary|8340/3
C0206683|T191|PT|MTHU003413|ICPC2ICD10ENG|adenocarcinoma; papillary with follicular|8340/3
C0206683|T191|PT|MTHU003414|ICPC2ICD10ENG|adenocarcinoma; papillary, follicular variant|8340/3
C0206683|T191|PT|MTHU014752|ICPC2ICD10ENG|carcinoma; follicular with papillary|8340/3
C0206683|T191|PT|MTHU014807|ICPC2ICD10ENG|carcinoma; papillary with follicular|8340/3
C0206683|T191|PT|MTHU014808|ICPC2ICD10ENG|carcinoma; papillary, follicular variant|8340/3
C0206683|T191|PT|MTHU029185|ICPC2ICD10ENG|follicular; adenocarcinoma with papillary|8340/3
C0206683|T191|PT|MTHU029193|ICPC2ICD10ENG|follicular; carcinoma, with papillary|8340/3
C0206683|T191|PT|MTHU057275|ICPC2ICD10ENG|papillary; adenocarcinoma with follicular|8340/3
C0206683|T191|PT|MTHU057276|ICPC2ICD10ENG|papillary; adenocarcinoma, follicular variant|8340/3
C0206683|T191|PT|MTHU057282|ICPC2ICD10ENG|papillary; carcinoma, follicular variant|8340/3
C0206683|T191|PT|MTHU057286|ICPC2ICD10ENG|papillary; carcinoma, with follicular|8340/3
C0206683|T191|MH|D018265|MSH|Carcinoma, Papillary, Follicular|8340/3
C0206683|T191|PN|NOCODE|MTH|Papillary and follicular adenocarcinoma|8340/3
C4745261|T191|PT|C7381|NCI|Follicular Variant Thyroid Gland Papillary Carcinoma, Infiltrative Subtype|8340/3
C0206683|T191|OP|C7380|NCI|Papillary and Follicular Adenocarcinoma|8340/3
C0206683|T191|OP|C7380|NCI|Papillary and Follicular Carcinoma|8340/3
C0206683|T191|OP|C7380|NCI|Thyroid Gland Papillary and Follicular Carcinoma|8340/3
C0206683|T191|PT|C7380|NCI|Thyroid Gland Papillary and Follicular Carcinoma|8340/3
C0206683|T191|AB|Xa98Q|RCD|Papill adenoca-follic variant|8340/3
C0206683|T191|OA|BB5f6|RCD|Papillary + follicular adenoca|8340/3
C0206683|T191|SY|Xa98Q|RCD|Papillary adenocarcinoma - follicular variant|8340/3
C0206683|T191|OP|BB5f6|RCD|Papillary and follicular adenocarcinoma|8340/3
C0206683|T191|AB|Xa98Q|RCD|Papillary and follicular ca|8340/3
C0206683|T191|SY|Xa98Q|RCD|Papillary and follicular carcinoma|8340/3
C0206683|T191|AB|Xa98Q|RCD|Papillary ca - follic variant|8340/3
C0206683|T191|PT|Xa98Q|RCD|Papillary carcinoma - follicular variant|8340/3
C0206683|T191|SY|21968007|SNOMEDCT_US|Papillary adenocarcinoma - follicular variant|8340/3
C0206683|T191|SY|21968007|SNOMEDCT_US|Papillary adenocarcinoma, follicular variant|8340/3
C0206683|T191|PT|189643000|SNOMEDCT_US|Papillary and follicular adenocarcinoma|8340/3
C0206683|T191|SY|21968007|SNOMEDCT_US|Papillary and follicular adenocarcinoma|8340/3
C0206683|T191|SY|21968007|SNOMEDCT_US|Papillary and follicular carcinoma|8340/3
C0206683|T191|SY|21968007|SNOMEDCT_US|Papillary carcinoma - follicular variant|8340/3
C1719806|T191|PT|421918000|SNOMEDCT_US|Papillary carcinoma, diffuse follicular|8340/3
C0206683|T191|PT|21968007|SNOMEDCT_US|Papillary carcinoma, follicular variant|8340/3
C1709457|T191|PT|236254|MEDCIN|papillary microcarcinoma of the thyroid gland|8341/3
C1709457|T191|SY|236254|MEDCIN|papillary microcarcinoma of thyroid gland|8341/3
C1709457|T191|NM|C563277|MSH|Papillary Thyroid Microcarcinoma|8341/3
C1709457|T191|SY|C46004|NCI|Papillary Microcarcinoma of the Thyroid|8341/3
C1709457|T191|SY|C46004|NCI|Papillary Microcarcinoma of the Thyroid Gland|8341/3
C1709457|T191|SY|C46004|NCI|Papillary Thyroid Gland Microcarcinoma|8341/3
C1709457|T191|SY|C46004|NCI|Papillary Thyroid Microcarcinoma|8341/3
C1709457|T191|PT|C46004|NCI|Thyroid Gland Papillary Microcarcinoma|8341/3
C1266051|T191|PT|128674003|SNOMEDCT_US|Papillary microcarcinoma|8341/3
C1709312|T191|PT|C46093|NCI|Oncocytic Variant Thyroid Gland Papillary Carcinoma|8342/3
C1709312|T191|SY|TCGA|NCI|Oncocytic Variant Thyroid Gland Papillary Carcinoma|8342/3
C1709312|T191|SY|C46093|NCI|Oxyphilic Variant Thyroid Gland Papillary Carcinoma|8342/3
C1709312|T191|DN|C46093|NCI_CTRP|Oncocytic Variant Thyroid Gland Papillary Cancer|8342/3
C1266052|T191|PT|128675002|SNOMEDCT_US|Papillary carcinoma, oxyphilic cell|8342/3
C1266053|T191|PN|NOCODE|MTH|Encapsulated papillary carcinoma|8343/3
C4745260|T191|PT|C66850|NCI|Follicular Variant Thyroid Gland Papillary Carcinoma, Encapsulated Subtype with Invasion|8343/3
C1266053|T191|PT|703545003|SNOMEDCT_US|Encapsulated papillary carcinoma|8343/3
C1266053|T191|SY|703545003|SNOMEDCT_US|Encysted papillary carcinoma|8343/3
C1266053|T191|SY|703545003|SNOMEDCT_US|Intracystic papillary adenocarcinoma|8343/3
C1266053|T191|SY|703545003|SNOMEDCT_US|Intracystic papillary carcinoma|8343/3
C1266053|T191|SY|703545003|SNOMEDCT_US|Non-infiltrating intracystic carcinoma|8343/3
C1266053|T191|SY|703545003|SNOMEDCT_US|Noninfiltrating intracystic carcinoma|8343/3
C1266053|T191|OAP|128676001|SNOMEDCT_US|Papillary carcinoma, encapsulated|8343/3
C1266054|T191|PN|NOCODE|MTH|Papillary carcinoma, columnar cell|8344/3
C2939464|T191|PN|NOCODE|MTH|Papillary carcinoma, tall cell|8344/3
C1333120|T191|SY|C35830|NCI|Columnar Cell Variant Papillary Carcinoma|8344/3
C1333120|T191|SY|C35830|NCI|Columnar Cell Variant Papillary Thyroid Gland Carcinoma|8344/3
C1333120|T191|PT|C35830|NCI|Columnar Cell Variant Thyroid Gland Papillary Carcinoma|8344/3
C1266054|T191|PT|128677005|SNOMEDCT_US|Papillary carcinoma, columnar cell|8344/3
C1266054|T191|SY|128677005|SNOMEDCT_US|Papillary carcinoma, tall cell|8344/3
C2939464|T191|PT|422198004|SNOMEDCT_US|Papillary carcinoma, tall cell|8344/3
C0334379|T191|PT|MTHU014793|ICPC2ICD10ENG|carcinoma; medullary with amyloid stroma, unspecified site|8345/3
C0334379|T191|PT|MTHU048008|ICPC2ICD10ENG|medullary; carcinoma with amyloid stroma, unspecified site|8345/3
C0334379|T191|SY|236232|MEDCIN|medullary carcinoma of thyroid gland with amyloid stroma|8345/3
C0334379|T191|SY|236232|MEDCIN|medullary carcinoma of thyroid with amyloid stroma|8345/3
C0334379|T191|PT|236232|MEDCIN|medullary thyroid carcinoma with amyloid stroma|8345/3
C0334379|T191|PN|NOCODE|MTH|Thyroid Gland Medullary Carcinoma with Amyloid Stroma|8345/3
C0334379|T191|SY|C4193|NCI|C Cell Adenocarcinoma with Amyloid Stroma|8345/3
C0334379|T191|SY|C4193|NCI|C Cell Carcinoma with Amyloid Stroma|8345/3
C0334379|T191|SY|C4193|NCI|Medullary Adenocarcinoma with Amyloid Stroma|8345/3
C0334379|T191|SY|C4193|NCI|Medullary Carcinoma with Amyloid Stroma|8345/3
C0334379|T191|SY|C4193|NCI|Medullary Thyroid Gland Carcinoma with Amyloid Stroma|8345/3
C0334379|T191|SY|C4193|NCI|Parafollicular Cell Adenocarcinoma with Amyloid Stroma|8345/3
C0334379|T191|SY|C4193|NCI|Parafollicular Cell Carcinoma with Amyloid Stroma|8345/3
C0334379|T191|PT|C4193|NCI|Thyroid Gland Medullary Carcinoma with Amyloid Stroma|8345/3
C0334379|T191|AB|BB9C.|RCD|Medullary ca + amyloid stroma|8345/3
C0334379|T191|PT|BB9C.|RCD|Medullary carcinoma with amyloid stroma|8345/3
C0334379|T191|OAP|36538001|SNOMEDCT_US|Medullary carcinoma with amyloid stroma|8345/3
C0334379|T191|PT|128916007|SNOMEDCT_US|Medullary carcinoma with amyloid stroma|8345/3
C0334379|T191|IS|36538001|SNOMEDCT_US|Medullary carcinoma with amyloid stroma -RETIRED-|8345/3
C0334379|T191|OF|36538001|SNOMEDCT_US|Medullary carcinoma with amyloid stroma -RETIRED-|8345/3
C1710414|T191|SY|236234|MEDCIN|mixed medullary-papillary carcinoma of thyroid gland|8346/3
C1710414|T191|PT|236234|MEDCIN|mixed medullary-papillary thyroid carcinoma|8346/3
C1710414|T191|PN|NOCODE|MTH|Thyroid Gland Mixed Medullary and Papillary Carcinoma|8346/3
C1710414|T191|AB|C46104|NCI|MMFTC|8346/3
C1710414|T191|PT|C46104|NCI|Thyroid Gland Mixed Medullary and Follicular Cell Carcinoma|8346/3
C1710414|T191|SY|C46104|NCI|Thyroid Gland Mixed Medullary and Papillary Carcinoma|8346/3
C1266055|T191|PT|128678000|SNOMEDCT_US|Mixed medullary-follicular carcinoma|8346/3
C1710414|T191|SY|236234|MEDCIN|mixed medullary-papillary carcinoma of thyroid gland|8347/3
C1710414|T191|PT|236234|MEDCIN|mixed medullary-papillary thyroid carcinoma|8347/3
C1710414|T191|PN|NOCODE|MTH|Thyroid Gland Mixed Medullary and Papillary Carcinoma|8347/3
C1710414|T191|AB|C46104|NCI|MMFTC|8347/3
C1710414|T191|PT|C46104|NCI|Thyroid Gland Mixed Medullary and Follicular Cell Carcinoma|8347/3
C1710414|T191|SY|C46104|NCI|Thyroid Gland Mixed Medullary and Papillary Carcinoma|8347/3
C1266056|T191|PT|128679008|SNOMEDCT_US|Mixed medullary-papillary carcinoma|8347/3
C0334330|T191|PT|MTHU003412|ICPC2ICD10ENG|adenocarcinoma; nonencapsulated sclerosing|8350/3
C0334330|T191|PT|MTHU014797|ICPC2ICD10ENG|carcinoma; nonencapsulated sclerosing|8350/3
C0334330|T191|PT|MTHU053295|ICPC2ICD10ENG|nonencapsulated sclerosing; carcinoma|8350/3
C0334330|T191|PT|MTHU053241|ICPC2ICD10ENG|nonencapsulated; sclerosing adenocarcinoma|8350/3
C0334330|T191|PT|MTHU053242|ICPC2ICD10ENG|nonencapsulated; sclerosing tumor|8350/3
C0334330|T191|PT|MTHU077107|ICPC2ICD10ENG|tumor; nonencapsulated sclerosing|8350/3
C0334330|T191|PT|C7427|NCI|Diffuse Sclerosing Variant Thyroid Gland Papillary Carcinoma|8350/3
C0334330|T191|SY|C7427|NCI|Nonencapsulated Sclerosing Adenocarcinoma|8350/3
C0334330|T191|SY|C7427|NCI|Nonencapsulated Sclerosing Carcinoma|8350/3
C0334330|T191|SY|C7427|NCI|Nonencapsulated Sclerosing Neoplasm|8350/3
C0334330|T191|SY|C7427|NCI|Nonencapsulated Sclerosing Papillary Thyroid Carcinoma|8350/3
C0334330|T191|SY|C7427|NCI|Nonencapsulated Sclerosing Tumor|8350/3
C0334330|T191|SY|C7427|NCI|Thyroid Gland Diffuse Sclerosing Papillary Carcinoma|8350/3
C0334330|T191|AB|BB5f7|RCD|Nonencapsul sclerosing adenoca|8350/3
C0334330|T191|AB|BB5f7|RCD|Nonencapsul sclerosing tumour|8350/3
C0334330|T191|SY|BB5f7|RCD|Nonencapsulated sclerosing adenocarcinoma|8350/3
C0334330|T191|AB|BB5f7|RCD|Nonencapsulated sclerosing ca|8350/3
C0334330|T191|PT|BB5f7|RCD|Nonencapsulated sclerosing carcinoma|8350/3
C0334330|T191|SY|BB5f7|RCD|Nonencapsulated sclerosing tumour|8350/3
C0334330|T191|AB|BB5f7|RCDAE|Nonencapsul sclerosing tumor|8350/3
C0334330|T191|SY|BB5f7|RCDAE|Nonencapsulated sclerosing tumor|8350/3
C0334330|T191|SY|62681000|SNOMEDCT_US|Nonencapsulated sclerosing adenocarcinoma|8350/3
C0334330|T191|PT|62681000|SNOMEDCT_US|Nonencapsulated sclerosing carcinoma|8350/3
C0334330|T191|SY|62681000|SNOMEDCT_US|Nonencapsulated sclerosing tumor|8350/3
C0334330|T191|SYGB|62681000|SNOMEDCT_US|Nonencapsulated sclerosing tumour|8350/3
C0334330|T191|SY|62681000|SNOMEDCT_US|Papillary carcinoma, diffuse sclerosing|8350/3
C0027662|T191|ET|0000004642|AOD|multiple endocrine neoplasm|8360/1
C0027662|T191|SY|0000008568|CHV|endocrine multiple neoplasia|8360/1
C0027662|T191|SY|0000008568|CHV|mea|8360/1
C0027662|T191|SY|0000008568|CHV|meas|8360/1
C0027662|T191|SY|0000008568|CHV|multiple endocrine adenoma|8360/1
C0027662|T191|SY|0000008568|CHV|multiple endocrine adenomatosis|8360/1
C0027662|T191|PT|0000008568|CHV|multiple endocrine neoplasia|8360/1
C0027662|T191|SY|0000008568|CHV|multiple endocrine neoplasias|8360/1
C0027662|T191|SY|0000008568|CHV|multiple endocrine neoplasm|8360/1
C0027662|T191|SY|0000008568|CHV|multiple endocrine neoplasms|8360/1
C0027662|T191|SY|0000008568|CHV|multiple endocrine tumasia|8360/1
C0027662|T191|ET|2009-6300|CSP|MEA|8360/1
C0027662|T191|ET|2009-6300|CSP|multiple endocrine adenopathy|8360/1
C0027662|T191|PT|2009-6300|CSP|multiple endocrine neoplasia|8360/1
C0027662|T191|SY|NOCODE|DXP|MEA SYNDROME|8360/1
C0027662|T191|ET|E31.2|ICD10CM|Multiple endocrine adenomatosis|8360/1
C0027662|T191|ET|E31.20|ICD10CM|Multiple endocrine adenomatosis NOS|8360/1
C0027662|T191|PT|sh85000844|LCH_NW|Adenomatosis, Familial endocrine|8360/1
C0027662|T191|LLT|10061299|MDR|Multiple endocrine adenomatosis|8360/1
C0027662|T191|LLT|10028189|MDR|Multiple endocrine adenomatosis NOS|8360/1
C0027662|T191|LLT|10051747|MDR|Multiple endocrine neoplasia|8360/1
C0027662|T191|PT|10051747|MDR|Multiple endocrine neoplasia|8360/1
C0027662|T191|HT|10028193|MDR|Multiple endocrine neoplasia syndromes|8360/1
C0027662|T191|HT|10028196|MDR|Multiple endocrine neoplasias|8360/1
C0027662|T191|PT|30455|MEDCIN|multiple endocrine neoplasia|8360/1
C0027662|T191|ET|475|MEDLINEPLUS|Multiple Endocrine Neoplasia|8360/1
C0027662|T191|ET|356|MEDLINEPLUS|Multiple Endocrine Neoplasia|8360/1
C0027662|T191|PM|D009377|MSH|Adenomatoses, Familial Endocrine|8360/1
C0027662|T191|PM|D009377|MSH|Adenomatoses, Multiple Endocrine|8360/1
C0027662|T191|ET|D009377|MSH|Adenomatosis, Familial Endocrine|8360/1
C0027662|T191|ET|D009377|MSH|Adenomatosis, Multiple Endocrine|8360/1
C0027662|T191|PM|D009377|MSH|Adenopathies, Multiple Endocrine|8360/1
C0027662|T191|PM|D009377|MSH|Adenopathy, Multiple Endocrine|8360/1
C0027662|T191|PM|D009377|MSH|Endocrine Adenomatoses, Familial|8360/1
C0027662|T191|PM|D009377|MSH|Endocrine Adenomatoses, Multiple|8360/1
C0027662|T191|PM|D009377|MSH|Endocrine Adenomatosis, Familial|8360/1
C0027662|T191|PM|D009377|MSH|Endocrine Adenomatosis, Multiple|8360/1
C0027662|T191|PM|D009377|MSH|Endocrine Adenopathies, Multiple|8360/1
C0027662|T191|PM|D009377|MSH|Endocrine Adenopathy, Multiple|8360/1
C0027662|T191|DEV|D009377|MSH|ENDOCRINE NEOPL MULTIPLE|8360/1
C0027662|T191|ET|D009377|MSH|Endocrine Neoplasia, Multiple|8360/1
C0027662|T191|PM|D009377|MSH|Endocrine Neoplasms, Multiple|8360/1
C0027662|T191|PM|D009377|MSH|Familial Endocrine Adenomatoses|8360/1
C0027662|T191|ET|D009377|MSH|Familial Endocrine Adenomatosis|8360/1
C0027662|T191|PM|D009377|MSH|Multiple Endocrine Adenomatoses|8360/1
C0027662|T191|ET|D009377|MSH|Multiple Endocrine Adenomatosis|8360/1
C0027662|T191|PM|D009377|MSH|Multiple Endocrine Adenopathies|8360/1
C0027662|T191|ET|D009377|MSH|Multiple Endocrine Adenopathy|8360/1
C0027662|T191|DEV|D009377|MSH|MULTIPLE ENDOCRINE NEOPL|8360/1
C0027662|T191|DEV|D009377|MSH|MULTIPLE ENDOCRINE NEOPL SYNDROMES|8360/1
C0027662|T191|MH|D009377|MSH|Multiple Endocrine Neoplasia|8360/1
C0027662|T191|ET|D009377|MSH|Multiple Endocrine Neoplasia Syndromes|8360/1
C0027662|T191|ET|D009377|MSH|Multiple Endocrine Neoplasms|8360/1
C0027662|T191|DEV|D009377|MSH|NEOPL MULTIPLE ENDOCRINE|8360/1
C0027662|T191|ET|D009377|MSH|Neoplasia, Multiple Endocrine|8360/1
C0027662|T191|ET|D009377|MSH|Neoplasms, Multiple Endocrine|8360/1
C0027662|T191|PN|NOCODE|MTH|Multiple Endocrine Neoplasia|8360/1
C0027662|T191|ET|258.0|MTHICD9|MEN syndromes|8360/1
C0027662|T191|ET|258.0|MTHICD9|Multiple endocrine neoplasia syndromes|8360/1
C0027662|T191|AB|C6432|NCI|MEN|8360/1
C0027662|T191|SY|C6432|NCI|Multiple Endocrine Adenomatosis|8360/1
C0027662|T191|PT|C6432|NCI|Multiple Endocrine Neoplasia|8360/1
C0027662|T191|SY|C6432|NCI|Multiple Endocrine Neoplasia Syndrome|8360/1
C0027662|T191|DN|C6432|NCI_CTRP|Multiple Endocrine Neoplasia|8360/1
C0027662|T191|PT|CDR0000563964|NCI_NCI-GLOSS|MEN syndrome|8360/1
C0027662|T191|PT|CDR0000270863|NCI_NCI-GLOSS|multiple endocrine adenomatosis|8360/1
C0027662|T191|PT|CDR0000044551|NCI_NCI-GLOSS|multiple endocrine neoplasia syndrome|8360/1
C0027662|T191|SY|C6432|NCI_NICHD|MEN Syndromes|8360/1
C0027662|T191|AB|CDR0000042848|PDQ|MEN|8360/1
C0027662|T191|SY|CDR0000042848|PDQ|Multiple Endocrine Adenomatosis|8360/1
C0027662|T191|SY|CDR0000042848|PDQ|Multiple Endocrine Adenomatosis NOS|8360/1
C0027662|T191|PT|CDR0000042848|PDQ|multiple endocrine neoplasia|8360/1
C0027662|T191|SY|CDR0000042848|PDQ|Multiple Endocrine Neoplasia Syndrome|8360/1
C0027662|T191|SY|XE10q|RCD|Endocrine adenomatosis|8360/1
C0027662|T191|AB|XE10q|RCD|MEA - Multip endocr adenomatos|8360/1
C0027662|T191|SY|XE10q|RCD|MEA - Multiple endocrine adenomatosis|8360/1
C0027662|T191|SY|XE10q|RCD|MEN - Multiple endocrine neoplasia|8360/1
C0027662|T191|AB|XE10q|RCD|MEN-Multiple endocrine neoplas|8360/1
C0027662|T191|OP|BB5g.|RCD|Multiple endocrine adenomas|8360/1
C0027662|T191|SY|XE10q|RCD|Multiple endocrine adenomatosis|8360/1
C0027662|T191|PT|XE10q|RCD|Multiple endocrine neoplasia|8360/1
C0027662|T191|SY|XE10q|RCD|Multiple endocrine tumasia|8360/1
C0027662|T191|AB|XE10q|RCD|Multple endocrine adenomatosis|8360/1
C0027662|T191|SY|60549007|SNOMEDCT_US|Endocrine adenomatosis|8360/1
C0027662|T191|SY|46724008|SNOMEDCT_US|Familial polyendocrine adenomatosis|8360/1
C0027662|T191|SY|46724008|SNOMEDCT_US|MEA - Multiple endocrine adenomatosis|8360/1
C0027662|T191|SY|46724008|SNOMEDCT_US|MEN - Multiple endocrine neoplasia|8360/1
C0027662|T191|PT|60549007|SNOMEDCT_US|Multiple endocrine adenomas|8360/1
C0027662|T191|OAS|190566000|SNOMEDCT_US|Multiple endocrine adenomatosis|8360/1
C0027662|T191|SY|46724008|SNOMEDCT_US|Multiple endocrine neoplasia|8360/1
C0027662|T191|SY|46724008|SNOMEDCT_US|Multiple endocrine tumasia|8360/1
C0334331|T191|PT|MTHU040709|ICPC2ICD10ENG|juxtaglomerular; tumor|8361/0
C0334331|T191|PT|MTHU064212|ICPC2ICD10ENG|reninoma|8361/0
C0334331|T191|PT|MTHU077076|ICPC2ICD10ENG|tumor; juxtaglomerular|8361/0
C0334331|T191|PT|31530|MEDCIN|juxtaglomerular cell tumor of kidney|8361/0
C0334331|T191|SY|31530|MEDCIN|juxtoglomerular cell tumor|8361/0
C0334331|T191|PT|C4162|NCI|Juxtaglomerular Cell Tumor|8361/0
C0334331|T191|SY|C4162|NCI|Juxtaglomerular Neoplasm|8361/0
C0334331|T191|SY|C4162|NCI|Juxtaglomerular Tumor|8361/0
C0334331|T191|SY|C4162|NCI|Reninoma|8361/0
C0334331|T191|PT|XaBBG|RCD|Juxtaglomerular tumour|8361/0
C0334331|T191|SY|XaBBG|RCD|Reninoma|8361/0
C0334331|T191|PT|XaBBG|RCDAE|Juxtaglomerular tumor|8361/0
C0334331|T191|PT|BB5a1|RCDSA|Juxtaglomerular tumor|8361/0
C0334331|T191|PT|BB5a1|RCDSY|Juxtaglomerular tumour|8361/0
C0334331|T191|OAP|5175004|SNOMEDCT_US|Juxtaglomerular tumor|8361/0
C0334331|T191|PT|307618001|SNOMEDCT_US|Juxtaglomerular tumor|8361/0
C0334331|T191|PT|128860008|SNOMEDCT_US|Juxtaglomerular tumor|8361/0
C0334331|T191|IS|5175004|SNOMEDCT_US|Juxtaglomerular tumor -RETIRED-|8361/0
C0334331|T191|OF|5175004|SNOMEDCT_US|Juxtaglomerular tumor -RETIRED-|8361/0
C0334331|T191|OAP|5175004|SNOMEDCT_US|Juxtaglomerular tumour|8361/0
C0334331|T191|PTGB|307618001|SNOMEDCT_US|Juxtaglomerular tumour|8361/0
C0334331|T191|PTGB|128860008|SNOMEDCT_US|Juxtaglomerular tumour|8361/0
C0334331|T191|IS|5175004|SNOMEDCT_US|Juxtaglomerular tumour -RETIRED-|8361/0
C0334331|T191|SY|128860008|SNOMEDCT_US|Reninoma|8361/0
C0334331|T191|IS|5175004|SNOMEDCT_US|Reninoma|8361/0
C0334331|T191|SY|307618001|SNOMEDCT_US|Reninoma|8361/0
C0206667|T191|PT|0013562|CCPSS|ADRENAL ADENOMA|8370/0
C0206667|T191|SY|0000025374|CHV|adenoma adrenal|8370/0
C0206667|T191|SY|0000021007|CHV|adenoma adrenal cortex|8370/0
C0206667|T191|SY|0000021007|CHV|adenoma adrenal cortical|8370/0
C0206667|T191|SY|0000025374|CHV|adenomas adrenal|8370/0
C0206667|T191|PT|0000025374|CHV|adrenal adenoma|8370/0
C0206667|T191|PT|0000021007|CHV|adrenal cortical adenoma|8370/0
C0206667|T191|SY|0000021007|CHV|adrenocortical adenoma|8370/0
C0206667|T191|PT|U000083|COSTAR|ADRENAL ADENOMA|8370/0
C0206667|T191|PT|U000123|COSTAR|BENIGN ADRENAL ADENOMA|8370/0
C0206667|T191|GT|ADENOMA|CST|ADENOMA ADRENAL|8370/0
C0206667|T191|DI|U000044|DXP|ADRENAL CORTEX, ADENOMA|8370/0
C0206667|T191|PT|HP:0008256|HPO|Adrenocortical adenoma|8370/0
C0206667|T191|SY|HP:0008256|HPO|Adrenocortical adenomas|8370/0
C0206667|T191|PT|MTHU003479|ICPC2ICD10ENG|adenoma; adrenal|8370/0
C0206667|T191|PT|MTHU010756|ICPC2ICD10ENG|adrenal; adenoma|8370/0
C0206667|T191|PT|T73011|ICPC2P|Adenoma;adrenal|8370/0
C0206667|T191|PTN|T73011|ICPC2P|adrenal adenoma|8370/0
C0206667|T191|LLT|10001232|MDR|Adenoma adrenal|8370/0
C0206667|T191|LLT|10001323|MDR|Adrenal adenoma|8370/0
C0206667|T191|PT|10001323|MDR|Adrenal adenoma|8370/0
C0206667|T191|PT|91180|MEDCIN|adrenal cortical adenoma|8370/0
C0206667|T191|ET|D018246|MSH|Adenoma, Adrenal Cortical|8370/0
C0206667|T191|ET|D018246|MSH|Adenoma, Adrenocortical|8370/0
C0206667|T191|PM|D018246|MSH|Adenomas, Adrenal Cortical|8370/0
C0206667|T191|PM|D018246|MSH|Adenomas, Adrenocortical|8370/0
C0206667|T191|PM|D018246|MSH|Adrenal Cortical Adenoma|8370/0
C0206667|T191|PM|D018246|MSH|Adrenal Cortical Adenomas|8370/0
C0206667|T191|MH|D018246|MSH|Adrenocortical Adenoma|8370/0
C0206667|T191|PM|D018246|MSH|Adrenocortical Adenomas|8370/0
C0206667|T191|PN|NOCODE|MTH|Adrenal Cortical Adenoma|8370/0
C0206667|T191|SY|C9003|NCI|Adenoma of Adrenal Cortex|8370/0
C0206667|T191|SY|C9003|NCI|Adenoma of Adrenal Gland|8370/0
C0206667|T191|SY|C9003|NCI|Adenoma of the Adrenal Cortex|8370/0
C0206667|T191|SY|C9003|NCI|Adenoma of the Adrenal Gland|8370/0
C0206667|T191|SY|C9003|NCI|Adrenal Adenoma|8370/0
C0206667|T191|PT|C9003|NCI|Adrenal Cortex Adenoma|8370/0
C0206667|T191|SY|C9003|NCI|Adrenal Cortical Adenoma|8370/0
C0206667|T191|SY|C9003|NCI|Adrenal Gland Adenoma|8370/0
C0206667|T191|SY|C9003|NCI|Adrenocortical Adenoma|8370/0
C0206667|T191|SY|C9003|NCI|Benign Adenoma of Adrenal Gland|8370/0
C0206667|T191|SY|C9003|NCI|Benign Adenoma of the Adrenal Gland|8370/0
C0206667|T191|SY|C9003|NCI|Benign Adrenal Adenoma|8370/0
C0206667|T191|SY|C9003|NCI|Benign Adrenal Gland Adenoma|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Adenoma of Adrenal Cortex|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Adenoma of Adrenal Gland|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Adenoma of the Adrenal Cortex|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Adenoma of the Adrenal Gland|8370/0
C0206667|T191|PT|C9003|NCI_CDISC|ADENOMA, ADRENOCORTICAL, BENIGN|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Adrenal Adenoma|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Adrenal Cortical Adenoma|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Adrenal Gland Adenoma|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Adrenocortical Adenoma|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Benign Adenoma of Adrenal Gland|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Benign Adenoma of the Adrenal Gland|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Benign Adrenal Adenoma|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Benign Adrenal Gland Adenoma|8370/0
C0206667|T191|SY|C9003|NCI_CDISC|Cortical Cell Adenoma|8370/0
C0206667|T191|PT|X78ce|RCD|Adrenal adenoma|8370/0
C0206667|T191|PT|Xa98S|RCD|Adrenal cortical adenoma|8370/0
C0206667|T191|PT|XaBBL|RCD|Adrenal cortical adenoma - morphology|8370/0
C0206667|T191|AB|XaBBL|RCD|Adrenal cortical adenoma-morph|8370/0
C0206667|T191|OA|BB5h0|RCDSY|Adrenal cortic. adenoma NOS|8370/0
C0206667|T191|OP|BB5h0|RCDSY|Adrenal cortical adenoma NOS|8370/0
C0206667|T191|PT|255036008|SNOMEDCT_US|Adrenal adenoma|8370/0
C0206667|T191|IS|18365006|SNOMEDCT_US|Adrenal cortical adenoma|8370/0
C0206667|T191|PT|302826002|SNOMEDCT_US|Adrenal cortical adenoma|8370/0
C1444008|T191|PT|409703003|SNOMEDCT_US|Adrenal cortical adenoma - category|8370/0
C0206667|T191|OAP|134348000|SNOMEDCT_US|Adrenal cortical adenoma - morphology|8370/0
C0206667|T191|OF|134348000|SNOMEDCT_US|Adrenal cortical adenoma - morphology|8370/0
C0206667|T191|PT|18365006|SNOMEDCT_US|Adrenal cortical adenoma morphology|8370/0
C0206667|T191|SY|18365006|SNOMEDCT_US|Adrenal cortical adenoma, no ICD-O subtype|8370/0
C0206667|T191|SY|18365006|SNOMEDCT_US|Adrenal cortical adenoma, no International Classification of Diseases for Oncology subtype|8370/0
C0206667|T191|IS|18365006|SNOMEDCT_US|Adrenal cortical adenoma, NOS|8370/0
C0206667|T191|PT|1810|WHO|ADENOMA ADRENAL|8370/0
C0206686|T191|SY|0000021020|CHV|adenocarcinoma adrenal|8370/3
C0206686|T191|SY|0000021020|CHV|adrenal adenocarcinoma|8370/3
C0206686|T191|PT|0000021020|CHV|adrenal carcinoma|8370/3
C0206686|T191|SY|0000021020|CHV|adrenal carcinomas|8370/3
C0206686|T191|SY|0000021020|CHV|adrenal cortex carcinoma|8370/3
C0206686|T191|SY|0000021020|CHV|adrenal cortical carcinoma|8370/3
C0206686|T191|SY|0000021020|CHV|adrenocortical carcinoma|8370/3
C0206686|T191|SY|0000021020|CHV|carcinoma adrenal|8370/3
C0206686|T191|PT|U000084|COSTAR|ADRENAL CARCINOMA|8370/3
C0206686|T191|GT|CARCINOMA|CST|CARCINOMA ADRENAL|8370/3
C0206686|T191|SY|NOCODE|DXP|ADRENAL CORTEX CANCER, CARCINOMA|8370/3
C0206686|T191|DI|U000045|DXP|ADRENAL CORTEX, CARCINOMA|8370/3
C0206686|T191|SY|HP:0006744|HPO|Adrenal carcinoma|8370/3
C0206686|T191|SY|HP:0006744|HPO|Adrenal gland carinoma|8370/3
C0206686|T191|PT|HP:0006744|HPO|Adrenocortical carcinoma|8370/3
C0206686|T191|PT|MTHU003373|ICPC2ICD10ENG|adenocarcinoma; adrenal cortical|8370/3
C0206686|T191|PT|MTHU010827|ICPC2ICD10ENG|adrenal cortical; adenocarcinoma|8370/3
C0206686|T191|PT|MTHU010828|ICPC2ICD10ENG|adrenal cortical; carcinoma|8370/3
C0206686|T191|PT|MTHU014731|ICPC2ICD10ENG|carcinoma; adrenal cortical|8370/3
C0206686|T191|LLT|10055076|MDR|Adrenal adenocarcinoma|8370/3
C0206686|T191|LLT|10001326|MDR|Adrenal carcinoma|8370/3
C0206686|T191|LLT|10001327|MDR|Adrenal carcinoma NOS|8370/3
C0206686|T191|PT|10001388|MDR|Adrenocortical carcinoma|8370/3
C0206686|T191|LLT|10001388|MDR|Adrenocortical carcinoma|8370/3
C0206686|T191|LLT|10007285|MDR|Carcinoma adrenal|8370/3
C0206686|T191|PT|236329|MEDCIN|adenocarcinoma of adrenal gland|8370/3
C0206686|T191|SY|236329|MEDCIN|adrenal adenocarcinoma|8370/3
C0206686|T191|SY|236318|MEDCIN|adrenal carcinoma|8370/3
C0206686|T191|SY|30561|MEDCIN|adrenocortical carcinoma|8370/3
C0206686|T191|PT|30561|MEDCIN|adrenocortical carcinoma of adrenal gland|8370/3
C0206686|T191|PT|236318|MEDCIN|carcinoma of adrenal gland|8370/3
C0206686|T191|PM|D018268|MSH|Adrenal Cortical Carcinoma|8370/3
C0206686|T191|PM|D018268|MSH|Adrenal Cortical Carcinomas|8370/3
C0206686|T191|MH|D018268|MSH|Adrenocortical Carcinoma|8370/3
C0206686|T191|PM|D018268|MSH|Adrenocortical Carcinomas|8370/3
C0206686|T191|ET|D018268|MSH|Carcinoma, Adrenal Cortical|8370/3
C0206686|T191|ET|D018268|MSH|Carcinoma, Adrenocortical|8370/3
C0206686|T191|PM|D018268|MSH|Carcinomas, Adrenal Cortical|8370/3
C0206686|T191|PM|D018268|MSH|Carcinomas, Adrenocortical|8370/3
C0206686|T191|PN|NOCODE|MTH|Adrenocortical carcinoma|8370/3
C0206686|T191|SY|C9325|NCI|Adrenal Cortex Adenocarcinoma|8370/3
C0206686|T191|SY|C9325|NCI|Adrenal Cortex Cancer|8370/3
C0206686|T191|PT|C9325|NCI|Adrenal Cortex Carcinoma|8370/3
C0206686|T191|SY|TCGA|NCI|Adrenal Cortex Carcinoma|8370/3
C0206686|T191|SY|C9325|NCI|Adrenal Cortical Adenocarcinoma|8370/3
C0206686|T191|SY|C9325|NCI|Adrenal Cortical Carcinoma|8370/3
C0206686|T191|SY|C9325|NCI|Adrenocortical Carcinoma|8370/3
C0206686|T191|SY|C9325|NCI|Carcinoma of Adrenal Cortex|8370/3
C0206686|T191|SY|C9325|NCI|Carcinoma of the Adrenal Cortex|8370/3
C0206686|T191|SY|C9325|NCI_CDISC|Adenocarcinoma, Adrenocortical, Malignant|8370/3
C0206686|T191|SY|C9325|NCI_CDISC|Adrenal Cortex Adenocarcinoma|8370/3
C0206686|T191|SY|C9325|NCI_CDISC|Adrenal Cortex Cancer|8370/3
C0206686|T191|SY|C9325|NCI_CDISC|Adrenal Cortical Adenocarcinoma|8370/3
C0206686|T191|SY|C9325|NCI_CDISC|Adrenal Cortical Carcinoma|8370/3
C0206686|T191|SY|C9325|NCI_CDISC|Adrenocortical Carcinoma|8370/3
C0206686|T191|PT|C9325|NCI_CDISC|CARCINOMA, ADRENOCORTICAL, MALIGNANT|8370/3
C0206686|T191|SY|C9325|NCI_CDISC|Cortical Cell Carcinoma|8370/3
C0206686|T191|PT|C9325|NCI_CPTAC|Adrenal Cortex Carcinoma|8370/3
C0206686|T191|SY|10001327|NCI_CTEP-SDC|Adrenocortical carcinoma|8370/3
C0206686|T191|PT|10001327|NCI_CTEP-SDC|Adrenocortical carcinoma, NOS|8370/3
C0206686|T191|DN|C9325|NCI_CTRP|Adrenal Cortex Cancer|8370/3
C0206686|T191|PT|C9325|NCI_CTRP|Adrenal Cortex Cancer|8370/3
C0206686|T191|SY|C9325|NCI_CTRP|Adrenal Cortex Carcinoma|8370/3
C0206686|T191|PT|CDR0000457974|NCI_NCI-GLOSS|adrenocortical cancer|8370/3
C0206686|T191|PT|CDR0000446526|NCI_NCI-GLOSS|adrenocortical carcinoma|8370/3
C0206686|T191|PT|CDR0000457975|NCI_NCI-GLOSS|cancer of the adrenal cortex|8370/3
C0206686|T191|SY|CDR0000038758|PDQ|adrenal cortical carcinoma|8370/3
C0206686|T191|ET|CDR0000038758|PDQ|Adrenocortical carcinoma|8370/3
C0206686|T191|PSC|CDR0000038758|PDQ|adrenocortical carcinoma|8370/3
C0206686|T191|SY|CDR0000038758|PDQ|carcinoma, adrenocortical|8370/3
C0206686|T191|PT|X78ca|RCD|Adrenal carcinoma|8370/3
C0206686|T191|AB|X78ca|RCD|Adrenal cortical adenoca|8370/3
C0206686|T191|SY|X78ca|RCD|Adrenal cortical adenocarcinoma|8370/3
C0206686|T191|OP|BB5h1|RCD|Adrenal cortical carcinoma|8370/3
C0206686|T191|PT|255035007|SNOMEDCT_US|Adrenal carcinoma|8370/3
C0206686|T191|SY|255035007|SNOMEDCT_US|Adrenal cortical adenocarcinoma|8370/3
C0206686|T191|SY|2227007|SNOMEDCT_US|Adrenal cortical adenocarcinoma|8370/3
C0206686|T191|PT|2227007|SNOMEDCT_US|Adrenal cortical carcinoma|8370/3
C0334332|T191|PN|NOCODE|MTH|Compact Cell Adrenal Cortical Adenoma|8371/0
C0334332|T191|PT|C4163|NCI|Adrenal Cortex Compact Cell Adenoma|8371/0
C0334332|T191|SY|C4163|NCI|Compact Cell Adrenal Cortex Adenoma|8371/0
C0334332|T191|SY|C4163|NCI|Compact Cell Adrenal Cortical Adenoma|8371/0
C0334332|T191|SY|C4163|NCI|Compact Cell Adrenocortical Adenoma|8371/0
C0334332|T191|AB|BB5h2|RCD|Adren cort adenom-compact cell|8371/0
C0334332|T191|PT|BB5h2|RCD|Adrenal cortical adenoma - compact cell|8371/0
C0334332|T191|SY|63687009|SNOMEDCT_US|Adrenal cortical adenoma - compact cell|8371/0
C0334332|T191|PT|63687009|SNOMEDCT_US|Adrenal cortical adenoma, compact cell|8371/0
C0334333|T191|PT|MTHU003531|ICPC2ICD10ENG|adenoma; black|8372/0
C0334333|T191|PT|MTHU084139|ICPC2ICD10ENG|black; adenoma|8372/0
C0334333|T191|PN|NOCODE|MTH|Heavily Pigmented Adrenal Cortical Adenoma|8372/0
C0334333|T191|SY|C4164|NCI|Black Adenoma|8372/0
C0334333|T191|SY|C4164|NCI|Heavily Pigmented Adrenal Cortex Adenoma|8372/0
C0334333|T191|SY|C4164|NCI|Heavily Pigmented Adrenal Cortical Adenoma|8372/0
C0334333|T191|SY|C4164|NCI|Heavily Pigmented Adrenocortical Adenoma|8372/0
C0334333|T191|PT|C4164|NCI|Pigmented Adrenal Cortex Adenoma|8372/0
C0334333|T191|AB|BB5h3|RCD|Adr cort adenom-heavy pigment|8372/0
C0334333|T191|PT|BB5h3|RCD|Adrenal cortical adenoma - heavily pigmented variant|8372/0
C0334333|T191|SY|BB5h3|RCD|Black adenoma|8372/0
C0334333|T191|SY|37302003|SNOMEDCT_US|Adrenal cortical adenoma - heavily pigmented variant|8372/0
C0334333|T191|SY|37302003|SNOMEDCT_US|Adrenal cortical adenoma, heavily pigmented variant|8372/0
C0334333|T191|PT|37302003|SNOMEDCT_US|Adrenal cortical adenoma, pigmented|8372/0
C0334333|T191|SY|37302003|SNOMEDCT_US|Black adenoma|8372/0
C0334333|T191|SY|37302003|SNOMEDCT_US|Pigmented adenoma|8372/0
C0334334|T191|PN|NOCODE|MTH|Clear Cell Adrenal Cortical Adenoma|8373/0
C0334334|T191|PT|C4165|NCI|Adrenal Cortex Clear Cell Adenoma|8373/0
C0334334|T191|SY|C4165|NCI|Clear Cell Adrenal Cortex Adenoma|8373/0
C0334334|T191|SY|C4165|NCI|Clear Cell Adrenal Cortical Adenoma|8373/0
C0334334|T191|SY|C4165|NCI|Clear Cell Adrenocortical Adenoma|8373/0
C0334334|T191|AB|BB5h4|RCD|Adren cort adenoma-clear cell|8373/0
C0334334|T191|PT|BB5h4|RCD|Adrenal cortical adenoma - clear cell|8373/0
C0334334|T191|SY|18977007|SNOMEDCT_US|Adrenal cortical adenoma - clear cell|8373/0
C0334334|T191|PT|18977007|SNOMEDCT_US|Adrenal cortical adenoma, clear cell|8373/0
C0334335|T191|PN|NOCODE|MTH|Glomerulosa Cell Adrenal Cortical Adenoma|8374/0
C0334335|T191|PT|C4166|NCI|Adrenal Cortex Glomerulosa Cell Adenoma|8374/0
C0334335|T191|SY|C4166|NCI|Glomerulosa Cell Adrenal Cortex Adenoma|8374/0
C0334335|T191|SY|C4166|NCI|Glomerulosa Cell Adrenal Cortical Adenoma|8374/0
C0334335|T191|SY|C4166|NCI|Glomerulosa Cell Adrenocortical Adenoma|8374/0
C0334335|T191|AB|BB5h5|RCD|Adr cort aden-glomerulosa cell|8374/0
C0334335|T191|PT|BB5h5|RCD|Adrenal cortical adenoma - glomerulosa cell|8374/0
C0334335|T191|SY|19329008|SNOMEDCT_US|Adrenal cortical adenoma - glomerulosa cell|8374/0
C0334335|T191|PT|19329008|SNOMEDCT_US|Adrenal cortical adenoma, glomerulosa cell|8374/0
C0334336|T191|PN|NOCODE|MTH|Mixed Cell Adrenal Cortical Adenoma|8375/0
C0334336|T191|PT|C4167|NCI|Adrenal Cortex Mixed Cell Adenoma|8375/0
C0334336|T191|SY|C4167|NCI|Mixed Cell Adrenal Cortex Adenoma|8375/0
C0334336|T191|SY|C4167|NCI|Mixed Cell Adrenal Cortical Adenoma|8375/0
C0334336|T191|SY|C4167|NCI|Mixed Cell Adrenocortical Adenoma|8375/0
C0334336|T191|AB|BB5h6|RCD|Adren cort adenoma-mixed cell|8375/0
C0334336|T191|PT|BB5h6|RCD|Adrenal cortical adenoma - mixed cell|8375/0
C0334336|T191|SY|39720002|SNOMEDCT_US|Adrenal cortical adenoma - mixed cell|8375/0
C0334336|T191|PT|39720002|SNOMEDCT_US|Adrenal cortical adenoma, mixed cell|8375/0
C2212024|T191|PT|233198|MEDCIN|endometrioid adenofibroma of ovary|8380/0
C2212024|T191|PT|C27287|NCI|Ovarian Endometrioid Adenofibroma|8380/0
C0334337|T191|PT|Xa98U|RCD|Endometrioid adenoma|8380/0
C0334337|T191|SY|Xa98U|RCD|Endometrioid cystadenoma|8380/0
C0334337|T191|SY|Xa98U|RCDSY|Endometrioid adenoma NOS|8380/0
C0334337|T191|OAP|189650001|SNOMEDCT_US|Endometrioid adenoma|8380/0
C0334337|T191|OF|189650001|SNOMEDCT_US|Endometrioid adenoma|8380/0
C0334337|T191|PT|71106006|SNOMEDCT_US|Endometrioid adenoma|8380/0
C0334337|T191|IS|71106006|SNOMEDCT_US|Endometrioid adenoma, NOS|8380/0
C0334337|T191|SY|71106006|SNOMEDCT_US|Endometrioid cystadenoma|8380/0
C0334337|T191|IS|71106006|SNOMEDCT_US|Endometrioid cystadenoma, NOS|8380/0
C0334338|T191|PT|MTHU003426|ICPC2ICD10ENG|adenofibroma; endometrioid, borderline malignancy|8380/1
C0334338|T191|PT|MTHU012112|ICPC2ICD10ENG|borderline malignancy; endometrioid adenofibroma|8380/1
C0334338|T191|PT|MTHU012113|ICPC2ICD10ENG|borderline malignancy; endometrioid cystadenofibroma|8380/1
C0334338|T191|PT|MTHU020303|ICPC2ICD10ENG|cystadenofibroma; endometrioid, borderline malignancy|8380/1
C0334338|T191|PT|MTHU026102|ICPC2ICD10ENG|endometrioid; adenofibroma, borderline malignancy|8380/1
C0334338|T191|PT|MTHU026109|ICPC2ICD10ENG|endometrioid; cystadenofibroma, borderline malignancy|8380/1
C0334338|T191|SY|C7983|NCI|Borderline Endometrioid Neoplasm of Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Borderline Endometrioid Neoplasm of the Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Borderline Endometrioid Tumor of Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Borderline Endometrioid Tumor of the Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Borderline Ovarian Endometrioid Neoplasm|8380/1
C0334338|T191|SY|C7983|NCI|Borderline Ovarian Endometrioid Tumor|8380/1
C0334338|T191|PT|C7983|NCI|Borderline Ovarian Endometrioid Tumor/Atypical Proliferative Ovarian Endometrioid Tumor|8380/1
C0334338|T191|AB|C7983|NCI|EBT/APET|8380/1
C0334338|T191|SY|C7983|NCI|Endometrioid Neoplasm of Low Malignant Potential|8380/1
C0334338|T191|SY|C7983|NCI|Endometrioid Neoplasm with Proliferating Activity, Ovarian|8380/1
C0334338|T191|SY|C7983|NCI|Endometrioid Tumor of Low Malignant Potential|8380/1
C0334338|T191|SY|C7983|NCI|Endometrioid Tumor with Proliferating Activity, Ovarian|8380/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Endometrioid Neoplasm of Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Endometrioid Neoplasm of the Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Endometrioid Tumor of Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Endometrioid Tumor of the Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Ovarian Endometrioid Neoplasm|8380/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Ovarian Endometrioid Tumor|8380/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Borderline Neoplasm|8380/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Borderline Tumor|8380/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Neoplasm of Low Malignant Potential|8380/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Neoplasm with Proliferating Activity|8380/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Tumor of Low Malignant Potential|8380/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Tumor with Proliferating Activity|8380/1
C0334338|T191|SY|C7983|NCI|Proliferating Endometrioid Neoplasm of Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Proliferating Endometrioid Neoplasm of the Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Proliferating Endometrioid Tumor of Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Proliferating Endometrioid Tumor of the Ovary|8380/1
C0334338|T191|SY|C7983|NCI|Proliferating Ovarian Endometrioid Neoplasm|8380/1
C0334338|T191|SY|C7983|NCI|Proliferating Ovarian Endometrioid Tumor|8380/1
C0334338|T191|DN|C7983|NCI_CTRP|Borderline Ovarian Endometrioid Tumor/Atypical Proliferative Ovarian Endometrioid Tumor|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Adenofibroma|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Cystadenoma|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Neoplasm of Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Neoplasm of the Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Tumor of Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Tumor of the Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Malignancy Endometrioid Adenofibroma|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Malignancy Endometrioid Cystadenoma|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Ovarian Endometrioid Neoplasm|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Ovarian Endometrioid Tumor|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Endometrioid Neoplasm of Low Malignant Potential|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Endometrioid Neoplasm with Proliferating Activity, Ovarian|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Endometrioid Tumor of Low Malignant Potential|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|endometrioid tumor with proliferating activity, ovarian|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignancy Potential Endometrioid Cystadenoma|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Endometrioid Neoplasm of Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Endometrioid Neoplasm of the Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Endometrioid Tumor of Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Endometrioid Tumor of the Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Ovarian Endometrioid Neoplasm|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Ovarian Endometrioid Tumor|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Borderline Neoplasm|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Borderline Tumor|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Neoplasm of Low Malignant Potential|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Neoplasm with Proliferating Activity|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Tumor of Low Malignant Potential|8380/1
C0334338|T191|PT|CDR0000039965|PDQ|ovarian endometrioid tumor with proliferating activity|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Endometrioid Neoplasm of Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Endometrioid Neoplasm of the Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Endometrioid Tumor of Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Endometrioid Tumor of the Ovary|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Ovarian Endometrioid Neoplasm|8380/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Ovarian Endometrioid Tumor|8380/1
C0334338|T191|AB|BB5j4|RCD|Endom adenofibroma-bord malig|8380/1
C0334338|T191|AB|BB5j4|RCD|Endom cystadenofibrom-bord mal|8380/1
C0334338|T191|AB|BB5j1|RCD|Endom cystadoma-bordline malig|8380/1
C0334338|T191|AB|BB5j1|RCD|Endom tumour low malig potent|8380/1
C0334338|T191|AB|BB5j1|RCD|Endomet adenoma-bordline malig|8380/1
C0334338|T191|PT|BB5j4|RCD|Endometrioid adenofibroma - borderline malignancy|8380/1
C0334338|T191|PT|BB5j1|RCD|Endometrioid adenoma - borderline malignancy|8380/1
C0334338|T191|SY|BB5j4|RCD|Endometrioid cystadenofibroma - borderline malignancy|8380/1
C0334338|T191|SY|BB5j1|RCD|Endometrioid cystadenoma - borderline malignancy|8380/1
C0334338|T191|SY|BB5j1|RCD|Endometrioid tumour of low malignant potential|8380/1
C0334338|T191|AB|BB5j1|RCDAE|Endom tumor low malig potent|8380/1
C0334338|T191|SY|BB5j1|RCDAE|Endometrioid tumor of low malignant potential|8380/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Atypical proliferative endometrioid tumor|8380/1
C0334338|T191|SYGB|75987005|SNOMEDCT_US|Atypical proliferative endometrioid tumour|8380/1
C0334338|T191|SY|25874003|SNOMEDCT_US|Endometrioid adenofibroma - borderline malignancy|8380/1
C0334338|T191|PT|25874003|SNOMEDCT_US|Endometrioid adenofibroma, borderline malignancy|8380/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid adenoma - borderline malignancy|8380/1
C0334338|T191|PT|75987005|SNOMEDCT_US|Endometrioid adenoma, borderline malignancy|8380/1
C0334338|T191|SY|25874003|SNOMEDCT_US|Endometrioid cystadenofibroma - borderline malignancy|8380/1
C0334338|T191|SY|25874003|SNOMEDCT_US|Endometrioid cystadenofibroma, borderline malignancy|8380/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid cystadenoma - borderline malignancy|8380/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid cystadenoma, borderline malignancy|8380/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid tumor of low malignant potential|8380/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid tumor, borderline|8380/1
C0334338|T191|SYGB|75987005|SNOMEDCT_US|Endometrioid tumour of low malignant potential|8380/1
C0334338|T191|SYGB|75987005|SNOMEDCT_US|Endometrioid tumour, borderline|8380/1
C3812874|T191|LLT|10079951|MDR|Endometrioid intraepithelial neoplasia|8380/2
C3812874|T191|PN|NOCODE|MTH|Endometrioid intraepithelial neoplasia|8380/2
C3812874|T191|SY|703548001|SNOMEDCT_US|Atypical hyperplasia of the endometrium|8380/2
C3812874|T191|PT|703548001|SNOMEDCT_US|Endometrioid intraepithelial neoplasia|8380/2
C0206687|T191|PT|0011175|CCPSS|ENDOMETRIOID CARCINOMA|8380/3
C0206687|T191|SY|0000021021|CHV|carcinoma endometrioid|8380/3
C0206687|T191|SY|0000021021|CHV|endometrioid adenocarcinoma|8380/3
C0206687|T191|PT|0000021021|CHV|endometrioid carcinoma|8380/3
C0206687|T191|PT|MTHU014750|ICPC2ICD10ENG|carcinoma; endometrioid, unspecified site, female|8380/3
C0206687|T191|PT|MTHU026105|ICPC2ICD10ENG|endometrioid; carcinoma, unspecified site, female|8380/3
C0206687|T191|PT|271450|MEDCIN|endometrioid carcinoma|8380/3
C0206687|T191|MH|D018269|MSH|Carcinoma, Endometrioid|8380/3
C0206687|T191|PM|D018269|MSH|Carcinomas, Endometrioid|8380/3
C0206687|T191|PM|D018269|MSH|Endometrioid Carcinoma|8380/3
C0206687|T191|PM|D018269|MSH|Endometrioid Carcinomas|8380/3
C0206687|T191|PN|NOCODE|MTH|Carcinoma, Endometrioid|8380/3
C0206687|T191|PT|C3769|NCI|Endometrioid Adenocarcinoma|8380/3
C0206687|T191|SY|TCGA|NCI|Endometrioid Adenocarcinoma|8380/3
C0206687|T191|SY|C3769|NCI|Endometrioid Carcinoma|8380/3
C0206687|T191|SY|C3769|NCI|Endometrioid Carcinoma of Female Reproductive System|8380/3
C0206687|T191|SY|C3769|NCI|Endometrioid Carcinoma of the Female Reproductive System|8380/3
C0206687|T191|SY|C3769|NCI|Female Reproductive Endometrioid Carcinoma|8380/3
C0206687|T191|PT|BB5j2|RCD|Endometrioid carcinoma|8380/3
C0206687|T191|PT|30289006|SNOMEDCT_US|Endometrioid carcinoma|8380/3
C0334339|T191|PT|MTHU003425|ICPC2ICD10ENG|adenofibroma; endometrioid|8381/0
C0334339|T191|PT|MTHU020302|ICPC2ICD10ENG|cystadenofibroma; endometrioid|8381/0
C0334339|T191|PT|MTHU026101|ICPC2ICD10ENG|endometrioid; adenofibroma|8381/0
C0334339|T191|PT|MTHU026108|ICPC2ICD10ENG|endometrioid; cystadenofibroma|8381/0
C2212024|T191|PT|233198|MEDCIN|endometrioid adenofibroma of ovary|8381/0
C2212024|T191|PT|C27287|NCI|Ovarian Endometrioid Adenofibroma|8381/0
C0334339|T191|PT|Xa98V|RCD|Endometrioid adenofibroma|8381/0
C0334339|T191|SY|Xa98V|RCD|Endometrioid cystadenofibroma|8381/0
C0334339|T191|OA|BB5j3|RCDSY|Endometrioid adenofibr.NOS|8381/0
C0334339|T191|OP|BB5j3|RCDSY|Endometrioid adenofibroma NOS|8381/0
C0334339|T191|PT|20829008|SNOMEDCT_US|Endometrioid adenofibroma|8381/0
C0334339|T191|IS|20829008|SNOMEDCT_US|Endometrioid adenofibroma, NOS|8381/0
C0334339|T191|SY|20829008|SNOMEDCT_US|Endometrioid cystadenofibroma|8381/0
C0334339|T191|IS|20829008|SNOMEDCT_US|Endometrioid cystadenofibroma, NOS|8381/0
C0334338|T191|PT|MTHU003426|ICPC2ICD10ENG|adenofibroma; endometrioid, borderline malignancy|8381/1
C0334338|T191|PT|MTHU012112|ICPC2ICD10ENG|borderline malignancy; endometrioid adenofibroma|8381/1
C0334338|T191|PT|MTHU012113|ICPC2ICD10ENG|borderline malignancy; endometrioid cystadenofibroma|8381/1
C0334338|T191|PT|MTHU020303|ICPC2ICD10ENG|cystadenofibroma; endometrioid, borderline malignancy|8381/1
C0334338|T191|PT|MTHU026102|ICPC2ICD10ENG|endometrioid; adenofibroma, borderline malignancy|8381/1
C0334338|T191|PT|MTHU026109|ICPC2ICD10ENG|endometrioid; cystadenofibroma, borderline malignancy|8381/1
C0334338|T191|SY|C7983|NCI|Borderline Endometrioid Neoplasm of Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Borderline Endometrioid Neoplasm of the Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Borderline Endometrioid Tumor of Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Borderline Endometrioid Tumor of the Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Borderline Ovarian Endometrioid Neoplasm|8381/1
C0334338|T191|SY|C7983|NCI|Borderline Ovarian Endometrioid Tumor|8381/1
C0334338|T191|PT|C7983|NCI|Borderline Ovarian Endometrioid Tumor/Atypical Proliferative Ovarian Endometrioid Tumor|8381/1
C0334338|T191|AB|C7983|NCI|EBT/APET|8381/1
C0334338|T191|SY|C7983|NCI|Endometrioid Neoplasm of Low Malignant Potential|8381/1
C0334338|T191|SY|C7983|NCI|Endometrioid Neoplasm with Proliferating Activity, Ovarian|8381/1
C0334338|T191|SY|C7983|NCI|Endometrioid Tumor of Low Malignant Potential|8381/1
C0334338|T191|SY|C7983|NCI|Endometrioid Tumor with Proliferating Activity, Ovarian|8381/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Endometrioid Neoplasm of Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Endometrioid Neoplasm of the Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Endometrioid Tumor of Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Endometrioid Tumor of the Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Ovarian Endometrioid Neoplasm|8381/1
C0334338|T191|SY|C7983|NCI|Low Malignant Potential Ovarian Endometrioid Tumor|8381/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Borderline Neoplasm|8381/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Borderline Tumor|8381/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Neoplasm of Low Malignant Potential|8381/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Neoplasm with Proliferating Activity|8381/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Tumor of Low Malignant Potential|8381/1
C0334338|T191|SY|C7983|NCI|Ovarian Endometrioid Tumor with Proliferating Activity|8381/1
C0334338|T191|SY|C7983|NCI|Proliferating Endometrioid Neoplasm of Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Proliferating Endometrioid Neoplasm of the Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Proliferating Endometrioid Tumor of Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Proliferating Endometrioid Tumor of the Ovary|8381/1
C0334338|T191|SY|C7983|NCI|Proliferating Ovarian Endometrioid Neoplasm|8381/1
C0334338|T191|SY|C7983|NCI|Proliferating Ovarian Endometrioid Tumor|8381/1
C0334338|T191|DN|C7983|NCI_CTRP|Borderline Ovarian Endometrioid Tumor/Atypical Proliferative Ovarian Endometrioid Tumor|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Adenofibroma|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Cystadenoma|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Neoplasm of Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Neoplasm of the Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Tumor of Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Endometrioid Tumor of the Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Malignancy Endometrioid Adenofibroma|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Malignancy Endometrioid Cystadenoma|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Ovarian Endometrioid Neoplasm|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Borderline Ovarian Endometrioid Tumor|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Endometrioid Neoplasm of Low Malignant Potential|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Endometrioid Neoplasm with Proliferating Activity, Ovarian|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Endometrioid Tumor of Low Malignant Potential|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|endometrioid tumor with proliferating activity, ovarian|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignancy Potential Endometrioid Cystadenoma|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Endometrioid Neoplasm of Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Endometrioid Neoplasm of the Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Endometrioid Tumor of Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Endometrioid Tumor of the Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Ovarian Endometrioid Neoplasm|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Low Malignant Potential Ovarian Endometrioid Tumor|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Borderline Neoplasm|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Borderline Tumor|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Neoplasm of Low Malignant Potential|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Neoplasm with Proliferating Activity|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Ovarian Endometrioid Tumor of Low Malignant Potential|8381/1
C0334338|T191|PT|CDR0000039965|PDQ|ovarian endometrioid tumor with proliferating activity|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Endometrioid Neoplasm of Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Endometrioid Neoplasm of the Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Endometrioid Tumor of Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Endometrioid Tumor of the Ovary|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Ovarian Endometrioid Neoplasm|8381/1
C0334338|T191|SY|CDR0000039965|PDQ|Proliferating Ovarian Endometrioid Tumor|8381/1
C0334338|T191|AB|BB5j4|RCD|Endom adenofibroma-bord malig|8381/1
C0334338|T191|AB|BB5j4|RCD|Endom cystadenofibrom-bord mal|8381/1
C0334338|T191|AB|BB5j1|RCD|Endom cystadoma-bordline malig|8381/1
C0334338|T191|AB|BB5j1|RCD|Endom tumour low malig potent|8381/1
C0334338|T191|AB|BB5j1|RCD|Endomet adenoma-bordline malig|8381/1
C0334338|T191|PT|BB5j4|RCD|Endometrioid adenofibroma - borderline malignancy|8381/1
C0334338|T191|PT|BB5j1|RCD|Endometrioid adenoma - borderline malignancy|8381/1
C0334338|T191|SY|BB5j4|RCD|Endometrioid cystadenofibroma - borderline malignancy|8381/1
C0334338|T191|SY|BB5j1|RCD|Endometrioid cystadenoma - borderline malignancy|8381/1
C0334338|T191|SY|BB5j1|RCD|Endometrioid tumour of low malignant potential|8381/1
C0334338|T191|AB|BB5j1|RCDAE|Endom tumor low malig potent|8381/1
C0334338|T191|SY|BB5j1|RCDAE|Endometrioid tumor of low malignant potential|8381/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Atypical proliferative endometrioid tumor|8381/1
C0334338|T191|SYGB|75987005|SNOMEDCT_US|Atypical proliferative endometrioid tumour|8381/1
C0334338|T191|SY|25874003|SNOMEDCT_US|Endometrioid adenofibroma - borderline malignancy|8381/1
C0334338|T191|PT|25874003|SNOMEDCT_US|Endometrioid adenofibroma, borderline malignancy|8381/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid adenoma - borderline malignancy|8381/1
C0334338|T191|PT|75987005|SNOMEDCT_US|Endometrioid adenoma, borderline malignancy|8381/1
C0334338|T191|SY|25874003|SNOMEDCT_US|Endometrioid cystadenofibroma - borderline malignancy|8381/1
C0334338|T191|SY|25874003|SNOMEDCT_US|Endometrioid cystadenofibroma, borderline malignancy|8381/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid cystadenoma - borderline malignancy|8381/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid cystadenoma, borderline malignancy|8381/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid tumor of low malignant potential|8381/1
C0334338|T191|SY|75987005|SNOMEDCT_US|Endometrioid tumor, borderline|8381/1
C0334338|T191|SYGB|75987005|SNOMEDCT_US|Endometrioid tumour of low malignant potential|8381/1
C0334338|T191|SYGB|75987005|SNOMEDCT_US|Endometrioid tumour, borderline|8381/1
C0334341|T191|PT|MTHU003427|ICPC2ICD10ENG|adenofibroma; endometrioid, malignant|8381/3
C0334341|T191|PT|MTHU020304|ICPC2ICD10ENG|cystadenofibroma; endometrioid, malignant|8381/3
C0334341|T191|PT|MTHU026103|ICPC2ICD10ENG|endometrioid; adenofibroma, malignant|8381/3
C0334341|T191|PT|MTHU026110|ICPC2ICD10ENG|endometrioid; cystadenofibroma, malignant|8381/3
C1518711|T191|PT|C40060|NCI|Ovarian Endometrioid Adenocarcinofibroma|8381/3
C1518711|T191|OP|C40060|NCI|Ovarian Endometrioid Adenocarcinofibroma|8381/3
C1518711|T191|OP|C40060|NCI|Ovarian Endometrioid Malignant Adenofibroma|8381/3
C0334341|T191|AB|BB5j5|RCD|Malig endomet cystadenofibroma|8381/3
C0334341|T191|AB|BB5j5|RCD|Malig endometr adenofibroma|8381/3
C0334341|T191|PT|BB5j5|RCD|Malignant endometrioid adenofibroma|8381/3
C0334341|T191|SY|BB5j5|RCD|Malignant endometrioid cystadenofibroma|8381/3
C0334341|T191|PT|18105004|SNOMEDCT_US|Endometrioid adenofibroma, malignant|8381/3
C0334341|T191|SY|18105004|SNOMEDCT_US|Endometrioid cystadenofibroma, malignant|8381/3
C0334341|T191|SY|18105004|SNOMEDCT_US|Malignant endometrioid adenofibroma|8381/3
C0334341|T191|SY|18105004|SNOMEDCT_US|Malignant endometrioid cystadenofibroma|8381/3
C1336907|T191|PT|C27839|NCI|Endometrial Endometrioid Adenocarcinoma, Secretory Variant|8382/3
C1336907|T191|SY|C27839|NCI|Secretory Uterine Corpus Endometrioid Adenocarcinoma|8382/3
C1266057|T191|PT|128680006|SNOMEDCT_US|Endometrioid adenocarcinoma, secretory variant|8382/3
C1336906|T191|SY|C27848|NCI|Ciliated Uterine Corpus Endometrioid Adenocarcinoma|8383/3
C1336906|T191|PT|C27848|NCI|Endometrial Endometrioid Adenocarcinoma, Ciliated Variant|8383/3
C1266058|T191|PT|128681005|SNOMEDCT_US|Endometrioid adenocarcinoma, ciliated cell variant|8383/3
C1272765|T191|PT|355656|MEDCIN|Adenoma malignum|8384/3
C1272765|T191|SY|355656|MEDCIN|cervical adenocarcinoma adenoma malignum|8384/3
C1266059|T191|PT|C66951|NCI|Adenocarcinoma, Endocervical Type|8384/3
C1266059|T191|PT|128682003|SNOMEDCT_US|Adenocarcinoma, endocervical type|8384/3
C1272765|T191|PT|385478001|SNOMEDCT_US|Adenoma malignum|8384/3
C1272765|T191|SY|388986005|SNOMEDCT_US|Adenoma malignum|8384/3
C1272765|T191|PT|388986005|SNOMEDCT_US|Minimal deviation adenocarcinoma of endocervical type|8384/3
C0334342|T191|PT|0000029959|CHV|adnexal tumor|8390/0
C0334342|T191|SY|0000029959|CHV|adnexal tumors|8390/0
C0334342|T191|SY|0000029959|CHV|adnexal tumour|8390/0
C0334342|T191|SY|0000029959|CHV|adnexal tumours|8390/0
C0334342|T191|SY|C7580|NCI|Adenoma of Adnexa|8390/0
C0334342|T191|SY|C7580|NCI|Adenoma of Skin Appendage|8390/0
C0334342|T191|SY|C7580|NCI|Adnexal Adenoma|8390/0
C0334342|T191|PT|C7580|NCI|Skin Appendage Adenoma|8390/0
C0334342|T191|SY|C7580|NCI_CDISC|Adenoma of Adnexa|8390/0
C0334342|T191|SY|C7580|NCI_CDISC|Adenoma of Skin Appendage|8390/0
C0334342|T191|PT|C7580|NCI_CDISC|ADENOMA, ADNEXAL, BENIGN|8390/0
C0334342|T191|SY|C7580|NCI_CDISC|Adnexal Adenoma|8390/0
C0334342|T191|SY|XM1FH|RCD|Adnexal tumour|8390/0
C0334342|T191|PT|XM1FH|RCD|Skin appendage adenoma|8390/0
C0334342|T191|SY|XM1FH|RCDAE|Adnexal tumor|8390/0
C0334342|T191|OP|BB600|RCDSY|Skin appendage adenoma|8390/0
C0334342|T191|SY|55681005|SNOMEDCT_US|Adnexal tumor|8390/0
C0334342|T191|SYGB|55681005|SNOMEDCT_US|Adnexal tumour|8390/0
C0334342|T191|PT|55681005|SNOMEDCT_US|Skin appendage adenoma|8390/0
C0206697|T191|PT|0000021029|CHV|adnexal carcinoma|8390/3
C0206697|T191|PT|231625|MEDCIN|skin appendage carcinoma|8390/3
C0206697|T191|PM|D018280|MSH|Appendage Carcinoma, Skin|8390/3
C0206697|T191|PM|D018280|MSH|Appendage Carcinomas, Skin|8390/3
C0206697|T191|MH|D018280|MSH|Carcinoma, Skin Appendage|8390/3
C0206697|T191|PM|D018280|MSH|Carcinomas, Skin Appendage|8390/3
C0206697|T191|PM|D018280|MSH|Skin Appendage Carcinoma|8390/3
C0206697|T191|PM|D018280|MSH|Skin Appendage Carcinomas|8390/3
C0206697|T191|PT|C3775|NCI|Adnexal Carcinoma|8390/3
C0206697|T191|SY|C3775|NCI|Carcinoma of Adnexa|8390/3
C0206697|T191|SY|C3775|NCI|Carcinoma of Skin Appendage|8390/3
C0206697|T191|SY|C3775|NCI|Skin Appendage Carcinoma|8390/3
C0206697|T191|SY|C3775|NCI_CDISC|Carcinoma of Adnexa|8390/3
C0206697|T191|SY|C3775|NCI_CDISC|Carcinoma of Skin Appendage|8390/3
C0206697|T191|PT|C3775|NCI_CDISC|CARCINOMA, ADNEXAL, MALIGNANT|8390/3
C0206697|T191|SY|C3775|NCI_CDISC|Skin Appendage Carcinoma|8390/3
C0206697|T191|SY|XM1FI|RCD|Adnexal carcinoma|8390/3
C0206697|T191|PT|XM1FI|RCD|Skin appendage carcinoma|8390/3
C0206697|T191|OP|BB601|RCDSY|Skin appendage carcinoma|8390/3
C0206697|T191|SY|64000002|SNOMEDCT_US|Adnexal carcinoma|8390/3
C0206697|T191|PT|64000002|SNOMEDCT_US|Skin appendage carcinoma|8390/3
C0346011|T191|SY|0000031040|CHV|fibrofolliculoma|8391/0
C0346011|T191|PT|0000031040|CHV|fibrofolliculomas|8391/0
C0346011|T191|SY|0000031040|CHV|trichodiscoma|8391/0
C0346011|T191|PT|HP:0030436|HPO|Fibrofolliculoma|8391/0
C0346011|T191|SY|HP:0030436|HPO|Fibrofolliculomas|8391/0
C0346011|T191|PN|NOCODE|MTH|Fibrofolliculoma|8391/0
C0346011|T191|PT|C43331|NCI|Fibrofolliculoma|8391/0
C0346011|T191|PT|X78SP|RCD|Fibrofolliculoma|8391/0
C0346011|T191|PT|254699007|SNOMEDCT_US|Fibrofolliculoma|8391/0
C0346011|T191|SY|128683008|SNOMEDCT_US|Fibrofolliculoma|8391/0
C0346011|T191|OAP|110984002|SNOMEDCT_US|Fibrofolliculoma|8391/0
C0346011|T191|PT|128683008|SNOMEDCT_US|Follicular fibroma|8391/0
C1266060|T191|SY|HP:0031018|HPO|Acrosyringeal adenomatosis|8392/0
C1266060|T191|PT|HP:0031018|HPO|Eccrine syringofibroadenoma|8392/0
C1266060|T191|SY|HP:0031018|HPO|Eccrine syringofibroadenomatous hyperplasia|8392/0
C1266060|T191|SY|HP:0031018|HPO|Syringofibroadenoma|8392/0
C1266060|T191|PEP|D057091|MSH|Syringofibroadenoma|8392/0
C1266060|T191|PM|D057091|MSH|Syringofibroadenomas|8392/0
C1266060|T191|SY|C43356|NCI|Acrosyringeal Adenomatosis|8392/0
C1266060|T191|SY|C43356|NCI|Acrosyringeal Nevus|8392/0
C1266060|T191|SY|C43356|NCI|Eccrine Poromatosis|8392/0
C1266060|T191|PT|C43356|NCI|Eccrine Syringofibroadenoma|8392/0
C1266060|T191|SY|C43356|NCI|Eccrine Syringofibroadenoma of Mascaro|8392/0
C1266060|T191|SY|C43356|NCI|Linear Eccrine Poroma|8392/0
C1266060|T191|SY|C43356|NCI|Nevus Syringoadenomatosus Papilliferum|8392/0
C1266060|T191|SY|C43356|NCI|Syringofibroadenoma|8392/0
C1266060|T191|PT|X50Jb|RCD|Acrosyringeal naevus|8392/0
C1266060|T191|PT|X50Jb|RCDAE|Acrosyringeal nevus|8392/0
C1266060|T191|PTGB|239117002|SNOMEDCT_US|Acrosyringeal naevus|8392/0
C1266060|T191|PT|239117002|SNOMEDCT_US|Acrosyringeal nevus|8392/0
C1266060|T191|PT|403936002|SNOMEDCT_US|Eccrine syringofibroadenoma|8392/0
C1266060|T191|SY|403936002|SNOMEDCT_US|Eccrine syringofibroadenoma of skin|8392/0
C1266060|T191|PT|128684002|SNOMEDCT_US|Syringofibroadenoma|8392/0
C1266060|T191|SY|403936002|SNOMEDCT_US|Syringofibroadenoma|8392/0
C0019522|T191|PT|0000006132|CHV|hidradenoma|8400/0
C0019522|T191|SY|0000006132|CHV|syringadenoma|8400/0
C0019522|T191|MH|D006607|MSH|Adenoma, Sweat Gland|8400/0
C0019522|T191|PM|D006607|MSH|Adenomas, Sweat Gland|8400/0
C0019522|T191|PM|D006607|MSH|Sweat Gland Adenoma|8400/0
C0019522|T191|PM|D006607|MSH|Sweat Gland Adenomas|8400/0
C0019522|T191|ET|D006607|MSH|Syringadenoma|8400/0
C0019522|T191|PM|D006607|MSH|Syringadenomas|8400/0
C0019522|T191|PN|NOCODE|MTH|Adenoma, Sweat Gland|8400/0
C0019522|T191|SY|C7563|NCI|Acrospiroma|8400/0
C0019522|T191|SY|C7560|NCI|Adenoma of Sweat Gland|8400/0
C0019522|T191|SY|C7560|NCI|Adenoma of the Sweat Gland|8400/0
C0019522|T191|SY|C7563|NCI|Eccrine Acrospiroma|8400/0
C0019522|T191|PT|C7563|NCI|Hidradenoma|8400/0
C0019522|T191|PT|C7560|NCI|Sweat Gland Adenoma|8400/0
C0019522|T191|SY|C7560|NCI_CDISC|Adenoma of Sweat Gland|8400/0
C0019522|T191|SY|C7560|NCI_CDISC|Adenoma of the Sweat Gland|8400/0
C0019522|T191|PT|C7560|NCI_CDISC|ADENOMA, SWEAT GLAND, BENIGN|8400/0
C0019522|T191|IS|X78Ss|RCD|Acrospiradenoma|8400/0
C0019522|T191|IS|X78Ss|RCD|Acrospiroma|8400/0
C0019522|T191|PT|X77nm|RCD|Hidradenoma|8400/0
C0019522|T191|PT|XaBA1|RCD|Hidradenoma morphology|8400/0
C0019522|T191|PT|XM1FJ|RCD|Sweat gland adenoma|8400/0
C0019522|T191|SY|X77nm|RCD|Syringadenoma|8400/0
C0019522|T191|IS|X78Ss|RCD|Syringadenoma|8400/0
C0019522|T191|OP|X78ob|RCD|Syringoadenoma|8400/0
C0019522|T191|SY|XaBA1|RCDSY|Sweat gland adenoma|8400/0
C0019522|T191|OAS|254719003|SNOMEDCT_US|Acrospiradenoma|8400/0
C0019522|T191|SY|400099008|SNOMEDCT_US|Acrospiradenoma|8400/0
C0019522|T191|OAS|254719003|SNOMEDCT_US|Acrospiroma|8400/0
C0019522|T191|SY|400099008|SNOMEDCT_US|Acrospiroma|8400/0
C0019522|T191|PT|253020008|SNOMEDCT_US|Hidradenoma|8400/0
C0019522|T191|SY|81393009|SNOMEDCT_US|Hidradenoma|8400/0
C0019522|T191|OF|307574003|SNOMEDCT_US|Hidradenoma morphology|8400/0
C0019522|T191|OAP|189664001|SNOMEDCT_US|Hidradenoma morphology|8400/0
C0019522|T191|OAP|307574003|SNOMEDCT_US|Hidradenoma morphology|8400/0
C0019522|T191|OF|189664001|SNOMEDCT_US|Hidradenoma morphology|8400/0
C0019522|T191|SY|253020008|SNOMEDCT_US|Hidradenoma of skin|8400/0
C0019522|T191|IS|81393009|SNOMEDCT_US|Hidradenoma, NOS|8400/0
C0019522|T191|PT|81393009|SNOMEDCT_US|Sweat gland adenoma|8400/0
C0019522|T191|OAS|254719003|SNOMEDCT_US|Syringadenoma|8400/0
C0019522|T191|SY|81393009|SNOMEDCT_US|Syringadenoma|8400/0
C0019522|T191|SY|253020008|SNOMEDCT_US|Syringadenoma|8400/0
C0019522|T191|IS|81393009|SNOMEDCT_US|Syringadenoma, NOS|8400/0
C0019522|T191|OAS|189051001|SNOMEDCT_US|Syringoadenoma|8400/0
C0019522|T191|OAP|255182002|SNOMEDCT_US|Syringoadenoma|8400/0
C0038987|T191|SY|0000011950|CHV|gland neoplasm sweat|8400/1
C0038987|T191|SY|0000011950|CHV|gland sweat neoplasms|8400/1
C0038987|T191|SY|0000011950|CHV|gland sweat tumor|8400/1
C0038987|T191|SY|0000011950|CHV|gland sweat tumors|8400/1
C0038987|T191|PT|0000011950|CHV|sweat gland tumor|8400/1
C0038987|T191|SY|0000011950|CHV|sweat gland tumour|8400/1
C0038987|T191|MTH_PT|10042658|MDR|Sweat gland tumor|8400/1
C0038987|T191|LLT|10042657|MDR|Sweat gland tumor|8400/1
C0038987|T191|MTH_LLT|10042659|MDR|Sweat gland tumor NOS|8400/1
C0038987|T191|LLT|10042658|MDR|Sweat gland tumour|8400/1
C0038987|T191|PT|10042658|MDR|Sweat gland tumour|8400/1
C0038987|T191|LLT|10042659|MDR|Sweat gland tumour NOS|8400/1
C0038987|T191|SY|354927|MEDCIN|neoplasm of integumentary system sweat gland|8400/1
C0038987|T191|PT|354927|MEDCIN|Neoplasm of sweat gland|8400/1
C0038987|T191|DEV|D013544|MSH|NEOPL SWEAT GLAND|8400/1
C0038987|T191|PM|D013544|MSH|Neoplasm, Sweat Gland|8400/1
C0038987|T191|ET|D013544|MSH|Neoplasms, Sweat Gland|8400/1
C0038987|T191|DEV|D013544|MSH|SWEAT GLAND NEOPL|8400/1
C0038987|T191|PM|D013544|MSH|Sweat Gland Neoplasm|8400/1
C0038987|T191|MH|D013544|MSH|Sweat Gland Neoplasms|8400/1
C0038987|T191|SY|C3398|NCI|Neoplasm of Sweat Gland|8400/1
C0038987|T191|SY|C3398|NCI|Neoplasm of the Sweat Gland|8400/1
C0038987|T191|PT|C3398|NCI|Sweat Gland Neoplasm|8400/1
C0038987|T191|SY|C3398|NCI|Sweat Gland Neoplasms|8400/1
C0038987|T191|SY|C3398|NCI|Sweat Gland Tumor|8400/1
C0038987|T191|SY|C3398|NCI|Tumor of Sweat Gland|8400/1
C0038987|T191|SY|C3398|NCI|Tumor of the Sweat Gland|8400/1
C0038987|T191|PT|Xa98g|RCD|Sweat gland tumour|8400/1
C0038987|T191|PT|X78Sc|RCD|Tumour of skin with eccrine differentiation|8400/1
C0038987|T191|AB|X78Sc|RCD|Tumour skin with eccrine diffn|8400/1
C0038987|T191|PT|Xa98g|RCDAE|Sweat gland tumor|8400/1
C0038987|T191|PT|X78Sc|RCDAE|Tumor of skin with eccrine differentiation|8400/1
C0038987|T191|AB|X78Sc|RCDAE|Tumor skin with eccrine diffn|8400/1
C0038987|T191|OP|BB611|RCDSA|Sweat gland tumor NOS|8400/1
C0038987|T191|OP|BB611|RCDSY|Sweat gland tumour NOS|8400/1
C0038987|T191|PT|126490003|SNOMEDCT_US|Neoplasm of sweat gland|8400/1
C0038987|T191|PT|12933008|SNOMEDCT_US|Sweat gland tumor|8400/1
C0038987|T191|IS|12933008|SNOMEDCT_US|Sweat gland tumor, NOS|8400/1
C0038987|T191|PTGB|12933008|SNOMEDCT_US|Sweat gland tumour|8400/1
C0038987|T191|SY|126490003|SNOMEDCT_US|Tumor of skin with eccrine differentiation|8400/1
C0038987|T191|SYGB|126490003|SNOMEDCT_US|Tumour of skin with eccrine differentiation|8400/1
C0334344|T191|SY|0000029960|CHV|digital papillary adenocarcinoma|8400/3
C0334344|T191|SY|0000029960|CHV|hidradenocarcinoma|8400/3
C0334344|T191|SY|0000029960|CHV|malignant nodular hidradenoma|8400/3
C0334344|T191|PT|0000029960|CHV|sweat gland carcinoma|8400/3
C0334344|T191|PT|10073088|MDR|Hidradenocarcinoma|8400/3
C0334344|T191|LLT|10073088|MDR|Hidradenocarcinoma|8400/3
C0334344|T191|PT|231626|MEDCIN|adenocarcinoma of sweat gland|8400/3
C0334344|T191|PN|NOCODE|MTH|Sweat gland adenocarcinoma|8400/3
C1412016|T191|PN|NOCODE|MTH|Sweat gland carcinoma|8400/3
C1412016|T191|SY|C6938|NCI|Carcinoma of Sweat Gland|8400/3
C1412016|T191|SY|C6938|NCI|Carcinoma of the Sweat Gland|8400/3
C0334344|T191|SY|C54664|NCI|Clear Cell Eccrine Carcinoma|8400/3
C0334344|T191|PT|C54664|NCI|Hidradenocarcinoma|8400/3
C1412016|T191|PT|C6938|NCI|Sweat Gland Carcinoma|8400/3
C1412016|T191|SY|C6938|NCI_CDISC|Carcinoma of Sweat Gland|8400/3
C1412016|T191|SY|C6938|NCI_CDISC|Carcinoma of the Sweat Gland|8400/3
C1412016|T191|PT|C6938|NCI_CDISC|CARCINOMA, SWEAT GLAND, MALIGNANT|8400/3
C0334344|T191|SY|X78Se|RCD|Hidradenocarcinoma|8400/3
C0334344|T191|SY|X78Sf|RCD|Hidradenocarcinoma|8400/3
C0334344|T191|PT|X78Sf|RCD|Sweat gland adenocarcinoma|8400/3
C1412016|T191|SY|X78Sd|RCD|Sweat gland carcinoma|8400/3
C1412016|T191|SY|X78Se|RCD|Sweat gland carcinoma|8400/3
C0334344|T191|OP|BB612|RCDSY|Sweat gland adenocarcinoma|8400/3
C0334344|T191|SY|254709009|SNOMEDCT_US|Hidradenocarcinoma|8400/3
C0334344|T191|SY|128894005|SNOMEDCT_US|Hidradenocarcinoma|8400/3
C0334344|T191|IS|254708001|SNOMEDCT_US|Hidradenocarcinoma|8400/3
C0334344|T191|PT|128894005|SNOMEDCT_US|Nodular hidradenoma, malignant|8400/3
C0334344|T191|SY|254709009|SNOMEDCT_US|Sweat gland adenocarcinoma|8400/3
C0334344|T191|OAP|254721008|SNOMEDCT_US|Sweat gland adenocarcinoma|8400/3
C0334344|T191|OF|254721008|SNOMEDCT_US|Sweat gland adenocarcinoma|8400/3
C0334344|T191|PT|32272007|SNOMEDCT_US|Sweat gland adenocarcinoma|8400/3
C1412016|T191|SY|254707006|SNOMEDCT_US|Sweat gland carcinoma|8400/3
C1412016|T191|SY|32272007|SNOMEDCT_US|Sweat gland carcinoma|8400/3
C1412016|T191|IS|254708001|SNOMEDCT_US|Sweat gland carcinoma|8400/3
C0334345|T191|SY|0000029961|CHV|adenoma apocrine|8401/0
C0334345|T191|SY|0000029961|CHV|apocrine cystadenoma|8401/0
C0334345|T191|PT|0000029961|CHV|apocrine hidrocystoma|8401/0
C0334345|T191|LLT|10072669|MDR|Tubular apocrine adenoma|8401/0
C0334345|T191|PN|NOCODE|MTH|Apocrine adenoma|8401/0
C0334345|T191|PT|C4168|NCI|Apocrine Adenoma|8401/0
C0334345|T191|PT|C27527|NCI|Tubular Apocrine Adenoma|8401/0
C0334345|T191|PT|XaBAq|RCD|Apocrine adenoma|8401/0
C0334345|T191|SY|XaBAq|RCD|Tubular apocrine adenoma|8401/0
C0334345|T191|PT|BB620|RCDSY|Apocrine adenoma|8401/0
C0334345|T191|PT|307596009|SNOMEDCT_US|Apocrine adenoma|8401/0
C0334345|T191|PT|36318001|SNOMEDCT_US|Apocrine adenoma|8401/0
C0334345|T191|SY|307596009|SNOMEDCT_US|Tubular apocrine adenoma|8401/0
C0334346|T191|PT|MTHU003370|ICPC2ICD10ENG|adenocarcinoma; apocrine, unspecified site|8401/3
C0334346|T191|PT|MTHU007557|ICPC2ICD10ENG|apocrine; adenocarcinoma, unspecified site|8401/3
C0334346|T191|PT|271480|MEDCIN|apocrine adenocarcinoma|8401/3
C1706827|T191|PT|C4169|NCI|Apocrine Carcinoma|8401/3
C1706827|T191|SY|C4169|NCI|Apocrine Gland Carcinoma|8401/3
C1706827|T191|SY|C4169|NCI|Carcinoma of Apocrine Gland|8401/3
C0334346|T191|PT|BB621|RCD|Apocrine adenocarcinoma|8401/3
C0334346|T191|PT|57141000|SNOMEDCT_US|Apocrine adenocarcinoma|8401/3
C0206671|T191|SY|0000021009|CHV|clear cell hidradenoma|8402/0
C0206671|T191|SY|0000021009|CHV|eccrine acrospiroma|8402/0
C0206671|T191|PT|0000021009|CHV|nodular hidradenoma|8402/0
C1370701|T191|PT|MTHU016916|ICPC2ICD10ENG|clear cell; hidradenoma|8402/0
C1370701|T191|PT|MTHU035117|ICPC2ICD10ENG|hidradenoma; clear cell|8402/0
C0206671|T191|PEP|D018250|MSH|Acrospiroma, Eccrine|8402/0
C0206671|T191|ET|D018250|MSH|Eccrine Acrospiroma|8402/0
C0206671|T191|PM|D018250|MSH|Eccrine Acrospiromas|8402/0
C0206671|T191|ET|D018250|MSH|Eccrine Spiradenoma|8402/0
C0206671|T191|PM|D018250|MSH|Eccrine Spiradenomas|8402/0
C0206671|T191|PM|D018250|MSH|Spiradenoma, Eccrine|8402/0
C0206671|T191|PM|D018250|MSH|Spiradenomas, Eccrine|8402/0
C1370701|T191|PN|NOCODE|MTH|Clear cell hidradenoma|8402/0
C0206671|T191|PN|NOCODE|MTH|Eccrine acrospiroma|8402/0
C1370701|T191|PT|C7567|NCI|Clear Cell Hidradenoma|8402/0
C0206671|T191|PT|C7568|NCI|Nodular Hidradenoma|8402/0
C0206671|T191|SY|C7568|NCI|Solid and Cystic Hidradenoma|8402/0
C0206671|T191|IS|X78Ss|RCD|Apocrine nodular hidradenoma|8402/0
C1370701|T191|IS|X78Ss|RCD|Clear cell hidradenoma|8402/0
C1370701|T191|IS|X78Ss|RCD|Clear cell myoepithelioma|8402/0
C1370701|T191|IS|X78Ss|RCD|Clear cell sweat gland adenoma|8402/0
C0206671|T191|IS|X78Ss|RCD|Eccrine acrospiroma|8402/0
C0206671|T191|OP|X78Ss|RCD|Eccrine hidradenoma|8402/0
C0206671|T191|IS|X78Ss|RCD|Eccrine nodular hidradenoma|8402/0
C0206671|T191|IS|X78Ss|RCD|Nodular apocrine hidradenoma|8402/0
C0206671|T191|SY|X77nm|RCD|Nodular hidradenoma|8402/0
C0206671|T191|IS|X78Ss|RCD|Nodular hidradenoma|8402/0
C0206671|T191|IS|X78Ss|RCD|Solid - cystic hidradenoma|8402/0
C0206671|T191|IS|X78Ss|RCD|Solid-cystic hidradenoma|8402/0
C1370701|T191|SY|BB63.|RCDSY|Clear cell hidradenoma|8402/0
C0206671|T191|PT|BB63.|RCDSY|Eccrine acrospiroma|8402/0
C0206671|T191|OAS|254719003|SNOMEDCT_US|Apocrine nodular hidradenoma|8402/0
C0206671|T191|SY|400099008|SNOMEDCT_US|Apocrine nodular hidradenoma|8402/0
C1370701|T191|OAS|254719003|SNOMEDCT_US|Clear cell hidradenoma|8402/0
C1370701|T191|PT|81143000|SNOMEDCT_US|Clear cell hidradenoma|8402/0
C1370701|T191|SY|400099008|SNOMEDCT_US|Clear cell hidradenoma|8402/0
C1370701|T191|OAS|254719003|SNOMEDCT_US|Clear cell myoepithelioma|8402/0
C1370701|T191|SY|400099008|SNOMEDCT_US|Clear cell myoepithelioma|8402/0
C1370701|T191|OAS|254719003|SNOMEDCT_US|Clear cell sweat gland adenoma|8402/0
C1370701|T191|SY|400099008|SNOMEDCT_US|Clear cell sweat gland adenoma|8402/0
C0206671|T191|OAS|254719003|SNOMEDCT_US|Eccrine acrospiroma|8402/0
C0206671|T191|SY|400099008|SNOMEDCT_US|Eccrine acrospiroma|8402/0
C0206671|T191|SY|81143000|SNOMEDCT_US|Eccrine acrospiroma|8402/0
C0206671|T191|OAP|254719003|SNOMEDCT_US|Eccrine hidradenoma|8402/0
C0206671|T191|PT|400099008|SNOMEDCT_US|Eccrine hidradenoma|8402/0
C0206671|T191|SY|400099008|SNOMEDCT_US|Eccrine hidradenoma of skin|8402/0
C0206671|T191|SY|400099008|SNOMEDCT_US|Eccrine nodular hidradenoma|8402/0
C0206671|T191|OAS|254719003|SNOMEDCT_US|Eccrine nodular hidradenoma|8402/0
C0206671|T191|OAS|254719003|SNOMEDCT_US|Nodular apocrine hidradenoma|8402/0
C0206671|T191|OAS|254719003|SNOMEDCT_US|Nodular hidradenoma|8402/0
C0206671|T191|SY|81143000|SNOMEDCT_US|Nodular hidradenoma|8402/0
C0206671|T191|SY|253020008|SNOMEDCT_US|Nodular hidradenoma|8402/0
C0206671|T191|IS|400099008|SNOMEDCT_US|Nodular hidradenoma|8402/0
C0206671|T191|IS|81393009|SNOMEDCT_US|Nodular hidradenoma|8402/0
C0206671|T191|OAS|254719003|SNOMEDCT_US|Solid-cystic hidradenoma|8402/0
C0206671|T191|SY|400099008|SNOMEDCT_US|Solid-cystic hidradenoma|8402/0
C0334344|T191|SY|0000029960|CHV|digital papillary adenocarcinoma|8402/3
C0334344|T191|SY|0000029960|CHV|hidradenocarcinoma|8402/3
C0334344|T191|SY|0000029960|CHV|malignant nodular hidradenoma|8402/3
C0334344|T191|PT|0000029960|CHV|sweat gland carcinoma|8402/3
C0334344|T191|PT|10073088|MDR|Hidradenocarcinoma|8402/3
C0334344|T191|LLT|10073088|MDR|Hidradenocarcinoma|8402/3
C0334344|T191|PT|231626|MEDCIN|adenocarcinoma of sweat gland|8402/3
C1275213|T191|PT|357597|MEDCIN|Clear cell eccrine hidradenocarcinoma of skin|8402/3
C1260964|T191|PT|357595|MEDCIN|Eccrine ductal carcinoma of skin|8402/3
C1275213|T191|SY|357597|MEDCIN|skin neop malign adnexa w/ eccrine differentiation clear cell hidradenocarcinoma|8402/3
C1260964|T191|SY|357595|MEDCIN|skin neoplasm malignant adnexa with eccrine differentiation ductal carcinoma|8402/3
C0334344|T191|PN|NOCODE|MTH|Sweat gland adenocarcinoma|8402/3
C0334344|T191|SY|C54664|NCI|Clear Cell Eccrine Carcinoma|8402/3
C1260964|T191|PT|C43345|NCI|Ductal Eccrine Adenocarcinoma|8402/3
C1260964|T191|SY|C43345|NCI|Ductal Eccrine Carcinoma|8402/3
C0334344|T191|PT|C54664|NCI|Hidradenocarcinoma|8402/3
C0334344|T191|SY|X78Se|RCD|Hidradenocarcinoma|8402/3
C0334344|T191|SY|X78Sf|RCD|Hidradenocarcinoma|8402/3
C0334344|T191|PT|X78Sf|RCD|Sweat gland adenocarcinoma|8402/3
C0334344|T191|OP|BB612|RCDSY|Sweat gland adenocarcinoma|8402/3
C1260964|T191|SY|403939009|SNOMEDCT_US|Anaplastic syringoma|8402/3
C1275213|T191|PT|403940006|SNOMEDCT_US|Clear cell eccrine hidradenocarcinoma|8402/3
C1275213|T191|PT|400147009|SNOMEDCT_US|Clear cell eccrine hidradenocarcinoma|8402/3
C1275213|T191|SY|403940006|SNOMEDCT_US|Clear cell eccrine hidradenocarcinoma of skin|8402/3
C1260964|T191|PT|400208002|SNOMEDCT_US|Eccrine ductal carcinoma|8402/3
C1260964|T191|PT|403939009|SNOMEDCT_US|Eccrine ductal carcinoma|8402/3
C1260964|T191|SY|403939009|SNOMEDCT_US|Eccrine ductal carcinoma of skin|8402/3
C0334344|T191|IS|254708001|SNOMEDCT_US|Hidradenocarcinoma|8402/3
C0334344|T191|SY|254709009|SNOMEDCT_US|Hidradenocarcinoma|8402/3
C0334344|T191|SY|128894005|SNOMEDCT_US|Hidradenocarcinoma|8402/3
C1260964|T191|SY|403939009|SNOMEDCT_US|Malignant acrospiroma|8402/3
C1260964|T191|SY|403939009|SNOMEDCT_US|Malignant eccrine acrospiroma|8402/3
C0334344|T191|PT|128894005|SNOMEDCT_US|Nodular hidradenoma, malignant|8402/3
C0334344|T191|OAP|254721008|SNOMEDCT_US|Sweat gland adenocarcinoma|8402/3
C0334344|T191|OF|254721008|SNOMEDCT_US|Sweat gland adenocarcinoma|8402/3
C0334344|T191|PT|32272007|SNOMEDCT_US|Sweat gland adenocarcinoma|8402/3
C0334344|T191|SY|254709009|SNOMEDCT_US|Sweat gland adenocarcinoma|8402/3
C0334347|T191|SY|0000029962|CHV|eccrine spiradenoma|8403/0
C0334347|T191|PT|0000029962|CHV|spiradenoma|8403/0
C0334347|T191|LLT|10065278|MDR|Eccrine spiradenoma|8403/0
C0334347|T191|PN|NOCODE|MTH|Eccrine spiradenoma|8403/0
C0334347|T191|SY|C4170|NCI|Benign Eccrine Spiradenoma|8403/0
C0334347|T191|SY|C4170|NCI|Eccrine Spiradenoma|8403/0
C0334347|T191|PT|C4170|NCI|Spiradenoma|8403/0
C0334347|T191|PT|BB64.|RCD|Eccrine spiradenoma|8403/0
C0334347|T191|SY|BB64.|RCD|Spiradenoma|8403/0
C0334347|T191|PT|4977000|SNOMEDCT_US|Eccrine spiradenoma|8403/0
C0334347|T191|PT|403938001|SNOMEDCT_US|Eccrine spiradenoma|8403/0
C0334347|T191|SY|403938001|SNOMEDCT_US|Eccrine spiradenoma of skin|8403/0
C0334347|T191|SY|4977000|SNOMEDCT_US|Spiradenoma|8403/0
C0334347|T191|SY|403938001|SNOMEDCT_US|Spiradenoma|8403/0
C0334347|T191|SY|403938001|SNOMEDCT_US|Spiradenoma eccrine|8403/0
C0334347|T191|IS|4977000|SNOMEDCT_US|Spiradenoma, NOS|8403/0
C1266063|T191|PT|231629|MEDCIN|malignant eccrine spiradenoma of skin|8403/3
C1266063|T191|SY|C5117|NCI|Malignant Eccrine Spiradenoma|8403/3
C1266063|T191|SY|C5117|NCI|Malignant Spiradenoma|8403/3
C1266063|T191|PT|C5117|NCI|Spiradenocarcinoma|8403/3
C1266063|T191|PT|403942003|SNOMEDCT_US|Malignant eccrine spiradenoma|8403/3
C1266063|T191|PT|128895006|SNOMEDCT_US|Malignant eccrine spiradenoma|8403/3
C1266063|T191|SY|403942003|SNOMEDCT_US|Malignant eccrine spiradenoma of skin|8403/3
C1266063|T191|SY|403942003|SNOMEDCT_US|Malignant spiradenoma|8403/3
C0206672|T191|SY|0000021010|CHV|eccrine hidrocystoma|8404/0
C0206672|T191|PT|0000021010|CHV|hidrocystoma|8404/0
C0206672|T191|LLT|10059019|MDR|Hidrocystoma|8404/0
C0206672|T191|MH|D018251|MSH|Hidrocystoma|8404/0
C0206672|T191|PM|D018251|MSH|Hidrocystomas|8404/0
C0206672|T191|PN|NOCODE|MTH|Hidrocystoma|8404/0
C0206672|T191|PT|C3760|NCI|Hidrocystoma|8404/0
C0206672|T191|SY|C3760|NCI|Hydrocystoma|8404/0
C0206672|T191|PT|BB65.|RCD|Hidrocystoma|8404/0
C0206672|T191|PT|80549000|SNOMEDCT_US|Hidrocystoma|8404/0
C0334348|T191|SY|0000029963|CHV|hidradenoma papilliferum|8405/0
C0334348|T191|SY|0000029963|CHV|hydradenomas papillary|8405/0
C0334348|T191|PT|0000029963|CHV|papillary hidradenoma|8405/0
C0334348|T191|PT|MTHU035118|ICPC2ICD10ENG|hidradenoma; papillary|8405/0
C0334348|T191|PT|MTHU057308|ICPC2ICD10ENG|papillary; hidradenoma|8405/0
C0334348|T191|LLT|10020042|MDR|Hidradenoma papilliferum|8405/0
C0334348|T191|ET|D000074009|MSH|Anogenital Papillary Hidradenoma|8405/0
C0334348|T191|PM|D000074009|MSH|Anogenital Papillary Hidradenomas|8405/0
C0334348|T191|PEP|D000074009|MSH|Hidradenoma Papilliferum|8405/0
C0334348|T191|PM|D000074009|MSH|Hidradenoma Papilliferums|8405/0
C0334348|T191|PM|D000074009|MSH|Hidradenoma, Anogenital Papillary|8405/0
C0334348|T191|PM|D000074009|MSH|Hidradenoma, Papillary|8405/0
C0334348|T191|ET|D000074009|MSH|Papillary Hidradenoma|8405/0
C0334348|T191|PM|D000074009|MSH|Papillary Hidradenoma, Anogenital|8405/0
C0334348|T191|PM|D000074009|MSH|Papillary Hidradenomas|8405/0
C0334348|T191|PM|D000074009|MSH|Papilliferum, Hidradenoma|8405/0
C0334348|T191|SY|C4171|NCI|Hidradenoma Papilliferum|8405/0
C0334348|T191|PT|C4171|NCI|Papillary Hidradenoma|8405/0
C0334348|T191|SY|XaBAr|RCD|Hidradenoma papilliferum|8405/0
C0334348|T191|PT|XaBAr|RCD|Papillary hidradenoma|8405/0
C0334348|T191|PT|BB66.|RCDSY|Papillary hydradenoma|8405/0
C0334348|T191|SY|89791006|SNOMEDCT_US|Hidradenoma papilliferum|8405/0
C0334348|T191|SY|307597000|SNOMEDCT_US|Hidradenoma papilliferum|8405/0
C0334348|T191|PT|89791006|SNOMEDCT_US|Papillary hidradenoma|8405/0
C0334348|T191|PT|307597000|SNOMEDCT_US|Papillary hidradenoma|8405/0
C0406803|T191|PT|MTHU057310|ICPC2ICD10ENG|papillary; syringadenoma|8406/0
C0406803|T191|PT|MTHU057311|ICPC2ICD10ENG|papillary; syringocystadenoma|8406/0
C0406803|T191|PT|MTHU073160|ICPC2ICD10ENG|syringadenoma; papillary|8406/0
C0406803|T191|PT|MTHU073168|ICPC2ICD10ENG|syringocystadenoma; papillary|8406/0
C0406803|T191|LLT|10042926|MDR|Syringocystadenoma papilliferum|8406/0
C0406803|T191|ET|D000074009|MSH|Papillary Syringocystadenoma|8406/0
C0406803|T191|PM|D000074009|MSH|Papillary Syringocystadenomas|8406/0
C0406803|T191|PM|D000074009|MSH|Papilliferum, Syringocystadenoma|8406/0
C0406803|T191|PEP|D000074009|MSH|Syringocystadenoma Papilliferum|8406/0
C0406803|T191|PM|D000074009|MSH|Syringocystadenoma Papilliferums|8406/0
C0406803|T191|PM|D000074009|MSH|Syringocystadenoma, Papillary|8406/0
C0406803|T191|PN|NOCODE|MTH|Syringocystadenoma Papilliferum|8406/0
C0406803|T191|SY|C4172|NCI|Papillary Syringadenoma|8406/0
C0406803|T191|SY|C4172|NCI|Papillary Syringocystadenoma|8406/0
C0406803|T191|SY|C4172|NCI|Syringadenoma|8406/0
C0406803|T191|PT|C4172|NCI|Syringocystadenoma Papilliferum|8406/0
C0406803|T191|AB|X50Jf|RCD|Naev syringocystadeno papillif|8406/0
C0406803|T191|SY|X50Jf|RCD|Naevus syringocystadenomatosus papilliferus|8406/0
C0406803|T191|PT|BB67.|RCD|Papillary syringadenoma|8406/0
C0406803|T191|SY|BB67.|RCD|Papillary syringocystadenoma|8406/0
C0406803|T191|AB|X50Jf|RCD|Syringocystadenoma papillif|8406/0
C0406803|T191|PT|X50Jf|RCD|Syringocystadenoma papilliferum|8406/0
C0406803|T191|SY|X50Jf|RCDAE|Nevus syringocystadenomatosus papilliferus|8406/0
C0406803|T191|SYGB|239121009|SNOMEDCT_US|Naevus syringocystadenomatosus papilliferus|8406/0
C0406803|T191|SY|239121009|SNOMEDCT_US|Nevus syringocystadenomatosus papilliferus|8406/0
C0406803|T191|PT|8934006|SNOMEDCT_US|Papillary syringadenoma|8406/0
C0406803|T191|SY|8934006|SNOMEDCT_US|Papillary syringocystadenoma|8406/0
C3697936|T191|PT|733887006|SNOMEDCT_US|Sialadenoma papilliferum|8406/0
C3697936|T191|PT|699277009|SNOMEDCT_US|Sialadenoma papilliferum|8406/0
C0406803|T191|PT|239121009|SNOMEDCT_US|Syringocystadenoma papilliferum|8406/0
C0406803|T191|SY|8934006|SNOMEDCT_US|Syringocystadenoma papilliferum|8406/0
C0206673|T191|PT|0000021011|CHV|syringoma|8407/0
C0206673|T191|SY|0000021011|CHV|syringomas|8407/0
C0206673|T191|DI|U001809|DXP|SYRINGOMA|8407/0
C0206673|T191|LLT|10042927|MDR|Syringoma|8407/0
C0206673|T191|SY|275523|MEDCIN|benign syringoma|8407/0
C0206673|T191|PT|275523|MEDCIN|syringoma of skin|8407/0
C0206673|T191|MH|D018252|MSH|Syringoma|8407/0
C0206673|T191|PM|D018252|MSH|Syringomas|8407/0
C0206673|T191|SY|C3761|NCI|Eccrine Syringoma|8407/0
C0206673|T191|PT|C3761|NCI|Syringoma|8407/0
C0431093|T191|PT|Xa0By|RCD|Clear cell syringoma|8407/0
C0206673|T191|PT|Xa98h|RCD|Syringoma|8407/0
C0206673|T191|PT|BB68.|RCDSY|Syringoma NOS|8407/0
C0431093|T191|PT|403934004|SNOMEDCT_US|Clear cell syringoma|8407/0
C0431093|T191|PT|276736008|SNOMEDCT_US|Clear cell syringoma|8407/0
C3839745|T191|SY|703552001|SNOMEDCT_US|Infiltrating syringomatous adenoma of nipple|8407/0
C0206673|T191|PT|71244007|SNOMEDCT_US|Syringoma|8407/0
C0206673|T191|PT|302828001|SNOMEDCT_US|Syringoma|8407/0
C0206673|T191|OAS|189051001|SNOMEDCT_US|Syringoma|8407/0
C0206673|T191|SY|302828001|SNOMEDCT_US|Syringoma of skin|8407/0
C0206673|T191|IS|71244007|SNOMEDCT_US|Syringoma, NOS|8407/0
C3839745|T191|SY|703552001|SNOMEDCT_US|Syringomatous adenoma of nipple|8407/0
C3839745|T191|PT|703552001|SNOMEDCT_US|Syringomatous tumor of nipple|8407/0
C3839745|T191|PTGB|703552001|SNOMEDCT_US|Syringomatous tumour of nipple|8407/0
C0346027|T191|SY|0000031042|CHV|carcinomas syringomatous|8407/3
C0346027|T191|PT|0000031042|CHV|microcystic adnexal carcinoma|8407/3
C0346027|T191|LLT|10073091|MDR|Microcystic adnexal carcinoma|8407/3
C0346027|T191|PT|231630|MEDCIN|sclerosing carcinoma of sweat duct|8407/3
C0346027|T191|SY|231630|MEDCIN|sclerosing sweat duct carcinoma|8407/3
C0346027|T191|NM|C000632664|MSH|Microcystic adnexal carcinoma|8407/3
C0346027|T191|SY|C7581|NCI|Eccrine Epithelioma|8407/3
C0346027|T191|PT|C7581|NCI|Microcystic Adnexal Carcinoma|8407/3
C0346027|T191|SY|C7581|NCI|Syringomatous Carcinoma|8407/3
C0346027|T191|PT|X78Sx|RCD|Eccrine epithelioma|8407/3
C0346027|T191|SY|X78Si|RCD|Malignant syringoma|8407/3
C0346027|T191|PT|X78Si|RCD|Microcystic adnexal carcinoma|8407/3
C0346027|T191|AB|X78Si|RCD|Sclerosing sweat duct carcinom|8407/3
C0346027|T191|SY|X78Si|RCD|Sclerosing sweat duct carcinoma|8407/3
C0346027|T191|SY|X78Si|RCD|Syringoid eccrine carcinoma|8407/3
C0346027|T191|AB|X78Si|RCD|Syringomat sweat duct carcinom|8407/3
C0346027|T191|SY|X78Si|RCD|Syringomatous sweat duct carcinoma|8407/3
C0346027|T191|PT|400135003|SNOMEDCT_US|Eccrine epithelioma|8407/3
C0346027|T191|PT|254722001|SNOMEDCT_US|Eccrine epithelioma|8407/3
C0346027|T191|SY|254722001|SNOMEDCT_US|Eccrine epithelioma of skin|8407/3
C0346027|T191|SY|254712007|SNOMEDCT_US|Malignant syringoma|8407/3
C0346027|T191|PT|254712007|SNOMEDCT_US|Microcystic adnexal carcinoma|8407/3
C0346027|T191|SY|128896007|SNOMEDCT_US|Microcystic adnexal carcinoma|8407/3
C0346027|T191|SY|254712007|SNOMEDCT_US|Microcystic adnexal carcinoma of skin|8407/3
C0346027|T191|PT|128896007|SNOMEDCT_US|Sclerosing sweat duct carcinoma|8407/3
C0346027|T191|SY|254712007|SNOMEDCT_US|Sclerosing sweat duct carcinoma|8407/3
C0346027|T191|SY|254712007|SNOMEDCT_US|Syringoid eccrine carcinoma|8407/3
C0346027|T191|SY|128896007|SNOMEDCT_US|Syringomatous carcinoma|8407/3
C0346027|T191|SY|254712007|SNOMEDCT_US|Syringomatous sweat duct carcinoma|8407/3
C0334350|T191|OP|C4173|NCI|Eccrine Papillary Adenoma|8408/0
C0334350|T191|OP|C4173|NCI|Papillary Eccrine Adenoma|8408/0
C0334350|T191|PT|C4173|NCI|Papillary Eccrine Adenoma|8408/0
C0334350|T191|AB|XaBA2|RCD|Eccrine papillary adenom morph|8408/0
C0334350|T191|PT|X77nn|RCD|Eccrine papillary adenoma|8408/0
C0334350|T191|PT|XaBA2|RCD|Eccrine papillary adenoma morphology|8408/0
C0334350|T191|OP|BB6B.|RCDSY|Eccrine papillary adenoma|8408/0
C0334350|T191|PT|253021007|SNOMEDCT_US|Eccrine papillary adenoma|8408/0
C0334350|T191|PT|10060008|SNOMEDCT_US|Eccrine papillary adenoma|8408/0
C0334350|T191|OAP|134345002|SNOMEDCT_US|Eccrine papillary adenoma morphology|8408/0
C0334350|T191|SY|253021007|SNOMEDCT_US|Eccrine papillary adenoma of skin|8408/0
C1367789|T191|LLT|10079286|MDR|Digital papillary carcinoma|8408/1
C1367789|T191|PN|NOCODE|MTH|Digital papillary eccrine carcinoma of skin|8408/1
C1367789|T191|PT|C27534|NCI|Aggressive Digital Papillary Adenocarcinoma|8408/1
C1266064|T191|PT|C162848|NCI|Aggressive Digital Papillary Adenoma|8408/1
C1367789|T191|SY|C27534|NCI|Digital Papillary Carcinoma|8408/1
C1367789|T191|CSN|C27534|NCI|Digital Papillary Eccrine Carcinoma|8408/1
C1367789|T191|SY|C27534|NCI|Papillary Digital Eccrine Carcinoma|8408/1
C1367789|T191|AB|X78Sf|RCD|Papill digit eccrine carcinom|8408/1
C1367789|T191|SY|X78Sf|RCD|Papillary digital eccrine carcinoma|8408/1
C1266064|T191|PT|128897003|SNOMEDCT_US|Aggressive digital papillary adenoma|8408/1
C1367789|T191|SY|254709009|SNOMEDCT_US|Digital papillary adenocarcinoma|8408/1
C1367789|T191|PT|254709009|SNOMEDCT_US|Digital papillary eccrine carcinoma of skin|8408/1
C1367789|T191|SY|254709009|SNOMEDCT_US|Papillary digital eccrine carcinoma|8408/1
C1367789|T191|LLT|10079286|MDR|Digital papillary carcinoma|8408/3
C1367789|T191|PN|NOCODE|MTH|Digital papillary eccrine carcinoma of skin|8408/3
C1367774|T191|PN|NOCODE|MTH|Eccrine Papillary Adenocarcinoma|8408/3
C1367789|T191|PT|C27534|NCI|Aggressive Digital Papillary Adenocarcinoma|8408/3
C1367789|T191|SY|C27534|NCI|Digital Papillary Carcinoma|8408/3
C1367789|T191|CSN|C27534|NCI|Digital Papillary Eccrine Carcinoma|8408/3
C1367789|T191|SY|C27534|NCI|Papillary Digital Eccrine Carcinoma|8408/3
C1367789|T191|AB|X78Sf|RCD|Papill digit eccrine carcinom|8408/3
C1367789|T191|SY|X78Sf|RCD|Papillary digital eccrine carcinoma|8408/3
C1367774|T191|SY|128898008|SNOMEDCT_US|Digital papillary adenocarcinoma|8408/3
C1367789|T191|SY|254709009|SNOMEDCT_US|Digital papillary adenocarcinoma|8408/3
C1367789|T191|PT|254709009|SNOMEDCT_US|Digital papillary eccrine carcinoma of skin|8408/3
C1367774|T191|PT|128898008|SNOMEDCT_US|Eccrine papillary adenocarcinoma|8408/3
C1367789|T191|SY|254709009|SNOMEDCT_US|Papillary digital eccrine carcinoma|8408/3
C1533161|T191|PT|0000058008|CHV|eccrine poroma|8409/0
C1533161|T191|LLT|10014083|MDR|Eccrine poroma|8409/0
C1533161|T191|PEP|D057091|MSH|Eccrine Poroma|8409/0
C1533161|T191|PM|D057091|MSH|Eccrine Poromas|8409/0
C1533161|T191|PM|D057091|MSH|Poroma, Eccrine|8409/0
C1533161|T191|PN|NOCODE|MTH|Eccrine Poroma|8409/0
C1533161|T191|SY|C27273|NCI|Eccrine Poroma|8409/0
C1533161|T191|PT|C27273|NCI|Poroma|8409/0
C1533161|T191|IS|X78Ss|RCD|Eccrine poroma|8409/0
C1533161|T191|SY|BB63.|RCDSY|Eccrine poroma|8409/0
C1533161|T191|OAS|254719003|SNOMEDCT_US|Eccrine poroma|8409/0
C1533161|T191|PT|399985004|SNOMEDCT_US|Eccrine poroma|8409/0
C1533161|T191|PT|128915006|SNOMEDCT_US|Eccrine poroma|8409/0
C1533161|T191|IS|81143000|SNOMEDCT_US|Eccrine poroma|8409/0
C1533161|T191|SY|399985004|SNOMEDCT_US|Eccrine poroma of skin|8409/0
C1266065|T191|SY|0000056681|CHV|malignant eccrine poroma|8409/3
C1266065|T191|PT|0000056681|CHV|porocarcinoma|8409/3
C1266065|T191|LLT|10063609|MDR|Porocarcinoma|8409/3
C1266065|T191|PT|10063609|MDR|Porocarcinoma|8409/3
C1266065|T191|PT|357599|MEDCIN|Eccrine porocarcinoma of skin|8409/3
C1266065|T191|SY|357599|MEDCIN|skin neop malignant adnexa w/ eccrine differentiation porocarcinoma|8409/3
C1266065|T191|MH|D057090|MSH|Eccrine Porocarcinoma|8409/3
C1266065|T191|PM|D057090|MSH|Eccrine Porocarcinomas|8409/3
C1266065|T191|PM|D057090|MSH|Eccrine Poroma, Malignant|8409/3
C1266065|T191|PM|D057090|MSH|Eccrine Poromas, Malignant|8409/3
C1266065|T191|ET|D057090|MSH|Malignant Eccrine Poroma|8409/3
C1266065|T191|PM|D057090|MSH|Malignant Eccrine Poromas|8409/3
C1266065|T191|PM|D057090|MSH|Porocarcinoma, Eccrine|8409/3
C1266065|T191|PM|D057090|MSH|Porocarcinomas, Eccrine|8409/3
C1266065|T191|PM|D057090|MSH|Poroma, Malignant Eccrine|8409/3
C1266065|T191|PM|D057090|MSH|Poromas, Malignant Eccrine|8409/3
C1266065|T191|PN|NOCODE|MTH|Eccrine porocarcinoma|8409/3
C1266065|T191|PT|C5560|NCI|Eccrine Porocarcinoma|8409/3
C1266065|T191|SY|C5560|NCI|Epidermotropic Eccrine Carcinoma|8409/3
C1266065|T191|SY|C5560|NCI|Malignant Eccrine Poroma|8409/3
C1266065|T191|PT|X78Se|RCD|Eccrine porocarcinoma|8409/3
C1266065|T191|PT|254708001|SNOMEDCT_US|Eccrine porocarcinoma|8409/3
C1266065|T191|SY|254708001|SNOMEDCT_US|Eccrine porocarcinoma of skin|8409/3
C1266065|T191|PT|128685001|SNOMEDCT_US|Eccrine poroma, malignant|8409/3
C1266065|T191|SY|128685001|SNOMEDCT_US|Porocarcinoma|8409/3
C1368816|T191|PT|0000030021|CHV|sebaceous adenoma|8410/0
C1368816|T191|SY|HP:0009720|HPO|Sebaceous adenoma|8410/0
C1368816|T191|ET|HP:0009720|HPO|Sebaceous adenomas|8410/0
C1368816|T191|LLT|10062919|MDR|Sebaceous adenoma|8410/0
C1368816|T191|PT|10062919|MDR|Sebaceous adenoma|8410/0
C1368816|T191|PN|NOCODE|MTH|Sebaceous adenoma|8410/0
C1368816|T191|SY|C4174|NCI|Adenoma of Sebaceous Gland|8410/0
C1368816|T191|SY|C4174|NCI|Adenoma of the Sebaceous Gland|8410/0
C1368816|T191|PT|C4174|NCI|Sebaceous Adenoma|8410/0
C1368816|T191|SY|C4174|NCI|Sebaceous Gland Adenoma|8410/0
C1368816|T191|SY|C4174|NCI|Skin Appendage Sebaceous Adenoma|8410/0
C1368816|T191|SY|C4174|NCI_CDISC|Adenoma of Sebaceous Gland|8410/0
C1368816|T191|SY|C4174|NCI_CDISC|Adenoma of the Sebaceous Gland|8410/0
C1368816|T191|SY|C4174|NCI_CDISC|Adenoma, Sebaceous Cell|8410/0
C1368816|T191|PT|C4174|NCI_CDISC|ADENOMA, SEBACEOUS, BENIGN|8410/0
C1368816|T191|SY|C4174|NCI_CDISC|Sebaceous Gland Adenoma|8410/0
C1368816|T191|SY|C4174|NCI_CDISC|Skin Appendage Sebaceous Adenoma|8410/0
C1368816|T191|SY|BB690|RCD|Sebaceous adenoma|8410/0
C4518353|T191|PT|734049008|SNOMEDCT_US|Cystic sebaceous neoplasm|8410/0
C4518557|T191|PT|733036009|SNOMEDCT_US|Non-sebaceous lymphadenoma|8410/0
C1368816|T191|PT|78424008|SNOMEDCT_US|Sebaceous adenoma|8410/0
C4518582|T191|PT|733102000|SNOMEDCT_US|Sebaceous lymphadenoma|8410/0
C0206684|T191|SY|0000021018|CHV|adenocarcinoma sebaceous|8410/3
C0206684|T191|PT|0000021018|CHV|sebaceous carcinoma|8410/3
C0206684|T191|SY|0000021018|CHV|sebaceous gland carcinoma|8410/3
C0206684|T191|SY|HP:0030410|HPO|Sebaceous carcinoma|8410/3
C0206684|T191|PT|HP:0030410|HPO|Sebaceous gland carcinoma|8410/3
C0206684|T191|LLT|10068784|MDR|Sebaceous carcinoma|8410/3
C0206684|T191|PT|10068784|MDR|Sebaceous carcinoma|8410/3
C0206684|T191|SY|356679|MEDCIN|malignant sebaceous adenocarcinoma|8410/3
C0206684|T191|PT|356679|MEDCIN|sebaceous adenocarcinoma|8410/3
C0206684|T191|MH|D018266|MSH|Adenocarcinoma, Sebaceous|8410/3
C0206684|T191|PM|D018266|MSH|Adenocarcinomas, Sebaceous|8410/3
C0206684|T191|PM|D018266|MSH|Sebaceous Adenocarcinoma|8410/3
C0206684|T191|PM|D018266|MSH|Sebaceous Adenocarcinomas|8410/3
C0206684|T191|PN|NOCODE|MTH|Sebaceous Adenocarcinoma|8410/3
C0206684|T191|SY|C40310|NCI|Carcinoma of Sebaceous Gland|8410/3
C0206684|T191|SY|C40310|NCI|Carcinoma of the Sebaceous Gland|8410/3
C0206684|T191|PT|C40310|NCI|Sebaceous Carcinoma|8410/3
C0206684|T191|SY|C40310|NCI|Sebaceous Gland Carcinoma|8410/3
C0206684|T191|PT|C40310|NCI_CDISC|ADENOCARCINOMA, SEBACEOUS, MALIGNANT|8410/3
C0206684|T191|SY|C40310|NCI_CDISC|Carcinoma of Sebaceous Gland|8410/3
C0206684|T191|SY|C40310|NCI_CDISC|Carcinoma of the Sebaceous Gland|8410/3
C0206684|T191|SY|C40310|NCI_CDISC|Carcinoma, Sebaceous Cell|8410/3
C0206684|T191|SY|C40310|NCI_CDISC|Sebaceous Gland Carcinoma|8410/3
C0206684|T191|DN|C40310|NCI_CTRP|Sebaceous Cancer|8410/3
C0206684|T191|SY|CDR0000636561|PDQ|Carcinoma of Sebaceous Gland|8410/3
C0206684|T191|SY|CDR0000636561|PDQ|Carcinoma of the Sebaceous Gland|8410/3
C0206684|T191|SY|CDR0000636561|PDQ|Sebaceous Carcinoma|8410/3
C0206684|T191|PT|CDR0000636561|PDQ|sebaceous gland carcinoma|8410/3
C0206684|T191|SY|XaBAt|RCD|Carcinoma of sebaceous gland|8410/3
C0206684|T191|PT|XaBAt|RCD|Sebaceous adenocarcinoma|8410/3
C0206684|T191|SY|XaBAt|RCD|Sebaceous carcinoma|8410/3
C0206684|T191|PT|BB691|RCDSY|Sebaceous adenocarcinoma|8410/3
C0206684|T191|SY|307599002|SNOMEDCT_US|Carcinoma of sebaceous gland|8410/3
C0206684|T191|PT|54734006|SNOMEDCT_US|Sebaceous adenocarcinoma|8410/3
C0206684|T191|PT|307599002|SNOMEDCT_US|Sebaceous adenocarcinoma|8410/3
C0206684|T191|SY|54734006|SNOMEDCT_US|Sebaceous carcinoma|8410/3
C0206684|T191|SY|307599002|SNOMEDCT_US|Sebaceous carcinoma|8410/3
C4518359|T191|PT|734055003|SNOMEDCT_US|Sebaceous lymphadenocarcinoma|8410/3
C1302864|T191|LLT|10069680|MDR|Eccrine carcinoma|8413/3
C1302864|T191|PT|10069680|MDR|Eccrine carcinoma|8413/3
C1302864|T191|PT|357594|MEDCIN|Eccrine carcinoma of skin|8413/3
C1302864|T191|SY|357594|MEDCIN|skin neoplasm malignant adnexa with eccrine differentiation carcinoma|8413/3
C1302864|T191|PT|C27255|NCI|Eccrine Carcinoma|8413/3
C1302864|T191|PT|C27255|NCI_CDISC|CARCINOMA, ECCRINE GLAND, MALIGNANT|8413/3
C1302864|T191|DN|C27255|NCI_CTRP|Eccrine Carcinoma|8413/3
C1302864|T191|SY|CDR0000559689|PDQ|Eccrine Carcinoma|8413/3
C1302864|T191|PT|CDR0000559689|PDQ|eccrine carcinoma of the skin|8413/3
C1266066|T191|PT|128686000|SNOMEDCT_US|Eccrine adenocarcinoma|8413/3
C1302864|T191|PT|400173004|SNOMEDCT_US|Eccrine carcinoma of skin|8413/3
C0334352|T191|SY|HP:0040097|HPO|Adenoma of the ceruminous gland|8420/0
C0334352|T191|SY|HP:0040097|HPO|Ceruminoma|8420/0
C0334352|T191|SY|HP:0040097|HPO|Ceruminous adenoma|8420/0
C0334352|T191|PT|HP:0040097|HPO|Neoplasm of the ceruminal gland|8420/0
C0334352|T191|PT|MTHU003486|ICPC2ICD10ENG|adenoma; ceruminous|8420/0
C0334352|T191|PT|MTHU015732|ICPC2ICD10ENG|ceruminous; adenoma|8420/0
C0334352|T191|PN|NOCODE|MTH|Ceruminous adenoma|8420/0
C1333488|T191|PN|NOCODE|MTH|External Auditory Canal Ceruminous Adenoma|8420/0
C1333488|T191|SY|C6088|NCI|Ceruminoma|8420/0
C1333488|T191|SY|C6088|NCI|Ceruminous Adenoma|8420/0
C1333488|T191|SY|C6088|NCI|Ceruminous Adenoma of External Auditory Canal|8420/0
C1333488|T191|SY|C6088|NCI|Ceruminous Adenoma of the External Auditory Canal|8420/0
C1333488|T191|PT|C6088|NCI|External Auditory Canal Ceruminous Adenoma|8420/0
C1333488|T191|PT|C6088|NCI_CDISC|ADENOMA, CERUMINOUS GLAND, BENIGN|8420/0
C1333488|T191|SY|C6088|NCI_CDISC|Ceruminoma|8420/0
C1333488|T191|SY|C6088|NCI_CDISC|Ceruminous Adenoma|8420/0
C1333488|T191|SY|C6088|NCI_CDISC|Ceruminous Adenoma of External Auditory Canal|8420/0
C1333488|T191|SY|C6088|NCI_CDISC|Ceruminous Adenoma of the External Auditory Canal|8420/0
C0334352|T191|PT|BB6A0|RCD|Ceruminous adenoma|8420/0
C0334352|T191|PT|403945001|SNOMEDCT_US|Ceruminous adenoma|8420/0
C0334352|T191|PT|52707009|SNOMEDCT_US|Ceruminous adenoma|8420/0
C0334353|T191|PT|MTHU003374|ICPC2ICD10ENG|adenocarcinoma; ceruminous|8420/3
C0334353|T191|PT|MTHU014734|ICPC2ICD10ENG|carcinoma; ceruminous|8420/3
C0334353|T191|PT|MTHU015731|ICPC2ICD10ENG|ceruminous; adenocarcinoma|8420/3
C0334353|T191|PT|MTHU015733|ICPC2ICD10ENG|ceruminous; carcinoma|8420/3
C0334353|T191|PT|C4176|NCI|Ceruminous Adenocarcinoma|8420/3
C0334353|T191|PT|C4176|NCI_CDISC|CARCINOMA, CERUMINOUS GLAND, MALIGNANT|8420/3
C0334353|T191|PT|BB6A1|RCD|Ceruminous adenocarcinoma|8420/3
C0334353|T191|SY|BB6A1|RCD|Ceruminous carcinoma|8420/3
C0334353|T191|PT|58069009|SNOMEDCT_US|Ceruminous adenocarcinoma|8420/3
C0334353|T191|SY|58069009|SNOMEDCT_US|Ceruminous carcinoma|8420/3
C0206694|T191|PT|0000021026|CHV|mucoepidermoid carcinoma|8430/1
C0206694|T191|LLT|10057269|MDR|Mucoepidermoid carcinoma|8430/1
C0206694|T191|PT|10057269|MDR|Mucoepidermoid carcinoma|8430/1
C0206694|T191|PT|271429|MEDCIN|mucoepidermoid carcinoma|8430/1
C0206694|T191|MH|D018277|MSH|Carcinoma, Mucoepidermoid|8430/1
C0206694|T191|PM|D018277|MSH|Carcinomas, Mucoepidermoid|8430/1
C0206694|T191|PM|D018277|MSH|Mucoepidermoid Carcinoma|8430/1
C0206694|T191|PM|D018277|MSH|Mucoepidermoid Carcinomas|8430/1
C0206712|T191|MH|D018298|MSH|Mucoepidermoid Tumor|8430/1
C0206712|T191|PM|D018298|MSH|Mucoepidermoid Tumors|8430/1
C0206712|T191|PM|D018298|MSH|Tumor, Mucoepidermoid|8430/1
C0206712|T191|PM|D018298|MSH|Tumors, Mucoepidermoid|8430/1
C0206694|T191|PN|NOCODE|MTH|Mucoepidermoid Carcinoma|8430/1
C0206694|T191|AB|C3772|NCI|MEC|8430/1
C0206694|T191|SY|TCGA|NCI|Mucoepidermoid Carcinoma|8430/1
C0206694|T191|PT|C3772|NCI|Mucoepidermoid Carcinoma|8430/1
C0206694|T191|PT|BB71.|RCD|Mucoepidermoid carcinoma|8430/1
C0206712|T191|PT|BB70.|RCD|Mucoepidermoid tumour|8430/1
C0206712|T191|PT|BB70.|RCDAE|Mucoepidermoid tumor|8430/1
C0206712|T191|OP|BB7z.|RCDSY|Mucoepidermoid neoplasm NOS|8430/1
C0206712|T191|OP|BB7..|RCDSY|Mucoepidermoid neoplasms|8430/1
C0206694|T191|PT|4079000|SNOMEDCT_US|Mucoepidermoid carcinoma|8430/1
C0206712|T191|SY|127571003|SNOMEDCT_US|Mucoepidermoid neoplasm|8430/1
C0206712|T191|OP|39892006|SNOMEDCT_US|Mucoepidermoid tumor|8430/1
C0206712|T191|PT|39892006|SNOMEDCT_US|Mucoepidermoid tumor uncertain whether benign or malignant|8430/1
C0206712|T191|IS|39892006|SNOMEDCT_US|Mucoepidermoid tumor, uncertain whether benign or malignant|8430/1
C0206712|T191|OP|39892006|SNOMEDCT_US|Mucoepidermoid tumour|8430/1
C0206712|T191|PTGB|39892006|SNOMEDCT_US|Mucoepidermoid tumour uncertain whether benign or malignant|8430/1
C0206712|T191|IS|39892006|SNOMEDCT_US|Mucoepidermoid tumour, uncertain whether benign or malignant|8430/1
C0206694|T191|PT|0000021026|CHV|mucoepidermoid carcinoma|8430/3
C0206694|T191|LLT|10057269|MDR|Mucoepidermoid carcinoma|8430/3
C0206694|T191|PT|10057269|MDR|Mucoepidermoid carcinoma|8430/3
C0206694|T191|PT|271429|MEDCIN|mucoepidermoid carcinoma|8430/3
C0206694|T191|MH|D018277|MSH|Carcinoma, Mucoepidermoid|8430/3
C0206694|T191|PM|D018277|MSH|Carcinomas, Mucoepidermoid|8430/3
C0206694|T191|PM|D018277|MSH|Mucoepidermoid Carcinoma|8430/3
C0206694|T191|PM|D018277|MSH|Mucoepidermoid Carcinomas|8430/3
C0206694|T191|PN|NOCODE|MTH|Mucoepidermoid Carcinoma|8430/3
C0206694|T191|AB|C3772|NCI|MEC|8430/3
C0206694|T191|SY|TCGA|NCI|Mucoepidermoid Carcinoma|8430/3
C0206694|T191|PT|C3772|NCI|Mucoepidermoid Carcinoma|8430/3
C0206694|T191|PT|BB71.|RCD|Mucoepidermoid carcinoma|8430/3
C0206694|T191|PT|4079000|SNOMEDCT_US|Mucoepidermoid carcinoma|8430/3
C1301193|T191|PT|397081004|SNOMEDCT_US|Mucoepidermoid carcinoma, high grade|8430/3
C1301192|T191|PT|397080003|SNOMEDCT_US|Mucoepidermoid carcinoma, intermediate grade|8430/3
C1301191|T191|PT|397079001|SNOMEDCT_US|Mucoepidermoid carcinoma, low grade|8430/3
C5231078|T191|PT|822964002|SNOMEDCT_US|Sclerosing mucoepidermoid carcinoma with eosinophilia|8430/3
C5231078|T191|SY|822964002|SNOMEDCT_US|SMECE - sclerosing mucoepidermoid carcinoma with eosinophilia|8430/3
C0010633|T191|PT|1017483|CCPSS|CYSTADENOMA|8440/0
C0010633|T191|PT|0000003542|CHV|cystadenoma|8440/0
C0010633|T191|SY|0000003542|CHV|cystadenomas|8440/0
C0010633|T191|SY|0000003542|CHV|cystoma|8440/0
C0010633|T191|LLT|10011812|MDR|Cystoma|8440/0
C0010633|T191|MH|D003537|MSH|Cystadenoma|8440/0
C0010633|T191|PM|D003537|MSH|Cystadenomas|8440/0
C0010633|T191|PN|NOCODE|MTH|Cystadenoma|8440/0
C0010633|T191|PT|C2972|NCI|Cystadenoma|8440/0
C0010633|T191|SY|C2972|NCI|Cystoma|8440/0
C0010633|T191|PT|C2972|NCI_CDISC|CYSTADENOMA, BENIGN|8440/0
C0010633|T191|SY|C2972|NCI_CDISC|Cystoma|8440/0
C0010633|T191|PT|Xa98j|RCD|Cystadenoma|8440/0
C0010633|T191|SY|Xa98j|RCD|Cystoma|8440/0
C0010633|T191|SY|Xa98j|RCDSY|Cystadenoma NOS|8440/0
C0010633|T191|OAP|189680006|SNOMEDCT_US|Cystadenoma|8440/0
C0010633|T191|OF|189680006|SNOMEDCT_US|Cystadenoma|8440/0
C0010633|T191|PT|47620003|SNOMEDCT_US|Cystadenoma|8440/0
C0010633|T191|IS|47620003|SNOMEDCT_US|Cystadenoma, NOS|8440/0
C0010633|T191|SY|47620003|SNOMEDCT_US|Cystoma|8440/0
C0010633|T191|IS|47620003|SNOMEDCT_US|Cystoma, NOS|8440/0
C0010631|T191|PT|0000003541|CHV|cystadenocarcinoma|8440/3
C0010631|T191|SY|0000003541|CHV|cystadenocarcinomas|8440/3
C0010631|T191|LLT|10063387|MDR|Cystadenocarcinoma|8440/3
C0010631|T191|PT|271439|MEDCIN|cystadenocarcinoma|8440/3
C0010631|T191|MH|D003536|MSH|Cystadenocarcinoma|8440/3
C0010631|T191|PM|D003536|MSH|Cystadenocarcinomas|8440/3
C0010631|T191|PT|C2971|NCI|Cystadenocarcinoma|8440/3
C0010631|T191|SY|TCGA|NCI|Cystadenocarcinoma|8440/3
C0010631|T191|PT|C2971|NCI_CDISC|CYSTADENOCARCINOMA, MALIGNANT|8440/3
C0010631|T191|PT|Xa98k|RCD|Cystadenocarcinoma|8440/3
C0010631|T191|OP|BB801|RCDSY|Cystadenocarcinoma NOS|8440/3
C0010631|T191|PT|21008007|SNOMEDCT_US|Cystadenocarcinoma|8440/3
C0010631|T191|IS|21008007|SNOMEDCT_US|Cystadenocarcinoma, NOS|8440/3
C2960605|T191|PT|447011009|SNOMEDCT_US|Mixed serous and mucinous cystadenocarcinoma|8440/3
C0206709|T191|PT|0037527|CCPSS|CYSTADENOMA SEROUS|8441/0
C0206709|T191|SY|0000021038|CHV|cystadenoma serous|8441/0
C0206709|T191|PT|0000021038|CHV|serous cystadenoma|8441/0
C0206709|T191|SY|0000021038|CHV|serous cystoma|8441/0
C0206709|T191|PT|MTHU020860|ICPC2ICD10ENG|cystoma; serous, unspecified site|8441/0
C0206709|T191|PT|MTHU067559|ICPC2ICD10ENG|serous; cystoma, unspecified site|8441/0
C0206709|T191|MH|D018293|MSH|Cystadenoma, Serous|8441/0
C0206709|T191|PM|D018293|MSH|Cystadenomas, Serous|8441/0
C0206709|T191|PM|D018293|MSH|Serous Cystadenoma|8441/0
C0206709|T191|PM|D018293|MSH|Serous Cystadenomas|8441/0
C0206709|T191|PT|C3783|NCI|Serous Cystadenoma|8441/0
C0206709|T191|SY|C3783|NCI|Serous Cystoma|8441/0
C0206709|T191|PT|Xa98l|RCD|Serous cystadenoma|8441/0
C0206709|T191|SY|Xa98l|RCD|Serous cystoma|8441/0
C0206709|T191|OP|BB810|RCDSY|Serous cystadenoma NOS|8441/0
C0206709|T191|PT|51608009|SNOMEDCT_US|Serous cystadenoma|8441/0
C0206709|T191|IS|51608009|SNOMEDCT_US|Serous cystadenoma, NOS|8441/0
C0206709|T191|SY|51608009|SNOMEDCT_US|Serous cystoma|8441/0
C0206709|T191|SY|51608009|SNOMEDCT_US|Serous microcystic adenoma|8441/0
C3838709|T191|PT|703558002|SNOMEDCT_US|Serous intraepithelial carcinoma|8441/2
C0206701|T191|SY|0000021032|CHV|serous adenocarcinoma|8441/3
C0206701|T191|PT|0000021032|CHV|serous carcinoma|8441/3
C0206701|T191|SY|0000021032|CHV|serous cystadenocarcinoma|8441/3
C0206701|T191|MH|D018284|MSH|Cystadenocarcinoma, Serous|8441/3
C0206701|T191|PM|D018284|MSH|Cystadenocarcinomas, Serous|8441/3
C0206701|T191|PM|D018284|MSH|Serous Cystadenocarcinoma|8441/3
C0206701|T191|PM|D018284|MSH|Serous Cystadenocarcinomas|8441/3
C0206701|T191|PN|NOCODE|MTH|Serous Cystadenocarcinoma|8441/3
C0206701|T191|SY|C3778|NCI|Serous Adenocarcinoma|8441/3
C0206701|T191|PT|C40101|NCI|Serous Adenocarcinoma|8441/3
C0206701|T191|PT|C3778|NCI|Serous Cystadenocarcinoma|8441/3
C0206701|T191|SY|TCGA|NCI|Serous Cystadenocarcinoma|8441/3
C0206701|T191|SY|Xa98m|RCD|Serous adenocarcinoma|8441/3
C0206701|T191|PT|Xa98m|RCD|Serous cystadenocarcinoma|8441/3
C0206701|T191|OA|BB812|RCDSY|Serous cystadenocarcin.NOS|8441/3
C0206701|T191|OP|BB812|RCDSY|Serous cystadenocarcinoma, NOS|8441/3
C0206701|T191|SY|90725004|SNOMEDCT_US|Papillary serous adenocarcinoma|8441/3
C0206701|T191|SY|90725004|SNOMEDCT_US|Papillary serous cystadenocarcinoma|8441/3
C0206701|T191|SY|90725004|SNOMEDCT_US|Serous adenocarcinoma|8441/3
C0206701|T191|IS|90725004|SNOMEDCT_US|Serous adenocarcinoma, NOS|8441/3
C0206701|T191|SY|90725004|SNOMEDCT_US|Serous carcinoma|8441/3
C0206701|T191|PT|90725004|SNOMEDCT_US|Serous cystadenocarcinoma|8441/3
C0206701|T191|IS|90725004|SNOMEDCT_US|Serous cystadenocarcinoma, NOS|8441/3
C0206701|T191|SY|90725004|SNOMEDCT_US|Serous surface papillary carcinoma|8441/3
C0334355|T191|PN|NOCODE|MTH|Serous cystadenoma, borderline malignancy|8442/1
C0334355|T191|SY|C4177|NCI|Borderline Malignancy Serous Cystadenoma|8442/1
C0334355|T191|PT|C4177|NCI|Borderline Serous Cystadenoma|8442/1
C0334355|T191|SY|C4177|NCI|Low Malignancy Potential Serous Cystadenoma|8442/1
C0334355|T191|SY|C4177|NCI|Serous Tumor of Borderline Malignant Potential|8442/1
C0334355|T191|PT|BB811|RCD|Serous cystadenoma - borderline malignancy|8442/1
C0334355|T191|AB|BB811|RCD|Serous cystadenoma-bord malign|8442/1
C0334355|T191|AB|BB811|RCD|Serous tumour low malig potent|8442/1
C0334355|T191|SY|BB811|RCD|Serous tumour of low malignant potential|8442/1
C0334355|T191|AB|BB811|RCDAE|Serous tumor low malig potent|8442/1
C0334355|T191|SY|BB811|RCDAE|Serous tumor of low malignant potential|8442/1
C0334355|T191|AB|BB811|RCDSY|Ser cystaden, borderl malig|8442/1
C0334355|T191|SY|BB811|RCDSY|Serous cystadenoma, borderline malignancy|8442/1
C0334355|T191|SY|128849004|SNOMEDCT_US|Atypical proliferating serous tumor|8442/1
C0334355|T191|SYGB|128849004|SNOMEDCT_US|Atypical proliferating serous tumour|8442/1
C0334355|T191|SY|128849004|SNOMEDCT_US|Serous borderline tumor|8442/1
C0334355|T191|SYGB|128849004|SNOMEDCT_US|Serous borderline tumour|8442/1
C0334355|T191|OAP|189694007|SNOMEDCT_US|Serous cystadenoma - borderline malignancy|8442/1
C0334355|T191|OF|189694007|SNOMEDCT_US|Serous cystadenoma - borderline malignancy|8442/1
C0334355|T191|OAP|37529007|SNOMEDCT_US|Serous cystadenoma, borderline malignancy|8442/1
C0334355|T191|PT|128849004|SNOMEDCT_US|Serous cystadenoma, borderline malignancy|8442/1
C0334355|T191|IS|37529007|SNOMEDCT_US|Serous cystadenoma, borderline malignancy -RETIRED-|8442/1
C0334355|T191|OF|37529007|SNOMEDCT_US|Serous cystadenoma, borderline malignancy -RETIRED-|8442/1
C0334355|T191|SY|128849004|SNOMEDCT_US|Serous tumor of low malignant potential|8442/1
C0334355|T191|SY|128849004|SNOMEDCT_US|Serous tumor, atypical proliferative|8442/1
C0334355|T191|IS|37529007|SNOMEDCT_US|Serous tumor, NOS, of low malignant potential|8442/1
C0334355|T191|SYGB|128849004|SNOMEDCT_US|Serous tumour of low malignant potential|8442/1
C0334355|T191|SYGB|128849004|SNOMEDCT_US|Serous tumour, atypical proliferative|8442/1
C1880102|T191|PT|C65203|NCI|Clear Cell Papillary Cystadenoma|8443/0
C1266068|T191|PT|128687009|SNOMEDCT_US|Clear cell cystadenoma|8443/0
C1511260|T191|PT|C40083|NCI|Borderline Ovarian Clear Cell Cystadenofibroma|8444/1
C1266069|T191|SY|128688004|SNOMEDCT_US|Atypical proliferating clear cell tumor|8444/1
C1266069|T191|SYGB|128688004|SNOMEDCT_US|Atypical proliferating clear cell tumour|8444/1
C1266069|T191|PT|128688004|SNOMEDCT_US|Clear cell cystic tumor of borderline malignancy|8444/1
C1266069|T191|PTGB|128688004|SNOMEDCT_US|Clear cell cystic tumour of borderline malignancy|8444/1
C0010636|T191|PT|0000003544|CHV|papillary cystadenoma|8450/0
C0010636|T191|PT|MTHU020321|ICPC2ICD10ENG|cystadenoma; papillary, unspecified site|8450/0
C0010636|T191|PT|MTHU057299|ICPC2ICD10ENG|papillary; cystadenoma, unspecified site|8450/0
C0010636|T191|MH|D018292|MSH|Cystadenoma, Papillary|8450/0
C0010636|T191|PM|D018292|MSH|Cystadenomas, Papillary|8450/0
C0010636|T191|PM|D018292|MSH|Papillary Cystadenoma|8450/0
C0010636|T191|PM|D018292|MSH|Papillary Cystadenomas|8450/0
C0010636|T191|PT|C2974|NCI|Papillary Cystadenoma|8450/0
C0010636|T191|PT|C2974|NCI_CDISC|CYSTADENOMA, PAPILLARY, BENIGN|8450/0
C0010636|T191|PT|Xa98n|RCD|Papillary cystadenoma|8450/0
C0010636|T191|OP|BB813|RCDSY|Papillary cystadenoma NOS|8450/0
C0010636|T191|PT|32140001|SNOMEDCT_US|Papillary cystadenoma|8450/0
C0010636|T191|IS|32140001|SNOMEDCT_US|Papillary cystadenoma, NOS|8450/0
C0206700|T191|PT|MTHU020295|ICPC2ICD10ENG|cystadenocarcinoma; papillary, unspecified site|8450/3
C0206700|T191|PT|MTHU057290|ICPC2ICD10ENG|papillary; cystadenocarcinoma, unspecified site|8450/3
C0206700|T191|MH|D018283|MSH|Cystadenocarcinoma, Papillary|8450/3
C0206700|T191|PM|D018283|MSH|Cystadenocarcinomas, Papillary|8450/3
C0206700|T191|PM|D018283|MSH|Papillary Cystadenocarcinoma|8450/3
C0206700|T191|PM|D018283|MSH|Papillary Cystadenocarcinomas|8450/3
C0206700|T191|PT|C3777|NCI|Papillary Cystadenocarcinoma|8450/3
C0206700|T191|PT|C3777|NCI_CDISC|CYSTADENOCARCINOMA, PAPILLARY, MALIGNANT|8450/3
C0206700|T191|PT|Xa98o|RCD|Papillary cystadenocarcinoma|8450/3
C0206700|T191|SY|Xa98o|RCD|Papillocystic adenocarcinoma|8450/3
C0206700|T191|OA|BB815|RCDSY|Papillary cystadenoca. NOS|8450/3
C0206700|T191|OP|BB815|RCDSY|Papillary cystadenocarcinoma, NOS|8450/3
C0206700|T191|PT|2735009|SNOMEDCT_US|Papillary cystadenocarcinoma|8450/3
C0206700|T191|IS|2735009|SNOMEDCT_US|Papillary cystadenocarcinoma, NOS|8450/3
C0206700|T191|SY|2735009|SNOMEDCT_US|Papillocystic adenocarcinoma|8450/3
C0334356|T191|PT|MTHU012118|ICPC2ICD10ENG|borderline malignancy; papillary cystadenoma, unspecified site|8451/1
C0334356|T191|PT|MTHU020315|ICPC2ICD10ENG|cystadenoma; papillary, borderline malignancy, unspecified site|8451/1
C0334356|T191|PT|MTHU057293|ICPC2ICD10ENG|papillary; cystadenoma, borderline malignancy, unspecified site|8451/1
C0334356|T191|SY|C4178|NCI|Borderline Malignancy Papillary Cystadenoma|8451/1
C0334356|T191|PT|C4178|NCI|Borderline Papillary Cystadenoma|8451/1
C0334356|T191|SY|C4178|NCI|Low Malignancy Potential Papillary Cystadenoma|8451/1
C0334356|T191|AB|BB814|RCD|Papill cystadenoma-bord malign|8451/1
C0334356|T191|PT|BB814|RCD|Papillary cystadenoma - borderline malignancy|8451/1
C0334356|T191|SY|BB814|RCDSY|Papillary cystadenoma, borderline malignancy|8451/1
C0334356|T191|AB|BB814|RCDSY|Papl cystaden, bordrl malig|8451/1
C0334356|T191|OAP|189695008|SNOMEDCT_US|Papillary cystadenoma - borderline malignancy|8451/1
C0334356|T191|OF|189695008|SNOMEDCT_US|Papillary cystadenoma - borderline malignancy|8451/1
C0334356|T191|OAP|47741001|SNOMEDCT_US|Papillary cystadenoma, borderline malignancy|8451/1
C0334356|T191|PT|128850004|SNOMEDCT_US|Papillary cystadenoma, borderline malignancy|8451/1
C0334356|T191|IS|47741001|SNOMEDCT_US|Papillary cystadenoma, borderline malignancy -RETIRED-|8451/1
C0334356|T191|OF|47741001|SNOMEDCT_US|Papillary cystadenoma, borderline malignancy -RETIRED-|8451/1
C0334357|T191|PT|MTHU057312|ICPC2ICD10ENG|papillary; tumor, cystic|8452/1
C0334357|T191|PT|MTHU077127|ICPC2ICD10ENG|tumor; papillary cystic|8452/1
C1336030|T191|LLT|10069368|MDR|Solid pseudopapillary tumor of the pancreas|8452/1
C1336030|T191|MTH_PT|10069345|MDR|Solid pseudopapillary tumor of the pancreas|8452/1
C1336030|T191|LLT|10069345|MDR|Solid pseudopapillary tumour of the pancreas|8452/1
C1336030|T191|PT|10069345|MDR|Solid pseudopapillary tumour of the pancreas|8452/1
C1336030|T191|SY|38693|MEDCIN|solid pseudopapillary pancreatic neoplasm|8452/1
C1336030|T191|PT|38693|MEDCIN|solid pseudopapillary tumor of pancreas|8452/1
C1336030|T191|OP|C37212|NCI|Frantz Tumor|8452/1
C0334357|T191|PT|C4179|NCI|Papillary Cystic Neoplasm|8452/1
C0334357|T191|SY|C4179|NCI|Papillary Cystic Tumor|8452/1
C1336030|T191|PT|C37212|NCI|Solid Pseudopapillary Neoplasm of the Pancreas|8452/1
C1336030|T191|OP|C37212|NCI|Solid Pseudopapillary Tumor of the Pancreas|8452/1
C0334357|T191|PT|X77ns|RCD|Papillary cystic tumour|8452/1
C0334357|T191|PT|X77ns|RCDAE|Papillary cystic tumor|8452/1
C0334357|T191|OAP|189696009|SNOMEDCT_US|Papillary cystic tumor|8452/1
C0334357|T191|PT|27078002|SNOMEDCT_US|Papillary cystic tumor|8452/1
C0334357|T191|PTGB|27078002|SNOMEDCT_US|Papillary cystic tumour|8452/1
C0334357|T191|OAP|189696009|SNOMEDCT_US|Papillary cystic tumour|8452/1
C0334357|T191|OF|189696009|SNOMEDCT_US|Papillary cystic tumour|8452/1
C0334357|T191|SY|27078002|SNOMEDCT_US|Solid and cystic tumor|8452/1
C0334357|T191|SYGB|27078002|SNOMEDCT_US|Solid and cystic tumour|8452/1
C0334357|T191|SY|27078002|SNOMEDCT_US|Solid and papillary epithelial neoplasm|8452/1
C0334357|T191|SY|27078002|SNOMEDCT_US|Solid pseudopapillary tumor|8452/1
C0334357|T191|SYGB|27078002|SNOMEDCT_US|Solid pseudopapillary tumour|8452/1
C1336029|T191|PT|38725|MEDCIN|solid pseudopapillary carcinoma of pancreas|8452/3
C1336029|T191|OP|C5728|NCI|Pancreatic Solid Pseudopapillary Carcinoma|8452/3
C1336029|T191|OP|C5728|NCI|Solid Pseudopapillary Carcinoma of Pancreas|8452/3
C1336029|T191|OP|C5728|NCI|Solid Pseudopapillary Carcinoma of the Pancreas|8452/3
C1336029|T191|PT|C5728|NCI|Solid Pseudopapillary Carcinoma of the Pancreas|8452/3
C1336029|T191|SY|782697005|SNOMEDCT_US|Pancreatic solid pseudopapillary carcinoma|8452/3
C1266070|T191|PT|116061001|SNOMEDCT_US|Solid pseudopapillary carcinoma|8452/3
C1336029|T191|PT|782697005|SNOMEDCT_US|Solid pseudopapillary carcinoma of pancreas|8452/3
C1518868|T191|SY|38688|MEDCIN|intraductal pancreatic papillary mucinous adenoma|8453/0
C1518868|T191|PT|38688|MEDCIN|intraductal papillary-mucinous adenoma of pancreas|8453/0
C1335305|T191|PT|38692|MEDCIN|intraductal papillary-mucinous neoplasm of pancreas with moderate dysplasia|8453/0
C1335305|T191|SY|38692|MEDCIN|pancreatic intraductal papillary mucinous neoplasm with moderate dysplasia|8453/0
C1266071|T191|PN|NOCODE|MTH|Intraductal papillary-mucinous adenoma|8453/0
C1518868|T191|PN|NOCODE|MTH|Pancreatic Intraductal Papillary-Mucinous Adenoma|8453/0
C1335305|T191|SY|C5719|NCI|Intraductal Papillary-Mucinous Neoplasm of Pancreas with Moderate Dysplasia|8453/0
C1335305|T191|SY|C5719|NCI|Intraductal Papillary-Mucinous Neoplasm of the Pancreas with Moderate Dysplasia|8453/0
C1335305|T191|SY|C5719|NCI|Intraductal Papillary-Mucinous Tumor of Pancreas with Moderate Dysplasia|8453/0
C1335305|T191|SY|C5719|NCI|Intraductal Papillary-Mucinous Tumor of the Pancreas with Moderate Dysplasia|8453/0
C1335305|T191|OP|C5719|NCI|Pancreatic Borderline Intraductal Papillary-Mucinous Neoplasm|8453/0
C1335305|T191|SY|C5719|NCI|Pancreatic Intraductal Papillary Mucinous Neoplasm with Intermediate Grade Dysplasia|8453/0
C1518868|T191|SY|C41249|NCI|Pancreatic Intraductal Papillary Mucinous Neoplasm with Low Grade Dysplasia|8453/0
C1518868|T191|OP|C41249|NCI|Pancreatic Intraductal Papillary-Mucinous Adenoma|8453/0
C1335305|T191|PT|C5719|NCI|Pancreatic Intraductal Papillary-Mucinous Neoplasm with Intermediate Grade Dysplasia|8453/0
C1518868|T191|PT|C41249|NCI|Pancreatic Intraductal Papillary-Mucinous Neoplasm with Low Grade Dysplasia|8453/0
C1335305|T191|SY|C5719|NCI|Pancreatic Intraductal Papillary-Mucinous Neoplasm with Moderate Dysplasia|8453/0
C1335305|T191|SY|C5719|NCI|Pancreatic Intraductal Papillary-Mucinous Tumor with Moderate Dysplasia|8453/0
C1266071|T191|SY|128689007|SNOMEDCT_US|Benign intra-ductal papillary mucinous neoplasm|8453/0
C1518868|T191|PT|473418001|SNOMEDCT_US|Intraductal papillary mucinous adenoma of pancreas|8453/0
C1518868|T191|SY|473418001|SNOMEDCT_US|Intraductal papillary mucinous neoplasm with intermediate dysplasia of pancreas|8453/0
C1518868|T191|IS|473418001|SNOMEDCT_US|Intraductal papillary mucinous neoplasm with low grade dysplasia|8453/0
C1266071|T191|SY|128689007|SNOMEDCT_US|Intraductal papillary mucinous neoplasm with low grade dysplasia|8453/0
C1518868|T191|SY|473418001|SNOMEDCT_US|Intraductal papillary mucinous neoplasm with low grade dysplasia of pancreas|8453/0
C1266071|T191|SY|128689007|SNOMEDCT_US|Intraductal papillary mucinous neoplasm with moderate dysplasia|8453/0
C1518868|T191|SY|473418001|SNOMEDCT_US|Intraductal papillary mucinous neoplasm with moderate dysplasia of pancreas|8453/0
C1266071|T191|SY|128689007|SNOMEDCT_US|Intraductal papillary mucinous tumor with intermediate dysplasia|8453/0
C1266071|T191|SY|128689007|SNOMEDCT_US|Intraductal papillary mucinous tumor with low grade dysplasia|8453/0
C1266071|T191|SY|128689007|SNOMEDCT_US|Intraductal papillary mucinous tumor with moderate dysplasia|8453/0
C1266071|T191|SYGB|128689007|SNOMEDCT_US|Intraductal papillary mucinous tumour with intermediate dysplasia|8453/0
C1266071|T191|SYGB|128689007|SNOMEDCT_US|Intraductal papillary mucinous tumour with low grade dysplasia|8453/0
C1266071|T191|SYGB|128689007|SNOMEDCT_US|Intraductal papillary mucinous tumour with moderate dysplasia|8453/0
C1266071|T191|PT|128689007|SNOMEDCT_US|Intraductal papillary-mucinous adenoma|8453/0
C1335305|T191|PT|38692|MEDCIN|intraductal papillary-mucinous neoplasm of pancreas with moderate dysplasia|8453/1
C1335305|T191|SY|38692|MEDCIN|pancreatic intraductal papillary mucinous neoplasm with moderate dysplasia|8453/1
C1335305|T191|SY|C5719|NCI|Intraductal Papillary-Mucinous Neoplasm of Pancreas with Moderate Dysplasia|8453/1
C1335305|T191|SY|C5719|NCI|Intraductal Papillary-Mucinous Neoplasm of the Pancreas with Moderate Dysplasia|8453/1
C1335305|T191|SY|C5719|NCI|Intraductal Papillary-Mucinous Tumor of Pancreas with Moderate Dysplasia|8453/1
C1335305|T191|SY|C5719|NCI|Intraductal Papillary-Mucinous Tumor of the Pancreas with Moderate Dysplasia|8453/1
C1335305|T191|OP|C5719|NCI|Pancreatic Borderline Intraductal Papillary-Mucinous Neoplasm|8453/1
C1335305|T191|SY|C5719|NCI|Pancreatic Intraductal Papillary Mucinous Neoplasm with Intermediate Grade Dysplasia|8453/1
C1335305|T191|PT|C5719|NCI|Pancreatic Intraductal Papillary-Mucinous Neoplasm with Intermediate Grade Dysplasia|8453/1
C1335305|T191|SY|C5719|NCI|Pancreatic Intraductal Papillary-Mucinous Neoplasm with Moderate Dysplasia|8453/1
C1335305|T191|SY|C5719|NCI|Pancreatic Intraductal Papillary-Mucinous Tumor with Moderate Dysplasia|8453/1
C1266073|T191|PN|NOCODE|MTH|Intraductal papillary-mucinous carcinoma, non-invasive|8453/2
C1518873|T191|SY|C41251|NCI|Pancreatic Intraductal Papillary Mucinous Neoplasm with High Grade Dysplasia|8453/2
C1518873|T191|PT|C41251|NCI|Pancreatic Intraductal Papillary-Mucinous Neoplasm with High Grade Dysplasia|8453/2
C1518873|T191|OP|C41251|NCI|Pancreatic Non-Invasive Intraductal Papillary-Mucinous Carcinoma|8453/2
C1266073|T191|SY|128691004|SNOMEDCT_US|Intraductal papillary mucinous carcinoma in situ|8453/2
C1266073|T191|SY|128691004|SNOMEDCT_US|Intraductal papillary mucinous neoplasm with high grade dysplasia|8453/2
C1266073|T191|PT|128691004|SNOMEDCT_US|Intraductal papillary-mucinous carcinoma, non-invasive|8453/2
C1518871|T191|PT|38721|MEDCIN|intraductal papillary-mucinous carcinoma of the pancreas invasive|8453/3
C1518871|T191|SY|38721|MEDCIN|invasive intraductal papillary-mucinous carcinoma of pancreas|8453/3
C1518871|T191|SY|C5726|NCI|Pancreatic Intraductal Papillary Mucinous Neoplasm with an Associated Invasive Carcinoma|8453/3
C1518871|T191|PT|C5726|NCI|Pancreatic Intraductal Papillary-Mucinous Neoplasm with an Associated Invasive Carcinoma|8453/3
C1518871|T191|OP|C5726|NCI|Pancreatic Invasive Intraductal Papillary-Mucinous Carcinoma|8453/3
C1266074|T191|SY|128692006|SNOMEDCT_US|Intraductal papillary mucinous neoplasm with an associated invasive carcinoma|8453/3
C1266074|T191|PT|128692006|SNOMEDCT_US|Intraductal papillary-mucinous carcinoma, invasive|8453/3
C1518871|T191|PT|780821007|SNOMEDCT_US|Invasive intraductal papillary-mucinous carcinoma of pancreas|8453/3
C1266074|T191|SY|128692006|SNOMEDCT_US|Malignant intraductal papillary mucinous neoplasm|8453/3
C1266074|T191|SY|128692006|SNOMEDCT_US|Malignant intraductal papillary mucinous neoplasm with an associated invasive carcinoma|8453/3
C1518871|T191|SY|780821007|SNOMEDCT_US|Malignant intraductal papillary-mucinous carcinoma of pancreas|8453/3
C1266075|T191|SY|C45754|NCI|Benign Mesothelioma of Mahaim|8454/0
C1266075|T191|SY|C45754|NCI|Cystic Tumor of Atrioventricular Node|8454/0
C1266075|T191|PT|C45754|NCI|Cystic Tumor of the Atrioventricular Node|8454/0
C1266075|T191|SY|C45754|NCI|Endodermal Rest|8454/0
C1266075|T191|SY|C45754|NCI|Intracardiac Endodermal Heterotopia|8454/0
C1266075|T191|SY|C45754|NCI|Mesothelioma of Atrioventricular Node|8454/0
C1266075|T191|SY|C45754|NCI|Tawarian Node|8454/0
C1266075|T191|PT|128693001|SNOMEDCT_US|Cystic tumor of atrio-ventricular node|8454/0
C1266075|T191|PTGB|128693001|SNOMEDCT_US|Cystic tumour of atrio-ventricular node|8454/0
C0334358|T191|PT|MTHU020327|ICPC2ICD10ENG|cystadenoma; papillary, serous, unspecified site|8460/0
C0334358|T191|PT|MTHU020339|ICPC2ICD10ENG|cystadenoma; serous, papillary, unspecified site|8460/0
C0334358|T191|PT|MTHU057305|ICPC2ICD10ENG|papillary; cystadenoma, serous, unspecified site|8460/0
C0334358|T191|PT|MTHU067558|ICPC2ICD10ENG|serous; cystadenoma, papillary, unspecified site|8460/0
C0334358|T191|PT|C4180|NCI|Papillary Serous Cystadenoma|8460/0
C0334358|T191|PT|X77nt|RCD|Papillary serous cystadenoma|8460/0
C0334358|T191|OA|BB816|RCDSY|Papill.serous cystadeno.NOS|8460/0
C0334358|T191|OP|BB816|RCDSY|Papillary serous cystadenoma NOS|8460/0
C0334358|T191|PT|22116003|SNOMEDCT_US|Papillary serous cystadenoma|8460/0
C0334358|T191|IS|22116003|SNOMEDCT_US|Papillary serous cystadenoma, NOS|8460/0
C3839578|T191|PT|703559005|SNOMEDCT_US|Serous borderline tumor, micropapillary variant|8460/2
C3839578|T191|PTGB|703559005|SNOMEDCT_US|Serous borderline tumour, micropapillary variant|8460/2
C3839578|T191|SY|703559005|SNOMEDCT_US|Serous carcinoma, non-invasive, low grade|8460/2
C3839184|T191|SY|0000029964|CHV|adenocarcinomas papillary serous|8460/3
C3839184|T191|PT|0000029964|CHV|papillary serous adenocarcinoma|8460/3
C3839184|T191|SY|0000029964|CHV|serous papillary adenocarcinoma|8460/3
C3839184|T191|PN|NOCODE|MTH|Papillary Serous Cystadenocarcinoma|8460/3
C3839184|T191|PT|C6882|NCI|Micropapillary Serous Carcinoma|8460/3
C3839184|T191|SY|C8377|NCI|Papillary Serous Adenocarcinoma|8460/3
C3839184|T191|SY|C8377|NCI|Papillary Serous Carcinoma|8460/3
C3839184|T191|PT|C8377|NCI|Papillary Serous Cystadenocarcinoma|8460/3
C3839184|T191|PT|CDR0000044781|NCI_NCI-GLOSS|papillary serous carcinoma|8460/3
C3839184|T191|OA|BB818|RCD|Papillary serous adenoca|8460/3
C3839184|T191|IS|BB818|RCD|Papillary serous adenocarcinoma|8460/3
C3839184|T191|OA|BB818|RCD|Papillary serous cystadenoca|8460/3
C3839184|T191|OP|BB818|RCD|Papillary serous cystadenocarcinoma|8460/3
C3839184|T191|PT|703561001|SNOMEDCT_US|Low grade serous carcinoma|8460/3
C3839184|T191|OAS|90282004|SNOMEDCT_US|Micropapillary serous carcinoma|8460/3
C3839184|T191|SY|703561001|SNOMEDCT_US|Micropapillary serous carcinoma|8460/3
C3839184|T191|OAS|90282004|SNOMEDCT_US|Papillary serous adenocarcinoma|8460/3
C3839184|T191|OAP|90282004|SNOMEDCT_US|Papillary serous cystadenocarcinoma|8460/3
C0334360|T191|PT|C4181|NCI|Serous Surface Papilloma|8461/0
C0334360|T191|PT|Xa98p|RCD|Serous surface papilloma|8461/0
C0334360|T191|OA|BB819|RCDSY|Serous surface papill.NOS|8461/0
C0334360|T191|OP|BB819|RCDSY|Serous surface papilloma NOS|8461/0
C0334360|T191|PT|67073007|SNOMEDCT_US|Serous surface papilloma|8461/0
C0334360|T191|IS|67073007|SNOMEDCT_US|Serous surface papilloma, NOS|8461/0
C0334361|T191|PN|NOCODE|MTH|Extraovarian primary peritoneal carcinoma|8461/3
C0334361|T191|PT|C4182|NCI|Serous Surface Papillary Carcinoma|8461/3
C0334361|T191|AB|BB81B|RCD|Serous surface papillary ca|8461/3
C0334361|T191|PT|BB81B|RCD|Serous surface papillary carcinoma|8461/3
C0334361|T191|SY|716649003|SNOMEDCT_US|EOPPC - Extraovarian primary peritoneal carcinoma|8461/3
C0334361|T191|PT|716649003|SNOMEDCT_US|Extraovarian primary peritoneal carcinoma|8461/3
C3839280|T191|PT|703563003|SNOMEDCT_US|High grade serous carcinoma|8461/3
C0334361|T191|SY|716649003|SNOMEDCT_US|Primary peritoneal serous carcinoma|8461/3
C0334361|T191|OAP|15674004|SNOMEDCT_US|Serous surface papillary carcinoma|8461/3
C0334361|T191|SY|716649003|SNOMEDCT_US|Serous surface papillary carcinoma|8461/3
C0334362|T191|SY|C4183|NCI|Borderline Malignancy Papillary Serous Cystadenoma|8462/1
C0334362|T191|PT|C4183|NCI|Borderline Papillary Serous Cystadenoma|8462/1
C0334362|T191|SY|C4183|NCI|Low Malignancy Potential Papillary Serous Cystadenoma|8462/1
C0334362|T191|SY|C4183|NCI|Low Malignant Potential Papillary Serous Neoplasm|8462/1
C0334362|T191|SY|C4183|NCI|Low Malignant Potential Papillary Serous Tumor|8462/1
C0334362|T191|SY|C4183|NCI|Papillary Serous Neoplasm of Low Malignant Potential|8462/1
C0334362|T191|SY|C4183|NCI|Papillary Serous Tumor of Low Malignant Potential|8462/1
C0334362|T191|DN|C4183|NCI_CTRP|Borderline Papillary Serous Cystadenoma|8462/1
C0334362|T191|SY|CDR0000685855|PDQ|borderline malignancy papillary serous cystadenoma|8462/1
C0334362|T191|PT|CDR0000685855|PDQ|borderline papillary serous cystadenoma|8462/1
C0334362|T191|SY|CDR0000685855|PDQ|low malignancy potential papillary serous cystadenoma|8462/1
C0334362|T191|SY|CDR0000685855|PDQ|low malignant potential papillary serous neoplasm|8462/1
C0334362|T191|SY|CDR0000685855|PDQ|low malignant potential papillary serous tumor|8462/1
C0334362|T191|SY|CDR0000685855|PDQ|papillary serous neoplasm of low malignant potential|8462/1
C0334362|T191|SY|CDR0000685855|PDQ|papillary serous tumor of low malignant potential|8462/1
C0334362|T191|AB|BB817|RCD|Papill ser cystadenom-bord mal|8462/1
C0334362|T191|AB|BB817|RCD|Papill ser tum low malig poten|8462/1
C0334362|T191|PT|BB817|RCD|Papillary serous cystadenoma - borderline malignancy|8462/1
C0334362|T191|SY|BB817|RCD|Papillary serous tumour of low malignant potential|8462/1
C0334362|T191|SY|BB817|RCDAE|Papillary serous tumor of low malignant potential|8462/1
C0334362|T191|AB|BB817|RCDSY|Pap ser cystad, bordl malig|8462/1
C0334362|T191|SY|BB817|RCDSY|Papillary serous cystadenoma, borderline malignancy|8462/1
C0334362|T191|SY|128851000|SNOMEDCT_US|Atypical proliferative papillary serous tumor|8462/1
C0334362|T191|SYGB|128851000|SNOMEDCT_US|Atypical proliferative papillary serous tumour|8462/1
C0334362|T191|OAP|189697000|SNOMEDCT_US|Papillary serous cystadenoma - borderline malignancy|8462/1
C0334362|T191|OF|189697000|SNOMEDCT_US|Papillary serous cystadenoma - borderline malignancy|8462/1
C0334362|T191|SY|128851000|SNOMEDCT_US|Papillary serous cystadenoma, borderline malignancy|8462/1
C0334362|T191|OAP|112678007|SNOMEDCT_US|Papillary serous cystadenoma, borderline malignancy|8462/1
C0334362|T191|IS|112678007|SNOMEDCT_US|Papillary serous cystadenoma, borderline malignancy -RETIRED-|8462/1
C0334362|T191|OF|112678007|SNOMEDCT_US|Papillary serous cystadenoma, borderline malignancy -RETIRED-|8462/1
C0334362|T191|SY|128851000|SNOMEDCT_US|Papillary serous tumor of low malignant potential|8462/1
C0334362|T191|IS|112678007|SNOMEDCT_US|Papillary serous tumor of low malignant potential|8462/1
C0334362|T191|SYGB|128851000|SNOMEDCT_US|Papillary serous tumour of low malignant potential|8462/1
C0334362|T191|PT|128851000|SNOMEDCT_US|Serous papillary cystic tumor of borderline malignancy|8462/1
C0334362|T191|PTGB|128851000|SNOMEDCT_US|Serous papillary cystic tumour of borderline malignancy|8462/1
C1511269|T191|OP|C7315|NCI|Borderline Ovarian Serous Surface Papillary Neoplasm|8463/1
C1511269|T191|OP|C7315|NCI|Borderline Ovarian Serous Surface Papillary Tumor|8463/1
C1511269|T191|PT|C7315|NCI|Borderline Ovarian Serous Surface Papillary Tumor|8463/1
C1266076|T191|PT|128694007|SNOMEDCT_US|Serous surface papillary tumor of borderline malignancy|8463/1
C1266076|T191|PTGB|128694007|SNOMEDCT_US|Serous surface papillary tumour of borderline malignancy|8463/1
C0010635|T191|PT|0046144|CCPSS|CYSTADENOMA MUCINOUS|8470/0
C0010635|T191|SY|0000029965|CHV|adenoma mucinous|8470/0
C0010635|T191|SY|0000003543|CHV|cystadenoma mucinous|8470/0
C0010635|T191|PT|0000029965|CHV|mucinous adenoma|8470/0
C0010635|T191|PT|0000003543|CHV|mucinous cystadenoma|8470/0
C0010635|T191|SY|0000003543|CHV|mucinous cystadenomas|8470/0
C0010635|T191|PT|MTHU020311|ICPC2ICD10ENG|cystadenoma; mucinous, unspecified site|8470/0
C0010635|T191|PT|MTHU020330|ICPC2ICD10ENG|cystadenoma; pseudomucinous, unspecified site|8470/0
C0010635|T191|PT|MTHU020859|ICPC2ICD10ENG|cystoma; mucinous, unspecified site|8470/0
C0010635|T191|PT|MTHU050445|ICPC2ICD10ENG|mucinous; cystadenoma, unspecified site|8470/0
C0010635|T191|PT|MTHU050449|ICPC2ICD10ENG|mucinous; cystoma, unspecified site|8470/0
C0010635|T191|PT|MTHU062300|ICPC2ICD10ENG|pseudomucinous; cystadenoma, unspecified site|8470/0
C2063870|T191|PT|38691|MEDCIN|cystic mucinous tumor of pancreas with moderate dysplasia|8470/0
C2063870|T191|SY|38691|MEDCIN|mucinous cystic neoplasm with moderate dysplasia|8470/0
C0010635|T191|MH|D018291|MSH|Cystadenoma, Mucinous|8470/0
C0010635|T191|PM|D018291|MSH|Cystadenomas, Mucinous|8470/0
C0010635|T191|PM|D018291|MSH|Mucinous Cystadenoma|8470/0
C0010635|T191|PM|D018291|MSH|Mucinous Cystadenomas|8470/0
C0010635|T191|SY|C2973|NCI|Mucinous Adenoma|8470/0
C0010635|T191|PT|C2973|NCI|Mucinous Cystadenoma|8470/0
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Neoplasm of Pancreas with Moderate Dysplasia|8470/0
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Neoplasm of the Pancreas with Moderate Dysplasia|8470/0
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor of Pancreas with Moderate Dysplasia|8470/0
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor of the Pancreas with Moderate Dysplasia|8470/0
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor with Moderate Dysplasia|8470/0
C0010635|T191|SY|C2973|NCI|Mucinous Cystoma|8470/0
C2063870|T191|SY|C6883|NCI|Pancreatic Borderline Mucinous Cystic Neoplasm|8470/0
C2063870|T191|SY|C6883|NCI|Pancreatic Low Grade Malignant Mucinous Cystic Neoplasm|8470/0
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Intermediate Grade Dysplasia|8470/0
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Intermediate-Grade Dysplasia|8470/0
C2987179|T191|SY|C95483|NCI|Pancreatic Mucinous Cystic Neoplasm with Low Grade Dysplasia|8470/0
C2987179|T191|SY|C95483|NCI|Pancreatic Mucinous Cystic Neoplasm with Low-Grade Dysplasia|8470/0
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Moderate Dysplasia|8470/0
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Tumor with Moderate Dysplasia|8470/0
C2063870|T191|PT|C6883|NCI|Pancreatic Mucinous-Cystic Neoplasm with Intermediate Grade Dysplasia|8470/0
C2987179|T191|PT|C95483|NCI|Pancreatic Mucinous-Cystic Neoplasm with Low Grade Dysplasia|8470/0
C0010635|T191|SY|C2973|NCI|Pseudomucinous Cystadenoma|8470/0
C0010635|T191|PT|C2973|NCI_CDISC|ADENOMA, MUCINOUS, BENIGN|8470/0
C0010635|T191|SY|C2973|NCI_CDISC|Mucinous Adenoma|8470/0
C0010635|T191|SY|C2973|NCI_CDISC|Mucinous Cystoma|8470/0
C0010635|T191|SY|C2973|NCI_CDISC|Pseudomucinous Cystadenoma|8470/0
C0010635|T191|PT|BB820|RCD|Mucinous adenoma|8470/0
C0010635|T191|PT|Xa98q|RCD|Mucinous cystadenoma|8470/0
C0010635|T191|SY|Xa98q|RCD|Mucinous cystoma|8470/0
C0010635|T191|SY|Xa98q|RCD|Pseudomucinous cystadenoma|8470/0
C0010635|T191|SY|Xa98q|RCDSY|Mucinous cystadenoma NOS|8470/0
C0010635|T191|PT|33170000|SNOMEDCT_US|Mucinous adenoma|8470/0
C0010635|T191|OAP|189691004|SNOMEDCT_US|Mucinous cystadenoma|8470/0
C0010635|T191|OF|189691004|SNOMEDCT_US|Mucinous cystadenoma|8470/0
C0010635|T191|PT|67182003|SNOMEDCT_US|Mucinous cystadenoma|8470/0
C0010635|T191|IS|67182003|SNOMEDCT_US|Mucinous cystadenoma, NOS|8470/0
C4518358|T191|PT|734054004|SNOMEDCT_US|Mucinous cystic neoplasm with low-grade intraepithelial neoplasia|8470/0
C2063870|T191|OAP|128899000|SNOMEDCT_US|Mucinous cystic tumor with moderate dysplasia|8470/0
C2063870|T191|OAP|128899000|SNOMEDCT_US|Mucinous cystic tumour with moderate dysplasia|8470/0
C0010635|T191|SY|67182003|SNOMEDCT_US|Mucinous cystoma|8470/0
C0010635|T191|SY|67182003|SNOMEDCT_US|Pseudomucinous cystadenoma|8470/0
C0010635|T191|IS|67182003|SNOMEDCT_US|Pseudomucinous cystadenoma, NOS|8470/0
C2063870|T191|PT|38691|MEDCIN|cystic mucinous tumor of pancreas with moderate dysplasia|8470/1
C2063870|T191|SY|38691|MEDCIN|mucinous cystic neoplasm with moderate dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Neoplasm of Pancreas with Moderate Dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Neoplasm of the Pancreas with Moderate Dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor of Pancreas with Moderate Dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor of the Pancreas with Moderate Dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor with Moderate Dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Pancreatic Borderline Mucinous Cystic Neoplasm|8470/1
C2063870|T191|SY|C6883|NCI|Pancreatic Low Grade Malignant Mucinous Cystic Neoplasm|8470/1
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Intermediate Grade Dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Intermediate-Grade Dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Moderate Dysplasia|8470/1
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Tumor with Moderate Dysplasia|8470/1
C2063870|T191|PT|C6883|NCI|Pancreatic Mucinous-Cystic Neoplasm with Intermediate Grade Dysplasia|8470/1
C2063870|T191|OAP|128899000|SNOMEDCT_US|Mucinous cystic tumor with moderate dysplasia|8470/1
C2063870|T191|OAP|128899000|SNOMEDCT_US|Mucinous cystic tumour with moderate dysplasia|8470/1
C2987185|T191|SY|C95493|NCI|Pancreatic Mucinous Cystic Neoplasm with High Grade Dysplasia|8470/2
C2987185|T191|PT|C95493|NCI|Pancreatic Mucinous-Cystic Neoplasm with High Grade Dysplasia|8470/2
C1518874|T191|PT|C41245|NCI|Pancreatic Non-Invasive Mucinous Cystadenocarcinoma|8470/2
C1518874|T191|OP|C41245|NCI|Pancreatic Non-Invasive Mucinous Cystadenocarcinoma|8470/2
C1266078|T191|PT|128900005|SNOMEDCT_US|Mucinous cystadenocarcinoma, non-invasive|8470/2
C4518360|T191|PT|734056002|SNOMEDCT_US|Mucinous cystic neoplasm with high-grade intraepithelial neoplasia|8470/2
C0206699|T191|PT|0000021031|CHV|mucinous cystadenocarcinoma|8470/3
C0206699|T191|PT|MTHU020292|ICPC2ICD10ENG|cystadenocarcinoma; mucinous, unspecified site|8470/3
C0206699|T191|PT|MTHU020298|ICPC2ICD10ENG|cystadenocarcinoma; pseudomucinous, unspecified site|8470/3
C0206699|T191|PT|MTHU050440|ICPC2ICD10ENG|mucinous; cystadenocarcinoma, unspecified site|8470/3
C0206699|T191|PT|MTHU062296|ICPC2ICD10ENG|pseudomucinous; cystadenocarcinoma, unspecified site|8470/3
C0206699|T191|MH|D018282|MSH|Cystadenocarcinoma, Mucinous|8470/3
C0206699|T191|PM|D018282|MSH|Cystadenocarcinomas, Mucinous|8470/3
C0206699|T191|PM|D018282|MSH|Mucinous Cystadenocarcinoma|8470/3
C0206699|T191|PM|D018282|MSH|Mucinous Cystadenocarcinomas|8470/3
C0206699|T191|PT|C3776|NCI|Mucinous Cystadenocarcinoma|8470/3
C0206699|T191|SY|TCGA|NCI|Mucinous Cystadenocarcinoma|8470/3
C1518870|T191|OP|C41246|NCI|Pancreatic Invasive Mucinous Cystadenocarcinoma|8470/3
C1518870|T191|SY|C41246|NCI|Pancreatic Mucinous Cystic Neoplasm with an Associated Invasive Carcinoma|8470/3
C1518870|T191|PT|C41246|NCI|Pancreatic Mucinous-Cystic Neoplasm with an Associated Invasive Carcinoma|8470/3
C0206699|T191|SY|C3776|NCI|Pseudomucinous Adenocarcinoma|8470/3
C0206699|T191|SY|C3776|NCI|Pseudomucinous Cystadenocarcinoma|8470/3
C0206699|T191|PT|Xa98r|RCD|Mucinous cystadenocarcinoma|8470/3
C0206699|T191|SY|Xa98r|RCD|Pseudomucinous adenocarcinoma|8470/3
C0206699|T191|AB|Xa98r|RCD|Pseudomucinous cystadenoca|8470/3
C0206699|T191|SY|Xa98r|RCD|Pseudomucinous cystadenocarcinoma|8470/3
C0206699|T191|OA|BB81E|RCDSY|Mucinous cystadenoca. NOS|8470/3
C0206699|T191|OP|BB81E|RCDSY|Mucinous cystadenocarcinoma NOS|8470/3
C0206699|T191|PT|79143006|SNOMEDCT_US|Mucinous cystadenocarcinoma|8470/3
C0206699|T191|IS|79143006|SNOMEDCT_US|Mucinous cystadenocarcinoma, NOS|8470/3
C4518373|T191|PT|734074006|SNOMEDCT_US|Mucinous cystic neoplasm with invasive carcinoma|8470/3
C0206699|T191|SY|79143006|SNOMEDCT_US|Pseudomucinous adenocarcinoma|8470/3
C0206699|T191|SY|79143006|SNOMEDCT_US|Pseudomucinous cystadenocarcinoma|8470/3
C0206699|T191|IS|79143006|SNOMEDCT_US|Pseudomucinous cystadenocarcinoma, NOS|8470/3
C0334363|T191|PT|MTHU020314|ICPC2ICD10ENG|cystadenoma; mucinous, papillary, unspecified site|8471/0
C0334363|T191|PT|MTHU020320|ICPC2ICD10ENG|cystadenoma; papillary, mucinous, unspecified site|8471/0
C0334363|T191|PT|MTHU020324|ICPC2ICD10ENG|cystadenoma; papillary, pseudomucinous, unspecified site|8471/0
C0334363|T191|PT|MTHU020333|ICPC2ICD10ENG|cystadenoma; pseudomucinous, papillary, unspecified site|8471/0
C0334363|T191|PT|MTHU050448|ICPC2ICD10ENG|mucinous; cystadenoma, papillary, unspecified site|8471/0
C0334363|T191|PT|MTHU057298|ICPC2ICD10ENG|papillary; cystadenoma, mucinous, unspecified site|8471/0
C0334363|T191|PT|MTHU057302|ICPC2ICD10ENG|papillary; cystadenoma, pseudomucinous, unspecified site|8471/0
C0334363|T191|PT|MTHU062303|ICPC2ICD10ENG|pseudomucinous; cystadenoma, papillary, unspecified site|8471/0
C0334363|T191|PT|C4184|NCI|Papillary Mucinous Cystadenoma|8471/0
C0334363|T191|SY|C4184|NCI|Papillary Pseudomucinous Cystadenoma|8471/0
C0334363|T191|AB|Xa98s|RCD|Papill pseudomucin cystadenoma|8471/0
C0334363|T191|PT|Xa98s|RCD|Papillary mucinous cystadenoma|8471/0
C0334363|T191|SY|Xa98s|RCD|Papillary pseudomucinous cystadenoma|8471/0
C0334363|T191|OA|BB81F|RCDSY|Papill.mucin.cystaden. NOS|8471/0
C0334363|T191|OP|BB81F|RCDSY|Papillary mucinous cystadenoma NOS|8471/0
C0334363|T191|PT|36721002|SNOMEDCT_US|Papillary mucinous cystadenoma|8471/0
C0334363|T191|IS|36721002|SNOMEDCT_US|Papillary mucinous cystadenoma, NOS|8471/0
C0334363|T191|SY|36721002|SNOMEDCT_US|Papillary pseudomucinous cystadenoma|8471/0
C0334363|T191|IS|36721002|SNOMEDCT_US|Papillary pseudomucinous cystadenoma, NOS|8471/0
C0334364|T191|PT|MTHU020293|ICPC2ICD10ENG|cystadenocarcinoma; mucinous, papillary, unspecified site|8471/3
C0334364|T191|PT|MTHU020294|ICPC2ICD10ENG|cystadenocarcinoma; papillary, mucinous, unspecified site|8471/3
C0334364|T191|PT|MTHU050441|ICPC2ICD10ENG|mucinous; cystadenocarcinoma, papillary, unspecified site|8471/3
C0334364|T191|PT|MTHU057289|ICPC2ICD10ENG|papillary; cystadenocarcinoma, mucinous, unspecified site|8471/3
C0334364|T191|PT|C65204|NCI|Papillary Mucinous Cystadenocarcinoma|8471/3
C0334364|T191|AB|BB81H|RCD|Papillary mucinous cystadenoca|8471/3
C0334364|T191|PT|BB81H|RCD|Papillary mucinous cystadenocarcinoma|8471/3
C0334364|T191|AB|BB81H|RCD|Papillary pseudomucin adenoca|8471/3
C0334364|T191|SY|BB81H|RCD|Papillary pseudomucinous adenocarcinoma|8471/3
C0334364|T191|PT|68880006|SNOMEDCT_US|Papillary mucinous cystadenocarcinoma|8471/3
C0334364|T191|SY|68880006|SNOMEDCT_US|Papillary pseudomucinous adenocarcinoma|8471/3
C0334364|T191|SY|68880006|SNOMEDCT_US|Papillary pseudomucinous cystadenocarcinoma|8471/3
C2063870|T191|PT|38691|MEDCIN|cystic mucinous tumor of pancreas with moderate dysplasia|8472/1
C2063870|T191|SY|38691|MEDCIN|mucinous cystic neoplasm with moderate dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Neoplasm of Pancreas with Moderate Dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Neoplasm of the Pancreas with Moderate Dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor of Pancreas with Moderate Dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor of the Pancreas with Moderate Dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Mucinous Cystic Tumor with Moderate Dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Pancreatic Borderline Mucinous Cystic Neoplasm|8472/1
C2063870|T191|SY|C6883|NCI|Pancreatic Low Grade Malignant Mucinous Cystic Neoplasm|8472/1
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Intermediate Grade Dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Intermediate-Grade Dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Neoplasm with Moderate Dysplasia|8472/1
C2063870|T191|SY|C6883|NCI|Pancreatic Mucinous Cystic Tumor with Moderate Dysplasia|8472/1
C2063870|T191|PT|C6883|NCI|Pancreatic Mucinous-Cystic Neoplasm with Intermediate Grade Dysplasia|8472/1
C0334365|T191|AB|BB81D|RCD|Mucin cystadenom-bord malign|8472/1
C0334365|T191|PT|BB81D|RCD|Mucinous cystadenoma - borderline malignancy|8472/1
C0334365|T191|AB|BB81D|RCD|Mucinous tumour low malig pot|8472/1
C0334365|T191|SY|BB81D|RCD|Mucinous tumour of low malignant potential|8472/1
C0334365|T191|AB|BB81D|RCD|Pseudomuc cystadenom-bord mal|8472/1
C0334365|T191|SY|BB81D|RCD|Pseudomucinous cystadenoma - borderline malignancy|8472/1
C0334365|T191|AB|BB81D|RCDAE|Mucinous tumor low malig pot|8472/1
C0334365|T191|SY|BB81D|RCDAE|Mucinous tumor of low malignant potential|8472/1
C0334365|T191|SY|128852007|SNOMEDCT_US|Atypical proliferative mucinous tumor|8472/1
C0334365|T191|SYGB|128852007|SNOMEDCT_US|Atypical proliferative mucinous tumour|8472/1
C0334365|T191|SY|128852007|SNOMEDCT_US|Mucinous borderline tumor|8472/1
C0334365|T191|SYGB|128852007|SNOMEDCT_US|Mucinous borderline tumour|8472/1
C0334365|T191|SY|128852007|SNOMEDCT_US|Mucinous cystadenoma - borderline malignancy|8472/1
C0334365|T191|OAP|85842001|SNOMEDCT_US|Mucinous cystadenoma, borderline malignancy|8472/1
C0334365|T191|SY|128852007|SNOMEDCT_US|Mucinous cystadenoma, borderline malignancy|8472/1
C0334365|T191|IS|85842001|SNOMEDCT_US|Mucinous cystadenoma, borderline malignancy -RETIRED-|8472/1
C0334365|T191|OF|85842001|SNOMEDCT_US|Mucinous cystadenoma, borderline malignancy -RETIRED-|8472/1
C0334365|T191|PT|128852007|SNOMEDCT_US|Mucinous cystic tumor of borderline malignancy|8472/1
C2063870|T191|OAP|128899000|SNOMEDCT_US|Mucinous cystic tumor with moderate dysplasia|8472/1
C0334365|T191|PTGB|128852007|SNOMEDCT_US|Mucinous cystic tumour of borderline malignancy|8472/1
C2063870|T191|OAP|128899000|SNOMEDCT_US|Mucinous cystic tumour with moderate dysplasia|8472/1
C0334365|T191|SY|128852007|SNOMEDCT_US|Mucinous tumor of low malignant potential|8472/1
C0334365|T191|IS|85842001|SNOMEDCT_US|Mucinous tumor, NOS, of low malignant potential|8472/1
C0334365|T191|SYGB|128852007|SNOMEDCT_US|Mucinous tumour of low malignant potential|8472/1
C0334365|T191|SY|128852007|SNOMEDCT_US|Pseudomucinous cystadenoma - borderline malignancy|8472/1
C0334365|T191|IS|85842001|SNOMEDCT_US|Pseudomucinous cystadenoma, borderline malignancy|8472/1
C0334365|T191|SY|128852007|SNOMEDCT_US|Pseudomucinous cystadenoma, borderline malignancy|8472/1
C0334366|T191|PT|MTHU057314|ICPC2ICD10ENG|papillary; tumor, mucinous, of low malignant potential|8473/1
C0334366|T191|PT|MTHU077130|ICPC2ICD10ENG|tumor; papillary, mucinous, of low malignant potential|8473/1
C0334366|T191|PN|NOCODE|MTH|Papillary mucinous cystadenoma, borderline malignancy|8473/1
C0334366|T191|SY|C4186|NCI|Borderline Malignancy Papillary Mucinous Cystadenoma|8473/1
C0334366|T191|SY|C4186|NCI|Borderline Malignancy Papillary Pseudomucinous Cystadenoma|8473/1
C0334366|T191|PT|C4186|NCI|Borderline Papillary Mucinous Cystadenoma|8473/1
C0334366|T191|SY|C4186|NCI|Borderline Papillary Pseudomucinous Cystadenoma|8473/1
C0334366|T191|SY|C4186|NCI|Low Malignancy Potential Papillary Mucinous Cystadenoma|8473/1
C0334366|T191|SY|C4186|NCI|Low Malignancy Potential Papillary Pseudomucinous Cystadenoma|8473/1
C0334366|T191|SY|C4186|NCI|Papillary Mucinous Neoplasm of Low Malignant Potential|8473/1
C0334366|T191|SY|C4186|NCI|Papillary Mucinous Tumor of Low Malignant Potential|8473/1
C0334366|T191|AB|BB81G|RCD|Papill muc cystadenom-bord mal|8473/1
C0334366|T191|AB|BB81G|RCD|Papill muc tum low malig poten|8473/1
C0334366|T191|PT|BB81G|RCD|Papillary mucinous cystadenoma - borderline malignancy|8473/1
C0334366|T191|SY|BB81G|RCD|Papillary mucinous tumour of low malignant potential|8473/1
C0334366|T191|SY|BB81G|RCDAE|Papillary mucinous tumor of low malignant potential|8473/1
C0334366|T191|SY|128853002|SNOMEDCT_US|Papillary mucinous cystadenoma - borderline malignancy|8473/1
C0334366|T191|OAP|14278004|SNOMEDCT_US|Papillary mucinous cystadenoma, borderline malignancy|8473/1
C0334366|T191|PT|128853002|SNOMEDCT_US|Papillary mucinous cystadenoma, borderline malignancy|8473/1
C0334366|T191|IS|14278004|SNOMEDCT_US|Papillary mucinous cystadenoma, borderline malignancy -RETIRED-|8473/1
C0334366|T191|OF|14278004|SNOMEDCT_US|Papillary mucinous cystadenoma, borderline malignancy -RETIRED-|8473/1
C0334366|T191|IS|14278004|SNOMEDCT_US|Papillary mucinous tumor of low malignant potential|8473/1
C0334366|T191|SY|128853002|SNOMEDCT_US|Papillary mucinous tumor of low malignant potential|8473/1
C0334366|T191|SYGB|128853002|SNOMEDCT_US|Papillary mucinous tumour of low malignant potential|8473/1
C0334366|T191|IS|14278004|SNOMEDCT_US|Papillary pseudomucinous cystadenoma, borderline malignancy|8473/1
C0334366|T191|SY|128853002|SNOMEDCT_US|Papillary pseudomucinous cystadenoma, borderline malignancy|8473/1
C3840171|T191|PT|703564009|SNOMEDCT_US|Seromucinous cystadenoma|8474/0
C3839681|T191|PT|703565005|SNOMEDCT_US|Seromucinous borderline tumor|8474/1
C3839681|T191|PTGB|703565005|SNOMEDCT_US|Seromucinous borderline tumour|8474/1
C3839681|T191|SY|703565005|SNOMEDCT_US|Seromucinous tumor, atypical proliferative|8474/1
C3839681|T191|SYGB|703565005|SNOMEDCT_US|Seromucinous tumour, atypical proliferative|8474/1
C3840227|T191|PT|703568007|SNOMEDCT_US|Seromucinous carcinoma|8474/3
C0010635|T191|PT|0046144|CCPSS|CYSTADENOMA MUCINOUS|8480/0
C0010635|T191|SY|0000029965|CHV|adenoma mucinous|8480/0
C0010635|T191|SY|0000003543|CHV|cystadenoma mucinous|8480/0
C0010635|T191|PT|0000029965|CHV|mucinous adenoma|8480/0
C0010635|T191|PT|0000003543|CHV|mucinous cystadenoma|8480/0
C0010635|T191|SY|0000003543|CHV|mucinous cystadenomas|8480/0
C0010635|T191|PT|MTHU020311|ICPC2ICD10ENG|cystadenoma; mucinous, unspecified site|8480/0
C0010635|T191|PT|MTHU020330|ICPC2ICD10ENG|cystadenoma; pseudomucinous, unspecified site|8480/0
C0010635|T191|PT|MTHU020859|ICPC2ICD10ENG|cystoma; mucinous, unspecified site|8480/0
C0010635|T191|PT|MTHU050445|ICPC2ICD10ENG|mucinous; cystadenoma, unspecified site|8480/0
C0010635|T191|PT|MTHU050449|ICPC2ICD10ENG|mucinous; cystoma, unspecified site|8480/0
C0010635|T191|PT|MTHU062300|ICPC2ICD10ENG|pseudomucinous; cystadenoma, unspecified site|8480/0
C0010635|T191|MH|D018291|MSH|Cystadenoma, Mucinous|8480/0
C0010635|T191|PM|D018291|MSH|Cystadenomas, Mucinous|8480/0
C0010635|T191|PM|D018291|MSH|Mucinous Cystadenoma|8480/0
C0010635|T191|PM|D018291|MSH|Mucinous Cystadenomas|8480/0
C0010635|T191|SY|C2973|NCI|Mucinous Adenoma|8480/0
C0010635|T191|PT|C2973|NCI|Mucinous Cystadenoma|8480/0
C0010635|T191|SY|C2973|NCI|Mucinous Cystoma|8480/0
C0010635|T191|SY|C2973|NCI|Pseudomucinous Cystadenoma|8480/0
C0010635|T191|PT|C2973|NCI_CDISC|ADENOMA, MUCINOUS, BENIGN|8480/0
C0010635|T191|SY|C2973|NCI_CDISC|Mucinous Adenoma|8480/0
C0010635|T191|SY|C2973|NCI_CDISC|Mucinous Cystoma|8480/0
C0010635|T191|SY|C2973|NCI_CDISC|Pseudomucinous Cystadenoma|8480/0
C0010635|T191|PT|BB820|RCD|Mucinous adenoma|8480/0
C0010635|T191|PT|Xa98q|RCD|Mucinous cystadenoma|8480/0
C0010635|T191|SY|Xa98q|RCD|Mucinous cystoma|8480/0
C0010635|T191|SY|Xa98q|RCD|Pseudomucinous cystadenoma|8480/0
C0010635|T191|SY|Xa98q|RCDSY|Mucinous cystadenoma NOS|8480/0
C0010635|T191|PT|33170000|SNOMEDCT_US|Mucinous adenoma|8480/0
C0010635|T191|OAP|189691004|SNOMEDCT_US|Mucinous cystadenoma|8480/0
C0010635|T191|OF|189691004|SNOMEDCT_US|Mucinous cystadenoma|8480/0
C0010635|T191|PT|67182003|SNOMEDCT_US|Mucinous cystadenoma|8480/0
C0010635|T191|IS|67182003|SNOMEDCT_US|Mucinous cystadenoma, NOS|8480/0
C0010635|T191|SY|67182003|SNOMEDCT_US|Mucinous cystoma|8480/0
C0010635|T191|SY|67182003|SNOMEDCT_US|Pseudomucinous cystadenoma|8480/0
C0010635|T191|IS|67182003|SNOMEDCT_US|Pseudomucinous cystadenoma, NOS|8480/0
C1708747|T191|SY|C42598|NCI|Appendix Well Differentiated Mucinous Adenocarcinoma|8480/1
C1708747|T191|AB|C42598|NCI|LAMN|8480/1
C1708747|T191|SY|C42598|NCI|Low Grade Appendiceal Mucinous Neoplasm|8480/1
C1708747|T191|SY|C42598|NCI|Low Grade Appendix Mucinous Neoplasm|8480/1
C1708747|T191|PT|C42598|NCI|Low-Grade Appendiceal Mucinous Neoplasm|8480/1
C1708747|T191|SY|C42598|NCI|Low-Grade Appendix Mucinous Neoplasm|8480/1
C1708747|T191|PT|450896006|SNOMEDCT_US|Low grade appendiceal mucinous neoplasm|8480/1
C0007130|T191|PT|0024899|CCPSS|ADENOCARCINOMA MUCINOUS|8480/3
C0007130|T191|SY|0000002432|CHV|adenocarcinoma mucinous|8480/3
C0007130|T191|SY|0000002432|CHV|adenocarcinoma mucous|8480/3
C0007130|T191|SY|0000002432|CHV|colloid carcinoma|8480/3
C0007130|T191|PT|0000002432|CHV|mucinous adenocarcinoma|8480/3
C0007130|T191|SY|0000002432|CHV|mucinous carcinoma|8480/3
C0007130|T191|SY|0000002432|CHV|mucoid adenocarcinoma|8480/3
C0007130|T191|LA|LA26497-0|LNC|Colloid carcinoma|8480/3
C0007130|T191|LLT|10061564|MDR|Mucinous carcinoma|8480/3
C0007130|T191|PT|271463|MEDCIN|mucinous adenocarcinoma|8480/3
C0346020|T191|PT|357600|MEDCIN|Mucinous eccrine carcinoma of skin|8480/3
C0346020|T191|SY|357600|MEDCIN|skin neop malignant adnexa w/ eccrine differentiation mucinous carcinoma|8480/3
C0007130|T191|MH|D002288|MSH|Adenocarcinoma, Mucinous|8480/3
C0007130|T191|PM|D002288|MSH|Adenocarcinomas, Mucinous|8480/3
C0007130|T191|ET|D002288|MSH|Carcinoma, Colloid|8480/3
C0007130|T191|ET|D002288|MSH|Carcinoma, Mucinous|8480/3
C0007130|T191|PM|D002288|MSH|Carcinomas, Colloid|8480/3
C0007130|T191|PM|D002288|MSH|Carcinomas, Mucinous|8480/3
C0007130|T191|PM|D002288|MSH|Colloid Carcinoma|8480/3
C0007130|T191|PM|D002288|MSH|Colloid Carcinomas|8480/3
C0007130|T191|PM|D002288|MSH|Mucinous Adenocarcinoma|8480/3
C0007130|T191|PM|D002288|MSH|Mucinous Adenocarcinomas|8480/3
C0007130|T191|PM|D002288|MSH|Mucinous Carcinoma|8480/3
C0007130|T191|PM|D002288|MSH|Mucinous Carcinomas|8480/3
C0007130|T191|PN|NOCODE|MTH|Mucinous Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Colloid Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Colloid Carcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Gelatinous Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Gelatinous Carcinoma|8480/3
C0007130|T191|PT|C26712|NCI|Mucinous Adenocarcinoma|8480/3
C0007130|T191|SY|TCGA|NCI|Mucinous Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Mucinous Carcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Mucoid Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Mucoid Carcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Mucous Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI|Mucous Carcinoma|8480/3
C0007130|T191|PT|C26712|NCI_CDISC|ADENOCARCINOMA, MUCINOUS, MALIGNANT|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Colloid Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Colloid Carcinoma|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Gelatinous Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Gelatinous Carcinoma|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Mucinous Carcinoma|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Mucoid Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Mucoid Carcinoma|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Mucous Adenocarcinoma|8480/3
C0007130|T191|SY|C26712|NCI_CDISC|Mucous Carcinoma|8480/3
C0007130|T191|PT|CDR0000044289|NCI_NCI-GLOSS|mucinous carcinoma|8480/3
C0007130|T191|SY|BB821|RCD|Colloid adenocarcinoma|8480/3
C0007130|T191|SY|BB821|RCD|Colloid carcinoma|8480/3
C0007130|T191|SY|BB821|RCD|Gelatinous adenocarcinoma|8480/3
C0007130|T191|SY|BB821|RCD|Gelatinous carcinoma|8480/3
C0007130|T191|PT|BB821|RCD|Mucinous adenocarcinoma|8480/3
C0007130|T191|SY|BB821|RCD|Mucinous carcinoma|8480/3
C0346020|T191|AB|X78Sk|RCD|Mucinous ecc carcinoma of skin|8480/3
C0346020|T191|PT|X78Sk|RCD|Mucinous eccrine carcinoma|8480/3
C0346020|T191|SY|X78Sk|RCD|Mucinous eccrine carcinoma of skin|8480/3
C0007130|T191|SY|BB821|RCD|Mucoid adenocarcinoma|8480/3
C0007130|T191|SY|BB821|RCD|Mucoid carcinoma|8480/3
C0007130|T191|SY|BB821|RCD|Mucous adenocarcinoma|8480/3
C0007130|T191|SY|BB821|RCD|Mucous carcinoma|8480/3
C0346020|T191|AB|X78Sk|RCD|Primary mucinous carcinoma|8480/3
C0346020|T191|SY|X78Sk|RCD|Primary mucinous carcinoma of skin|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Colloid adenocarcinoma|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Colloid carcinoma|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Gelatinous adenocarcinoma|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Gelatinous carcinoma|8480/3
C0007130|T191|PT|72495009|SNOMEDCT_US|Mucinous adenocarcinoma|8480/3
C1302417|T191|PT|399449005|SNOMEDCT_US|Mucinous adenocarcinoma, intestinal type|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Mucinous carcinoma|8480/3
C0346020|T191|PT|254714008|SNOMEDCT_US|Mucinous eccrine carcinoma|8480/3
C0346020|T191|PT|399540006|SNOMEDCT_US|Mucinous eccrine carcinoma|8480/3
C0346020|T191|SY|254714008|SNOMEDCT_US|Mucinous eccrine carcinoma of skin|8480/3
C4518220|T191|PT|733884004|SNOMEDCT_US|Mucinous minimally invasive adenocarcinoma|8480/3
C4518375|T191|PT|734077004|SNOMEDCT_US|Mucinous tubular and spindle cell carcinoma|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Mucoid adenocarcinoma|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Mucoid carcinoma|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Mucous adenocarcinoma|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Mucous carcinoma|8480/3
C0346020|T191|SY|254714008|SNOMEDCT_US|Primary mucinous carcinoma of skin|8480/3
C0007130|T191|SY|72495009|SNOMEDCT_US|Pseudomyxoma peritonei with unknown primary site|8480/3
C0033822|T191|SY|0000010297|CHV|gelatinous ascites|8480/6
C0033822|T191|PT|0000050200|CHV|myxoma peritonei|8480/6
C0033822|T191|PT|0000010297|CHV|pseudomyxoma peritonei|8480/6
C0033822|T191|SY|NOCODE|DXP|PERITONITIS, MYXOMATOUS|8480/6
C0033822|T191|DI|U001608|DXP|PSEUDOMYXOMA PERITONEI|8480/6
C0033822|T191|PT|MTHU062307|ICPC2ICD10ENG|pseudomyxoma peritonei|8480/6
C0033822|T191|LLT|10028666|MDR|Myxoma peritonei|8480/6
C0033822|T191|LLT|10037138|MDR|Pseudomyxoma peritonei|8480/6
C0033822|T191|PT|10037138|MDR|Pseudomyxoma peritonei|8480/6
C0033822|T191|SY|31641|MEDCIN|pseudomyxoma peritonei|8480/6
C0033822|T191|PT|31641|MEDCIN|pseudomyxoma peritonei of peritoneum|8480/6
C0033822|T191|ET|D011553|MSH|Ascites, Gelatinous|8480/6
C0033822|T191|ET|D011553|MSH|Gelatinous Ascites|8480/6
C0033822|T191|MH|D011553|MSH|Pseudomyxoma Peritonei|8480/6
C0033822|T191|PM|D011553|MSH|Pseudomyxoma Peritonei Syndrome|8480/6
C0033822|T191|PM|D011553|MSH|Pseudomyxoma Peritonei Syndromes|8480/6
C0033822|T191|ET|D011553|MSH|Syndrome of Pseudomyxoma Peritonei|8480/6
C0033822|T191|PN|NOCODE|MTH|Pseudomyxoma Peritonei|8480/6
C0033822|T191|SY|C3345|NCI|Gelatinous Ascites|8480/6
C0033822|T191|SY|C3345|NCI|Mucinous Ascites|8480/6
C0033822|T191|SY|C3345|NCI|Myxoma Peritonei|8480/6
C0033822|T191|SY|C3345|NCI|Peritoneal Cavity Pseudomyxoma Peritonei|8480/6
C0033822|T191|PT|C3345|NCI|Pseudomyxoma Peritonei|8480/6
C0033822|T191|SY|C3345|NCI|Well Differentiated Peritoneal Mucinous Adenocarcinoma|8480/6
C0033822|T191|DN|C3345|NCI_CTRP|Pseudomyxoma Peritonei|8480/6
C0033822|T191|PT|CDR0000044256|NCI_NCI-GLOSS|pseudomyxoma peritonei|8480/6
C0033822|T191|SY|CDR0000040915|PDQ|malignant peritoneal pseudomyxoma peritonei|8480/6
C0033822|T191|SY|CDR0000040915|PDQ|malignant pseudomyxoma peritonei|8480/6
C0033822|T191|SY|CDR0000040915|PDQ|peritoneal cavity pseudomyxoma peritonei|8480/6
C0033822|T191|PSC|CDR0000040915|PDQ|pseudomyxoma peritonei|8480/6
C0033822|T191|PT|XaBAu|RCD|Pseudomyxoma peritonei|8480/6
C0033822|T191|PT|BB83.|RCDSY|Pseudomyxoma peritonei|8480/6
C0033822|T191|PT|307601000|SNOMEDCT_US|Pseudomyxoma peritonei|8480/6
C0033822|T191|PT|112679004|SNOMEDCT_US|Pseudomyxoma peritonei|8480/6
C0334368|T191|SY|0000029966|CHV|adenocarcinoma mucin secreting|8481/3
C0334368|T191|SY|0000029966|CHV|carcinoma mucin secreting|8481/3
C0334368|T191|PT|0000029966|CHV|mucin-producing adenocarcinoma|8481/3
C0334368|T191|PT|271464|MEDCIN|mucin-producing adenocarcinoma|8481/3
C0334368|T191|PT|C27379|NCI|Mucin-Producing Adenocarcinoma|8481/3
C0334368|T191|PT|C27825|NCI|Mucin-Producing Carcinoma|8481/3
C0334368|T191|PT|C27825|NCI_CPTAC|Mucin-Producing Carcinoma|8481/3
C0334368|T191|PT|BB84.|RCD|Mucin-producing adenocarcinoma|8481/3
C0334368|T191|SY|BB84.|RCD|Mucin-producing carcinoma|8481/3
C0334368|T191|SY|BB84.|RCD|Mucin-secreting adenocarcinoma|8481/3
C0334368|T191|SY|BB84.|RCD|Mucin-secreting carcinoma|8481/3
C0334368|T191|PT|900006|SNOMEDCT_US|Mucin-producing adenocarcinoma|8481/3
C0334368|T191|SY|900006|SNOMEDCT_US|Mucin-producing carcinoma|8481/3
C0334368|T191|SY|900006|SNOMEDCT_US|Mucin-secreting adenocarcinoma|8481/3
C0334368|T191|SY|900006|SNOMEDCT_US|Mucin-secreting carcinoma|8481/3
C1266079|T191|PT|C66953|NCI|Mucinous Adenocarcinoma, Endocervical Type|8482/3
C1266079|T191|PT|128695008|SNOMEDCT_US|Mucinous adenocarcinoma, endocervical type|8482/3
C3839471|T191|PT|703569004|SNOMEDCT_US|Mucinous adenocarcinoma, endocervical, gastric type|8482/3
C0206696|T191|SY|0000021028|CHV|adenocarcinoma cells ring signet|8490/3
C0206696|T191|SY|0000021028|CHV|carcinoma signet ring cell|8490/3
C0206696|T191|SY|0000021028|CHV|signet ring carcinoma|8490/3
C0206696|T191|PT|0000021028|CHV|signet ring cell carcinoma|8490/3
C0206696|T191|SY|0000021028|CHV|signet-ring cell carcinoma|8490/3
C4264447|T191|LA|LA26095-2|LNC|Poorly cohesive carcinoma|8490/3
C0206696|T191|LA|LA15444-5|LNC|Signet ring cell carcinoma|8490/3
C0206696|T191|LLT|10057266|MDR|Signet-ring cell carcinoma|8490/3
C0206696|T191|PT|10057266|MDR|Signet-ring cell carcinoma|8490/3
C1302700|T191|PT|355118|MEDCIN|Primary signet ring carcinoma of skin|8490/3
C0206696|T191|PT|271440|MEDCIN|signet ring cell carcinoma|8490/3
C1302700|T191|SY|355118|MEDCIN|skin neoplasm malignant w/apocrine differentiation primary signet ring carcinoma|8490/3
C0206696|T191|MH|D018279|MSH|Carcinoma, Signet Ring Cell|8490/3
C0206696|T191|ET|D018279|MSH|Signet Ring Cell Carcinoma|8490/3
C2987393|T191|PT|C95743|NCI|Gastric Poorly Cohesive Carcinoma|8490/3
C2987393|T191|SY|C95743|NCI|Poorly Cohesive Gastric Adenocarcinoma|8490/3
C2987393|T191|SY|C95743|NCI|Poorly Cohesive Gastric Carcinoma|8490/3
C0206696|T191|SY|C3774|NCI|Signet Ring Cell Adenocarcinoma|8490/3
C0206696|T191|PT|C3774|NCI|Signet Ring Cell Carcinoma|8490/3
C0206696|T191|SY|TCGA|NCI|Signet Ring Cell Carcinoma|8490/3
C0206696|T191|PT|CDR0000044297|NCI_NCI-GLOSS|signet ring cell carcinoma|8490/3
C1302700|T191|AB|Xa0C0|RCD|Prim signet ring carcinom-skin|8490/3
C1302700|T191|PT|Xa0C0|RCD|Primary signet ring carcinoma of skin|8490/3
C0206696|T191|SY|BB850|RCD|Signet ring carcinoma|8490/3
C0206696|T191|AB|BB850|RCD|Signet ring cell adenoca|8490/3
C0206696|T191|SY|BB850|RCD|Signet ring cell adenocarcinoma|8490/3
C0206696|T191|PT|BB850|RCD|Signet ring cell carcinoma|8490/3
C0206696|T191|OP|BB85z|RCDSY|Signet ring carcinoma NOS|8490/3
C4264447|T191|PT|725503008|SNOMEDCT_US|Poorly cohesive carcinoma|8490/3
C1302700|T191|PT|276738009|SNOMEDCT_US|Primary signet ring carcinoma of skin|8490/3
C0206696|T191|SY|87737001|SNOMEDCT_US|Signet ring carcinoma|8490/3
C1302700|T191|PT|399887008|SNOMEDCT_US|Signet ring carcinoma, primary cutaneous|8490/3
C0206696|T191|SY|87737001|SNOMEDCT_US|Signet ring cell adenocarcinoma|8490/3
C0206696|T191|PT|87737001|SNOMEDCT_US|Signet ring cell carcinoma|8490/3
C0206696|T191|OAP|189701002|SNOMEDCT_US|Signet ring cell carcinoma|8490/3
C0206696|T191|OF|189701002|SNOMEDCT_US|Signet ring cell carcinoma|8490/3
C1881801|T191|PN|NOCODE|MTH|Metastatic signet ring cell carcinoma|8490/6
C1881801|T191|PT|C66717|NCI|Metastatic Signet Ring Cell Carcinoma|8490/6
C1881801|T191|AB|BB851|RCD|Metastatic signet ring cell ca|8490/6
C1881801|T191|PT|BB851|RCD|Metastatic signet ring cell carcinoma|8490/6
C1881801|T191|PT|4305004|SNOMEDCT_US|Metastatic signet ring cell carcinoma|8490/6
C3273050|T191|PT|C96808|NCI|Bile Duct Papillary Neoplasm with Intermediate Grade Intraepithelial Neoplasia|850/30
C3273050|T191|SY|C96808|NCI|Intraductal Papillary Neoplasm with Intermediate Grade Intraepithelial Neoplasia|850/30
C0007124|T191|SY|0000002429|CHV|breast cancer intraductal|8500/2
C0007124|T191|SY|0000002429|CHV|breast carcinoma ductal situ|8500/2
C0007124|T191|SY|0000002429|CHV|breast ductal carcinoma in situ|8500/2
C0007124|T191|SY|0000002429|CHV|carcinoma ductal in situ|8500/2
C0007124|T191|SY|0000002429|CHV|carcinoma ductal situ|8500/2
C0007124|T191|SY|0000002429|CHV|carcinoma intraductal|8500/2
C0007124|T191|SY|0000002429|CHV|dci|8500/2
C0007124|T191|PT|0000002429|CHV|dcis|8500/2
C0007124|T191|SY|0000002429|CHV|ductal carcinoma in situ|8500/2
C0007124|T191|SY|0000002429|CHV|ductal carcinoma situ|8500/2
C0007124|T191|SY|0000002429|CHV|ductal in situ carcinoma|8500/2
C0007124|T191|SY|0000002429|CHV|in situ ductal carcinoma|8500/2
C0007124|T191|SY|0000002429|CHV|intraductal breast cancer|8500/2
C0007124|T191|SY|0000002429|CHV|intraductal carcinoma|8500/2
C0007124|T191|SY|0000002429|CHV|intraductal carcinoma breast|8500/2
C0007124|T191|ET|2016-0671|CSP|DCIS|8500/2
C0007124|T191|ET|2016-0671|CSP|ductal carcinoma in situ|8500/2
C0007124|T191|ET|2000-1867|CSP|intraductal carcinoma|8500/2
C0007124|T191|PT|HP:0030075|HPO|Ductal carcinoma in situ|8500/2
C0007124|T191|PT|D05.1|ICD10|Intraductal carcinoma in situ|8500/2
C0007124|T191|AB|D05.1|ICD10CM|Intraductal carcinoma in situ of breast|8500/2
C0007124|T191|HT|D05.1|ICD10CM|Intraductal carcinoma in situ of breast|8500/2
C0007124|T191|PT|MTHU003399|ICPC2ICD10ENG|adenocarcinoma; intraductal, noninfiltrating, breast|8500/2
C0007124|T191|PT|MTHU047381|ICPC2ICD10ENG|breast; carcinoma in situ, intraductal|8500/2
C0007124|T191|PT|MTHU047385|ICPC2ICD10ENG|breast; carcinoma, intraductal|8500/2
C0007124|T191|PT|MTHU047429|ICPC2ICD10ENG|breast; intraductal carcinoma|8500/2
C0007124|T191|PT|MTHU047428|ICPC2ICD10ENG|breast; intraductal carcinoma in situ|8500/2
C0007124|T191|PT|MTHU014710|ICPC2ICD10ENG|carcinoma in situ; intraductal, breast|8500/2
C0007124|T191|PT|MTHU014711|ICPC2ICD10ENG|carcinoma in situ; intraductal, unspecified site|8500/2
C0007124|T191|PT|MTHU014775|ICPC2ICD10ENG|carcinoma; intraductal, breast|8500/2
C0007124|T191|PT|MTHU014776|ICPC2ICD10ENG|carcinoma; intraductal, unspecified site|8500/2
C0007124|T191|PT|MTHU040055|ICPC2ICD10ENG|intraductal; carcinoma in situ, breast|8500/2
C0007124|T191|PT|MTHU040056|ICPC2ICD10ENG|intraductal; carcinoma in situ, unspecified site|8500/2
C0007124|T191|PT|MTHU040057|ICPC2ICD10ENG|intraductal; carcinoma, breast|8500/2
C0007124|T191|PT|MTHU040058|ICPC2ICD10ENG|intraductal; carcinoma, unspecified site|8500/2
C0007124|T191|LPN|LP57573-5|LNC|DCIS|8500/2
C0007124|T191|LLT|10007360|MDR|Carcinoma in situ of breast ductal|8500/2
C0007124|T191|LLT|10013806|MDR|Ductal carcinoma in situ|8500/2
C0007124|T191|SY|351623|MEDCIN|breast malignant carcinoma intraductal|8500/2
C0007124|T191|SY|361469|MEDCIN|breast neoplasm carcinoma in situ intraductal|8500/2
C0007124|T191|PT|361469|MEDCIN|Intraductal carcinoma in situ of breast|8500/2
C0007124|T191|PT|351623|MEDCIN|Intraductal carcinoma of breast|8500/2
C0007124|T191|ET|D002285|MSH|Carcinoma, Intraductal|8500/2
C0007124|T191|MH|D002285|MSH|Carcinoma, Intraductal, Noninfiltrating|8500/2
C0007124|T191|PM|D002285|MSH|Carcinoma, Noninfiltrating Intraductal|8500/2
C0007124|T191|PM|D002285|MSH|Carcinomas, Intraductal|8500/2
C0007124|T191|PM|D002285|MSH|Carcinomas, Noninfiltrating Intraductal|8500/2
C0007124|T191|ET|D002285|MSH|DCIS|8500/2
C0007124|T191|ET|D002285|MSH|Ductal Carcinoma In Situ|8500/2
C0007124|T191|PM|D002285|MSH|Intraductal Carcinoma|8500/2
C0007124|T191|ET|D002285|MSH|Intraductal Carcinoma, Noninfiltrating|8500/2
C0007124|T191|PM|D002285|MSH|Intraductal Carcinomas|8500/2
C0007124|T191|PM|D002285|MSH|Intraductal Carcinomas, Noninfiltrating|8500/2
C0007124|T191|PM|D002285|MSH|Noninfiltrating Intraductal Carcinoma|8500/2
C0007124|T191|PM|D002285|MSH|Noninfiltrating Intraductal Carcinomas|8500/2
C0007124|T191|PN|NOCODE|MTH|Noninfiltrating Intraductal Carcinoma|8500/2
C0007124|T191|AB|C2924|NCI|DCIS|8500/2
C0007124|T191|PT|C2924|NCI|Ductal Breast Carcinoma In Situ|8500/2
C0007124|T191|SY|C2924|NCI|Ductal Carcinoma In Situ|8500/2
C0007124|T191|SY|C2924|NCI|Ductal Carcinoma In Situ of Breast|8500/2
C0007124|T191|SY|C2924|NCI|Ductal Carcinoma In Situ of the Breast|8500/2
C0007124|T191|SY|C2924|NCI|Intraductal Breast Carcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Intraductal Carcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Intraductal Carcinoma of Breast|8500/2
C0007124|T191|SY|C2924|NCI|Intraductal Carcinoma of the Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Ductal Adenocarcinoma of Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Ductal Adenocarcinoma of the Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Ductal Breast Adenocarcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Ductal Breast Carcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Ductal Carcinoma of Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Ductal Carcinoma of the Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Intraductal Adenocarcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Intraductal Adenocarcinoma of Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Intraductal Adenocarcinoma of the Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Intraductal Breast Adenocarcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Non-Infiltrating Intraductal Carcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Ductal Adenocarcinoma of Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Ductal Adenocarcinoma of the Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Ductal Breast Adenocarcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Ductal Breast Carcinoma|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Ductal Carcinoma of Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Ductal Carcinoma of the Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Intraductal Adenocarcinoma of Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Intraductal Adenocarcinoma of the Breast|8500/2
C0007124|T191|SY|C2924|NCI|Non-Invasive Intraductal Breast Adenocarcinoma|8500/2
C0007124|T191|PT|C2924|NCI_CPTAC|Ductal Breast Carcinoma In Situ|8500/2
C0007124|T191|PT|10013806|NCI_CTEP-SDC|Ductal carcinoma in situ|8500/2
C0007124|T191|PT|CDR0000044394|NCI_NCI-GLOSS|DCIS|8500/2
C0007124|T191|PT|CDR0000045674|NCI_NCI-GLOSS|ductal carcinoma in situ|8500/2
C0007124|T191|PT|CDR0000046748|NCI_NCI-GLOSS|intraductal carcinoma|8500/2
C0007124|T191|AB|CDR0000039839|PDQ|DCIS|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|DCIS of the breast|8500/2
C0007124|T191|PT|CDR0000039839|PDQ|ductal breast carcinoma in situ|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|ductal cancer in situ of the breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|ductal carcinoma in situ|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Ductal Carcinoma in situ of Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|ductal carcinoma in situ of the breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|in situ ductal breast carcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|intraductal breast cancer|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|intraductal breast carcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Intraductal Carcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Intraductal Carcinoma of Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Intraductal Carcinoma of the Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Ductal Adenocarcinoma of Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Ductal Adenocarcinoma of the Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Ductal Breast Adenocarcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Ductal Breast Carcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Ductal Carcinoma of Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Ductal Carcinoma of the Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Intraductal Adenocarcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Intraductal Adenocarcinoma of Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Intraductal Adenocarcinoma of the Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Intraductal Breast Adenocarcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Infiltrating Intraductal Carcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Ductal Adenocarcinoma of Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Ductal Adenocarcinoma of the Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Ductal Breast Adenocarcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Ductal Breast Carcinoma|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Ductal Carcinoma of Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Ductal Carcinoma of the Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Intraductal Adenocarcinoma of Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Intraductal Adenocarcinoma of the Breast|8500/2
C0007124|T191|SY|CDR0000039839|PDQ|Non-Invasive Intraductal Breast Adenocarcinoma|8500/2
C0007124|T191|PT|Xa0bT|RCD|Intraduct carcinoma of breast|8500/2
C0007124|T191|AB|X78WW|RCD|Intraductal ca in situ breast|8500/2
C0007124|T191|SY|X77nz|RCD|Intraductal carcinoma|8500/2
C0007124|T191|PT|X78WW|RCD|Intraductal carcinoma in situ of breast|8500/2
C0007124|T191|AB|X77nz|RCD|Non-infiltr intraduct adenoca|8500/2
C0007124|T191|AB|X77nz|RCD|Non-infiltrat intraductal ca|8500/2
C0007124|T191|SY|X77nz|RCD|Non-infiltrating intraductal adenocarcinoma|8500/2
C0007124|T191|PT|X77nz|RCD|Non-infiltrating intraductal carcinoma|8500/2
C0007124|T191|OA|BB90.|RCDSY|Intraduct ca, noninfilt NOS|8500/2
C0007124|T191|OP|BB90.|RCDSY|Intraductal carcinoma, non-infiltrating NOS|8500/2
C1266081|T191|PT|128697000|SNOMEDCT_US|Cystic hypersecretory carcinoma|8500/2
C0007124|T191|SY|86616005|SNOMEDCT_US|DCIS|8500/2
C0007124|T191|SY|86616005|SNOMEDCT_US|Ductal carcinoma in situ|8500/2
C0007124|T191|IS|278053004|SNOMEDCT_US|Intraduct carcinoma of breast|8500/2
C0007124|T191|SY|86616005|SNOMEDCT_US|Intraductal adenocarcinoma, noninfiltrating|8500/2
C0007124|T191|IS|86616005|SNOMEDCT_US|Intraductal adenocarcinoma, noninfiltrating, NOS|8500/2
C0007124|T191|SY|86616005|SNOMEDCT_US|Intraductal carcinoma|8500/2
C0007124|T191|PT|109889007|SNOMEDCT_US|Intraductal carcinoma in situ of breast|8500/2
C0007124|T191|OAP|189338004|SNOMEDCT_US|Intraductal carcinoma in situ of breast|8500/2
C0007124|T191|OF|189338004|SNOMEDCT_US|Intraductal carcinoma in situ of breast|8500/2
C0007124|T191|OAP|278053004|SNOMEDCT_US|Intraductal carcinoma of breast|8500/2
C0007124|T191|PT|86616005|SNOMEDCT_US|Intraductal carcinoma, noninfiltrating|8500/2
C0007124|T191|SY|86616005|SNOMEDCT_US|Intraductal carcinoma, noninfiltrating, no ICD-O subtype|8500/2
C0007124|T191|SY|86616005|SNOMEDCT_US|Intraductal carcinoma, noninfiltrating, no International Classification of Diseases for Oncology subtype|8500/2
C0007124|T191|IS|86616005|SNOMEDCT_US|Intraductal carcinoma, noninfiltrating, NOS|8500/2
C0007124|T191|IS|86616005|SNOMEDCT_US|Intraductal carcinoma, NOS|8500/2
C0007124|T191|SY|86616005|SNOMEDCT_US|Non-infiltrating intraductal adenocarcinoma|8500/2
C0007124|T191|SY|86616005|SNOMEDCT_US|Non-infiltrating intraductal carcinoma|8500/2
C1134719|T191|PT|0042764|CCPSS|BREAST CANCER DUCTAL INFILTRATING|8500/3
C1134719|T191|SY|0000050852|CHV|breast cancer invasive ductal|8500/3
C1134719|T191|SY|0000056504|CHV|breast carcinoma ductal invasive|8500/3
C1134719|T191|SY|0000050852|CHV|cancer breast invasive ductal|8500/3
C1134719|T191|SY|0000054856|CHV|carcinoma ductal infiltrate|8500/3
C1134719|T191|SY|0000054856|CHV|carcinoma ductal infiltrated|8500/3
C1134719|T191|SY|0000056504|CHV|carcinoma infiltrating duct|8500/3
C1134719|T191|SY|0000054856|CHV|carcinomas ductal infiltrating|8500/3
C1134719|T191|SY|0000054856|CHV|ductal infiltrating carcinoma|8500/3
C1134719|T191|SY|0000050852|CHV|ductal invasive breast cancer|8500/3
C1134719|T191|PT|0000054856|CHV|infiltrating ductal carcinoma|8500/3
C1134719|T191|PT|0000050852|CHV|invasive ductal breast cancer|8500/3
C1134719|T191|PT|0000056504|CHV|invasive ductal breast carcinoma|8500/3
C1134719|T191|SY|0000056504|CHV|invasive ductal carcinoma breast|8500/3
C1134719|T191|PT|MTHU014743|ICPC2ICD10ENG|carcinoma; ductal, infiltrating, unspecified site|8500/3
C1134719|T191|PT|MTHU014744|ICPC2ICD10ENG|carcinoma; ductular, infiltrating, unspecified site|8500/3
C1134719|T191|PT|MTHU014770|ICPC2ICD10ENG|carcinoma; infiltrating duct, unspecified site|8500/3
C1134719|T191|PT|MTHU014771|ICPC2ICD10ENG|carcinoma; infiltrating ductular, unspecified site|8500/3
C1134719|T191|PT|MTHU024095|ICPC2ICD10ENG|ductal; carcinoma, infiltrating, unspecified site|8500/3
C1134719|T191|PT|MTHU024097|ICPC2ICD10ENG|ductular; carcinoma, infiltrating, unspecified site|8500/3
C1134719|T191|PT|MTHU039173|ICPC2ICD10ENG|infiltrating; ductal adenocarcinoma, unspecified site|8500/3
C1134719|T191|PT|MTHU039175|ICPC2ICD10ENG|infiltrating; ductal carcinoma, unspecified site|8500/3
C1134719|T191|PT|MTHU039176|ICPC2ICD10ENG|infiltrating; ductular carcinoma, unspecified site|8500/3
C1134719|T191|LLT|10006235|MDR|Breast ductal cancer infiltrating|8500/3
C1134719|T191|LLT|10006236|MDR|Breast ductal cancer invasive|8500/3
C1134719|T191|LLT|10021944|MDR|Infiltrating ductal breast cancer|8500/3
C1134719|T191|LLT|10022882|MDR|Invasive ductal breast cancer|8500/3
C1134719|T191|LLT|10073095|MDR|Invasive ductal breast carcinoma|8500/3
C1134719|T191|PT|10073095|MDR|Invasive ductal breast carcinoma|8500/3
C1134719|T191|PT|232310|MEDCIN|infiltrating ductal carcinoma of breast|8500/3
C1134719|T191|MH|D018270|MSH|Carcinoma, Ductal, Breast|8500/3
C1134719|T191|ET|D018270|MSH|Carcinoma, Infiltrating Duct|8500/3
C1134719|T191|ET|D018270|MSH|Carcinoma, Invasive Ductal, Breast|8500/3
C1134719|T191|PM|D018270|MSH|Carcinomas, Infiltrating Duct|8500/3
C1134719|T191|ET|D018270|MSH|Invasive Ductal Carcinoma, Breast|8500/3
C1412014|T191|PN|NOCODE|MTH|Infiltrating duct carcinoma|8500/3
C1134719|T191|PN|NOCODE|MTH|Invasive Ductal Breast Carcinoma|8500/3
C1301194|T191|SY|C5904|NCI|Carcinoma of Salivary Duct|8500/3
C1301194|T191|SY|C5904|NCI|Carcinoma of the Salivary Duct|8500/3
C1301194|T191|SY|C5904|NCI|High Grade Salivary Duct Carcinoma|8500/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Adenocarcinoma|8500/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Breast Carcinoma|8500/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Carcinoma|8500/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Carcinoma of Breast|8500/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Carcinoma of the Breast|8500/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Adenocarcinoma|8500/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Breast Carcinoma|8500/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma|8500/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma of Breast|8500/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma of the Breast|8500/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma, No Specific Type|8500/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma, NOS|8500/3
C1134719|T191|PT|C4194|NCI|Invasive Ductal Carcinoma, Not Otherwise Specified|8500/3
C1134719|T191|SY|TCGA|NCI|Invasive Ductal Carcinoma, Not Otherwise Specified|8500/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma, NST|8500/3
C1301194|T191|PT|C5904|NCI|Salivary Duct Carcinoma|8500/3
C1134719|T191|DN|C4194|NCI_CTRP|Invasive Ductal Carcinoma, NOS|8500/3
C1134719|T191|PT|CDR0000045099|NCI_NCI-GLOSS|infiltrating ductal carcinoma|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|ductal invasive breast carcinoma|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Adenocarcinoma|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Breast Carcinoma|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Carcinoma|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Carcinoma of Breast|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Carcinoma of the Breast|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Adenocarcinoma|8500/3
C1134719|T191|PT|CDR0000039843|PDQ|invasive ductal breast carcinoma|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma of Breast|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma of the Breast|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma, No Specific Type|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma, NOS|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma, Not Otherwise Specified|8500/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma, NST|8500/3
C1412014|T191|AB|BB91.|RCD|Infiltrating duct adenoca|8500/3
C1412014|T191|SY|BB91.|RCD|Infiltrating duct adenocarcinoma|8500/3
C1412014|T191|PT|BB91.|RCD|Infiltrating duct carcinoma|8500/3
C1134719|T191|AB|BB9G.|RCD|Infiltrating ductular ca|8500/3
C1134719|T191|PT|BB9G.|RCD|Infiltrating ductular carcinoma|8500/3
C3839330|T191|PT|703570003|SNOMEDCT_US|Adenocarcinoma of mammary gland type|8500/3
C1412014|T191|SY|82711006|SNOMEDCT_US|Infiltrating duct adenocarcinoma|8500/3
C1412014|T191|PT|82711006|SNOMEDCT_US|Infiltrating duct carcinoma|8500/3
C1134719|T191|PT|408643008|SNOMEDCT_US|Infiltrating duct carcinoma of breast|8500/3
C1134719|T191|SY|408643008|SNOMEDCT_US|Infiltrating ductal carcinoma of breast|8500/3
C1134719|T191|PT|58477004|SNOMEDCT_US|Infiltrating ductular carcinoma|8500/3
C1412014|T191|SY|82711006|SNOMEDCT_US|Invasive breast carcinoma of no special type|8500/3
C1134719|T191|SY|408643008|SNOMEDCT_US|Invasive duct carcinoma of breast|8500/3
C1134719|T191|SY|408643008|SNOMEDCT_US|Invasive ductal carcinoma of breast|8500/3
C1298749|T191|PT|373395001|SNOMEDCT_US|Invasive ductal carcinoma with an extensive intraductal component|8500/3
C1301194|T191|PT|397082006|SNOMEDCT_US|Salivary duct carcinoma|8500/3
C1334002|T191|LLT|10066275|MDR|Comedocarcinoma of breast|8501/2
C1334002|T191|PT|232311|MEDCIN|comedocarcinoma of breast|8501/2
C1334002|T191|PN|NOCODE|MTH|High Grade Ductal Breast Carcinoma In Situ|8501/2
C1334002|T191|SY|C7949|NCI|Breast Comedocarcinoma|8501/2
C1334002|T191|SY|C7949|NCI|DCIS Grade 3|8501/2
C1334002|T191|AB|C7949|NCI|DIN 3|8501/2
C1334002|T191|SY|C7949|NCI|Ductal Intraepithelial Neoplasia, Grade 3|8501/2
C1334002|T191|PT|C7949|NCI|High Grade Ductal Breast Carcinoma In Situ|8501/2
C1334002|T191|SY|C7949|NCI|High-Grade DCIS of Breast|8501/2
C1334002|T191|SY|C7949|NCI|High-Grade DCIS of the Breast|8501/2
C1334002|T191|SY|C7949|NCI|High-Grade Ductal Carcinoma In Situ of Breast|8501/2
C1334002|T191|DN|C7949|NCI_CTRP|High Grade Ductal Breast Carcinoma In Situ|8501/2
C1334002|T191|PT|CDR0000044330|NCI_NCI-GLOSS|comedo carcinoma|8501/2
C1334002|T191|SY|CDR0000039844|PDQ|Breast Comedocarcinoma|8501/2
C1334002|T191|PT|CDR0000039844|PDQ|comedo ductal breast carcinoma|8501/2
C1334002|T191|SY|CDR0000039844|PDQ|DCIS Grade 3|8501/2
C1334002|T191|AB|CDR0000039844|PDQ|DIN 3|8501/2
C1334002|T191|SY|CDR0000039844|PDQ|ductal comedo breast carcinoma|8501/2
C1334002|T191|SY|CDR0000039844|PDQ|Ductal Intraepithelial Neoplasia, Grade 3|8501/2
C1334002|T191|SY|CDR0000039844|PDQ|High Grade Ductal Breast Carcinoma In Situ|8501/2
C1334002|T191|SY|CDR0000039844|PDQ|High-Grade DCIS of Breast|8501/2
C1334002|T191|SY|CDR0000039844|PDQ|High-Grade DCIS of the Breast|8501/2
C1334002|T191|SY|CDR0000039844|PDQ|High-Grade Ductal Carcinoma In Situ of Breast|8501/2
C0334369|T191|OA|BB92.|RCD|Non-infiltrating comedoca|8501/2
C0334369|T191|OP|BB92.|RCD|Non-infiltrating comedocarcinoma|8501/2
C0334369|T191|PT|78197004|SNOMEDCT_US|Comedocarcinoma, noninfiltrating|8501/2
C0334369|T191|SY|78197004|SNOMEDCT_US|DCIS, comedo type|8501/2
C1334002|T191|SY|86616005|SNOMEDCT_US|DIN 3|8501/2
C0334369|T191|SY|78197004|SNOMEDCT_US|Ductal carcinoma in situ, comedo type|8501/2
C1334002|T191|SY|86616005|SNOMEDCT_US|Ductal intraepithelial neoplasia 3|8501/2
C0334369|T191|SY|78197004|SNOMEDCT_US|Non-infiltrating comedocarcinoma|8501/2
C0334370|T191|PN|NOCODE|MTH|Comedocarcinoma|8501/3
C0334370|T191|PT|C4188|NCI|Comedocarcinoma|8501/3
C0334370|T191|PT|C4188|NCI_CPTAC|Comedocarcinoma|8501/3
C0334370|T191|PT|Xa98u|RCD|Comedocarcinoma|8501/3
C0334370|T191|OP|BB93.|RCDSY|Comedocarcinoma NOS|8501/3
C0334370|T191|OAP|36425007|SNOMEDCT_US|Comedocarcinoma|8501/3
C4302718|T191|SY|722237009|SNOMEDCT_US|Comedocarcinoma, no ICD-O subtype|8501/3
C4302718|T191|PT|722237009|SNOMEDCT_US|Comedocarcinoma, no International Classification of Diseases for Oncology subtype|8501/3
C0334370|T191|IS|36425007|SNOMEDCT_US|Comedocarcinoma, NOS|8501/3
C0334371|T191|PT|232314|MEDCIN|hypersecretory cystic carcinoma of breast|8502/3
C0334371|T191|PT|232312|MEDCIN|secretory carcinoma of breast|8502/3
C0334371|T191|NM|C537535|MSH|Secretory breast carcinoma|8502/3
C0334371|T191|SY|C4189|NCI|Cystic Hypersecretory Breast Carcinoma|8502/3
C0334371|T191|SY|C4189|NCI|Cystic Hypersecretory Carcinoma of Breast|8502/3
C0334371|T191|SY|C4189|NCI|Cystic Hypersecretory Carcinoma of the Breast|8502/3
C0334371|T191|SY|C4189|NCI|Infiltrating Cystic Hypersecretory Duct Breast Carcinoma|8502/3
C0334371|T191|SY|C4189|NCI|Invasive Cystic Hypersecretory Duct Breast Carcinoma|8502/3
C0334371|T191|SY|C4189|NCI|Juvenile Breast Carcinoma|8502/3
C0334371|T191|SY|C4189|NCI|Juvenile Carcinoma of Breast|8502/3
C0334371|T191|SY|C4189|NCI|Juvenile Carcinoma of the Breast|8502/3
C0334371|T191|SY|C4189|NCI|Juvenile Secretory Breast Carcinoma|8502/3
C0334371|T191|SY|C4189|NCI|Juvenile Secretory Carcinoma of Breast|8502/3
C0334371|T191|SY|C4189|NCI|Juvenile Secretory Carcinoma of the Breast|8502/3
C0334371|T191|PT|C4189|NCI|Secretory Breast Carcinoma|8502/3
C0334371|T191|SY|C4189|NCI|Secretory Carcinoma|8502/3
C0334371|T191|SY|C4189|NCI|Secretory Carcinoma of Breast|8502/3
C0334371|T191|SY|C4189|NCI|Secretory Carcinoma of the Breast|8502/3
C0334371|T191|AB|BB94.|RCD|Juvenile carcinoma of breast|8502/3
C0334371|T191|PT|BB94.|RCD|Juvenile carcinoma of the breast|8502/3
C0334371|T191|AB|BB94.|RCD|Secretory carcinoma of breast|8502/3
C0334371|T191|SY|BB94.|RCD|Secretory carcinoma of the breast|8502/3
C0334371|T191|PT|41919003|SNOMEDCT_US|Juvenile carcinoma of the breast|8502/3
C0334371|T191|SY|41919003|SNOMEDCT_US|Secretory carcinoma of the breast|8502/3
C0206713|T191|SY|0000021040|CHV|duct adenoma|8503/0
C0206713|T191|SY|0000021040|CHV|ductal papilloma|8503/0
C0206713|T191|SY|0000021040|CHV|ductal papillomas|8503/0
C0206713|T191|PT|0000021040|CHV|intraductal papilloma|8503/0
C0206713|T191|SY|0000021040|CHV|intraductal papillomas|8503/0
C0206713|T191|SY|0000021040|CHV|papilloma intraductal|8503/0
C0206713|T191|PT|NOCODE|COSTAR|Intraductal Papilloma|8503/0
C3160815|T191|LLT|10070999|MDR|Intraductal papillary mucinous neoplasm|8503/0
C3160815|T191|PT|10070999|MDR|Intraductal papillary mucinous neoplasm|8503/0
C0206713|T191|PM|D018300|MSH|Intraductal Papilloma|8503/0
C0206713|T191|PM|D018300|MSH|Intraductal Papillomas|8503/0
C2987189|T191|ET|D000077779|MSH|Intraductal Tubulopapillary Neoplasm, Pancreatic|8503/0
C2987189|T191|PEP|D000077779|MSH|Pancreatic Intraductal Tubulopapillary Neoplasm|8503/0
C0206713|T191|MH|D018300|MSH|Papilloma, Intraductal|8503/0
C0206713|T191|PM|D018300|MSH|Papillomas, Intraductal|8503/0
C1879344|T191|PT|C6881|NCI|Bile Duct Papillary Neoplasm|8503/0
C3273049|T191|PT|C96807|NCI|Bile Duct Papillary Neoplasm with Low Grade Intraepithelial Neoplasia|8503/0
C1879344|T191|SY|C6881|NCI|Bile Duct Papillomatosis|8503/0
C1879344|T191|SY|C6881|NCI|Biliary Papillomatosis|8503/0
C0206713|T191|OP|C3785|NCI|Duct Adenoma|8503/0
C0206713|T191|SY|C3785|NCI|Ductal Papilloma|8503/0
C3273094|T191|PT|C96878|NCI|Gallbladder Papillary Neoplasm with Intermediate Grade Intraepithelial Neoplasia|8503/0
C3273093|T191|PT|C96877|NCI|Gallbladder Papillary Neoplasm with Low Grade Intraepithelial Neoplasia|8503/0
C3273094|T191|SY|C96878|NCI|Intracystic Papillary Neoplasm with Intermediate Grade Intraepithelial Neoplasia|8503/0
C3273093|T191|SY|C96877|NCI|Intracystic Papillary Neoplasm with Low Grade Intraepithelial Neoplasia|8503/0
C1879344|T191|SY|C6881|NCI|Intraductal Papillary Neoplasm|8503/0
C3273049|T191|SY|C96807|NCI|Intraductal Papillary Neoplasm with Low Grade Intraepithelial Neoplasia|8503/0
C0206713|T191|PT|C3785|NCI|Intraductal Papilloma|8503/0
C1879344|T191|AB|C6881|NCI|IPN|8503/0
C2987189|T191|AB|C95506|NCI|ITPN|8503/0
C2987189|T191|SY|C95506|NCI|Pancreatic Intraductal Tubular Neoplasm|8503/0
C2987189|T191|PT|C95506|NCI|Pancreatic Intraductal Tubulopapillary Neoplasm|8503/0
C2987189|T191|SY|C95506|NCI|Pancreatic ITPN|8503/0
C0206713|T191|PT|CDR0000430864|NCI_NCI-GLOSS|intraductal papilloma|8503/0
C0206713|T191|SY|BB95.|RCD|Duct adenoma|8503/0
C0206713|T191|SY|BB95.|RCD|Ductal papilloma|8503/0
C0206713|T191|PT|BB95.|RCD|Intraductal papilloma|8503/0
C1879344|T191|SY|128663007|SNOMEDCT_US|Biliary papillomatosis|8503/0
C0206713|T191|SY|5244003|SNOMEDCT_US|Duct adenoma|8503/0
C0206713|T191|IS|5244003|SNOMEDCT_US|Duct adenoma, NOS|8503/0
C0206713|T191|SY|5244003|SNOMEDCT_US|Ductal papilloma|8503/0
C3273093|T191|PT|734135002|SNOMEDCT_US|Intracystic papillary neoplasm with low grade intraepithelial neoplasia|8503/0
C3160815|T191|PT|726097000|SNOMEDCT_US|Intraductal papillary mucinous neoplasm|8503/0
C3273049|T191|PT|734091005|SNOMEDCT_US|Intraductal papillary neoplasm with low-grade intraepithelial neoplasia|8503/0
C0206713|T191|PT|5244003|SNOMEDCT_US|Intraductal papilloma|8503/0
C3840150|T191|PT|703575008|SNOMEDCT_US|Intraductal papilloma with atypical ductal hyperplasia|8503/0
C4518202|T191|PT|733846005|SNOMEDCT_US|Inverted ductal papilloma|8503/0
C0334372|T191|PT|MTHU003404|ICPC2ICD10ENG|adenocarcinoma; intraductal, papillary, breast|8503/2
C0334372|T191|PT|MTHU003415|ICPC2ICD10ENG|adenocarcinoma; papillary, intraductal, breast|8503/2
C0334372|T191|PT|MTHU047386|ICPC2ICD10ENG|breast; carcinoma, intraductal papillary|8503/2
C0334372|T191|PT|MTHU047430|ICPC2ICD10ENG|breast; intraductal papillary carcinoma|8503/2
C0334372|T191|PT|MTHU014778|ICPC2ICD10ENG|carcinoma; intraductal, papillary, breast|8503/2
C0334372|T191|PT|MTHU040060|ICPC2ICD10ENG|intraductal; carcinoma, papillary, breast|8503/2
C0334372|T191|PT|MTHU057277|ICPC2ICD10ENG|papillary; adenocarcinoma, intraductal, breast|8503/2
C2987189|T191|ET|D000077779|MSH|Intraductal Tubulopapillary Neoplasm, Pancreatic|8503/2
C2987189|T191|PEP|D000077779|MSH|Pancreatic Intraductal Tubulopapillary Neoplasm|8503/2
C3273051|T191|PT|C96809|NCI|Bile Duct Papillary Neoplasm with High Grade Intraepithelial Neoplasia|8503/2
C3273095|T191|PT|C96879|NCI|Gallbladder Papillary Neoplasm with High Grade Intraepithelial Neoplasia|8503/2
C3273095|T191|SY|C96879|NCI|Intracystic Papillary Neoplasm with High Grade Intraepithelial Neoplasia|8503/2
C0334372|T191|SY|C4190|NCI|Intraductal Papillary Adenocarcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Intraductal Papillary Breast Adenocarcinoma|8503/2
C0334372|T191|PT|C4190|NCI|Intraductal Papillary Breast Carcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Intraductal Papillary Carcinoma|8503/2
C3273051|T191|SY|C96809|NCI|Intraductal Papillary Neoplasm with High Grade Intraepithelial Neoplasia|8503/2
C2987189|T191|AB|C95506|NCI|ITPN|8503/2
C0334372|T191|SY|C4190|NCI|Non-Infiltrating Intraductal Papillary Adenocarcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Non-Infiltrating Intraductal Papillary Carcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Non-Infiltrating Papillary Breast Adenocarcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Non-Infiltrating Papillary Breast Carcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Non-Invasive Intraductal Papillary Adenocarcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Non-Invasive Intraductal Papillary Carcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Non-Invasive Papillary Breast Adenocarcinoma|8503/2
C0334372|T191|SY|C4190|NCI|Non-Invasive Papillary Breast Carcinoma|8503/2
C2987189|T191|SY|C95506|NCI|Pancreatic Intraductal Tubular Neoplasm|8503/2
C2987189|T191|PT|C95506|NCI|Pancreatic Intraductal Tubulopapillary Neoplasm|8503/2
C2987189|T191|SY|C95506|NCI|Pancreatic ITPN|8503/2
C0334372|T191|AB|BB96.|RCD|Intraductal papillary adenoca|8503/2
C0334372|T191|SY|BB96.|RCD|Intraductal papillary adenocarcinoma|8503/2
C0334372|T191|AB|BB96.|RCD|Intraductal papillary ca|8503/2
C0334372|T191|SY|BB96.|RCD|Intraductal papillary carcinoma|8503/2
C0334372|T191|AB|BB96.|RCD|Non-infil intraduc pap adenoca|8503/2
C0334372|T191|AB|BB96.|RCD|Non-infilt intraduct papill ca|8503/2
C0334372|T191|PT|BB96.|RCD|Non-infiltrating intraductal papillary adenocarcinoma|8503/2
C0334372|T191|SY|BB96.|RCD|Non-infiltrating intraductal papillary carcinoma|8503/2
C0334372|T191|SY|30566004|SNOMEDCT_US|DCIS, papillary|8503/2
C0334372|T191|SY|30566004|SNOMEDCT_US|Ductal carcinoma in situ, papillary|8503/2
C0334372|T191|SY|30566004|SNOMEDCT_US|Intraductal papillary adenocarcinoma|8503/2
C0334372|T191|IS|30566004|SNOMEDCT_US|Intraductal papillary adenocarcinoma, NOS|8503/2
C0334372|T191|SY|30566004|SNOMEDCT_US|Intraductal papillary carcinoma|8503/2
C0334372|T191|IS|30566004|SNOMEDCT_US|Intraductal papillary carcinoma, NOS|8503/2
C3273051|T191|PT|734133009|SNOMEDCT_US|Intraductal papillary neoplasm with high grade intraepithelial neoplasia|8503/2
C3839576|T191|SY|703576009|SNOMEDCT_US|Intraductal papilloma with DCIS|8503/2
C3839576|T191|PT|703576009|SNOMEDCT_US|Intraductal papilloma with ductal carcinoma in situ|8503/2
C0334372|T191|SY|30566004|SNOMEDCT_US|Non-infiltrating intraductal papillary adenocarcinoma|8503/2
C0334372|T191|SY|30566004|SNOMEDCT_US|Non-infiltrating intraductal papillary carcinoma|8503/2
C0334372|T191|PT|30566004|SNOMEDCT_US|Noninfiltrating intraductal papillary adenocarcinoma|8503/2
C0334372|T191|SY|30566004|SNOMEDCT_US|Noninfiltrating intraductal papillary carcinoma|8503/2
C1333753|T191|LLT|10073079|MDR|Gallbladder papillary adenocarcinoma|8503/3
C3812899|T191|LLT|10066207|MDR|Papillary breast carcinoma|8503/3
C1333753|T191|PT|39460|MEDCIN|papillary adenocarcinoma of gallbladder|8503/3
C3812899|T191|PT|232289|MEDCIN|papillary carcinoma of breast|8503/3
C1333753|T191|PT|218093|MEDCIN|papillary carcinoma of gallbladder|8503/3
C3273052|T191|PN|NOCODE|MTH|Bile Duct Papillary Neoplasm with an Associated Invasive Carcinoma|8503/3
C3273052|T191|SY|C96810|NCI|Bile Duct Papillary Adenocarcinoma|8503/3
C3273052|T191|PT|C96810|NCI|Bile Duct Papillary Neoplasm with an Associated Invasive Carcinoma|8503/3
C1333753|T191|PT|C5743|NCI|Gallbladder Papillary Neoplasm with an Associated Invasive Carcinoma|8503/3
C1333753|T191|SY|C5743|NCI|Intracystic Papillary Neoplasm with an Associated Invasive Carcinoma|8503/3
C0334373|T191|PT|C7439|NCI|Intraductal Papillary Adenocarcinoma with Invasion|8503/3
C3273052|T191|SY|C96810|NCI|Intraductal Papillary Neoplasm with an Associated Invasive Carcinoma|8503/3
C3812899|T191|PT|C9134|NCI|Papillary Breast Carcinoma|8503/3
C3812899|T191|SY|C9134|NCI|Papillary Carcinoma of Breast|8503/3
C1333753|T191|SY|C5743|NCI|Papillary Carcinoma of Gallbladder|8503/3
C3812899|T191|SY|C9134|NCI|Papillary Carcinoma of the Breast|8503/3
C1333753|T191|SY|C5743|NCI|Papillary Carcinoma of the Gallbladder|8503/3
C1333753|T191|DN|C5743|NCI_CTRP|Gallbladder Papillary Neoplasm with an Associated Invasive Cancer|8503/3
C3812899|T191|DN|C9134|NCI_CTRP|Papillary Breast Cancer|8503/3
C3812899|T191|SY|CDR0000039845|PDQ|ductal papillary breast carcinoma|8503/3
C3812899|T191|SY|CDR0000039845|PDQ|Papillary Breast Carcinoma|8503/3
C3812899|T191|SY|CDR0000039845|PDQ|Papillary Carcinoma of Breast|8503/3
C3812899|T191|SY|CDR0000039845|PDQ|Papillary Carcinoma of the Breast|8503/3
C3812899|T191|PT|CDR0000039845|PDQ|papillary ductal breast carcinoma|8503/3
C0334373|T191|AB|X77nu|RCD|Intraduc papill adenoca+invas|8503/3
C0334373|T191|PT|X77nu|RCD|Intraductal papillary adenocarcinoma with invasion|8503/3
C0334373|T191|AB|X77nu|RCDSY|Intrad papil adenoc+invason|8503/3
C0334373|T191|OAP|189706007|SNOMEDCT_US|Intraductal papillary adenocarcinoma with invasion|8503/3
C0334373|T191|OF|189706007|SNOMEDCT_US|Intraductal papillary adenocarcinoma with invasion|8503/3
C0334373|T191|PT|64524002|SNOMEDCT_US|Intraductal papillary adenocarcinoma with invasion|8503/3
C4518374|T191|PT|734075007|SNOMEDCT_US|Intraductal papillary neoplasm with invasive carcinoma|8503/3
C3812899|T191|PT|703577000|SNOMEDCT_US|Papillary carcinoma of the breast|8503/3
C0334374|T191|SY|C4191|NCI|Intracystic Papillary Adenoma|8504/0
C0334374|T191|PT|C4191|NCI|Intracystic Papilloma|8504/0
C0334374|T191|PT|BB97.|RCD|Intracystic papillary adenoma|8504/0
C0334374|T191|SY|BB97.|RCD|Intracystic papilloma|8504/0
C0334374|T191|PT|47488001|SNOMEDCT_US|Intracystic papillary adenoma|8504/0
C0334374|T191|SY|47488001|SNOMEDCT_US|Intracystic papilloma|8504/0
C0334376|T191|PT|232313|MEDCIN|intracystic carcinoma of breast|8504/2
C1266053|T191|PN|NOCODE|MTH|Encapsulated papillary carcinoma|8504/2
C0334376|T191|PN|NOCODE|MTH|Intracystic Papillary Breast Carcinoma|8504/2
C0334375|T191|PN|NOCODE|MTH|Noninfiltrating intracystic carcinoma|8504/2
C0334376|T191|SY|C7645|NCI|Intracystic Breast Carcinoma|8504/2
C0334376|T191|SY|C7645|NCI|Intracystic Papillary Adenocarcinoma|8504/2
C0334376|T191|PT|C7645|NCI|Intracystic Papillary Breast Carcinoma|8504/2
C0334376|T191|SY|C7645|NCI|Noninfiltrating Intracystic Breast Carcinoma|8504/2
C0334376|T191|PT|X77nv|RCD|Intracystic carcinoma|8504/2
C0334376|T191|AB|X77nv|RCD|Intracystic papillary adenoca|8504/2
C0334376|T191|SY|X77nv|RCD|Intracystic papillary adenocarcinoma|8504/2
C0334375|T191|AB|BB98.|RCD|Non-infiltrat intracystic ca|8504/2
C0334375|T191|PT|BB98.|RCD|Non-infiltrating intracystic carcinoma|8504/2
C0334376|T191|OP|BB9M.|RCDSY|Intracystic carcinoma NOS|8504/2
C1266053|T191|PT|703545003|SNOMEDCT_US|Encapsulated papillary carcinoma|8504/2
C1266053|T191|SY|703545003|SNOMEDCT_US|Encysted papillary carcinoma|8504/2
C0334376|T191|OAP|23746000|SNOMEDCT_US|Intracystic carcinoma|8504/2
C0334376|T191|IS|23746000|SNOMEDCT_US|Intracystic carcinoma, NOS|8504/2
C0334376|T191|OAS|23746000|SNOMEDCT_US|Intracystic papillary adenocarcinoma|8504/2
C1266053|T191|SY|703545003|SNOMEDCT_US|Intracystic papillary adenocarcinoma|8504/2
C1266053|T191|SY|703545003|SNOMEDCT_US|Intracystic papillary carcinoma|8504/2
C1266053|T191|SY|703545003|SNOMEDCT_US|Non-infiltrating intracystic carcinoma|8504/2
C0334375|T191|OAS|89277004|SNOMEDCT_US|Non-infiltrating intracystic carcinoma|8504/2
C0334375|T191|OAP|89277004|SNOMEDCT_US|Noninfiltrating intracystic carcinoma|8504/2
C1266053|T191|SY|703545003|SNOMEDCT_US|Noninfiltrating intracystic carcinoma|8504/2
C1266053|T191|OAP|128676001|SNOMEDCT_US|Papillary carcinoma, encapsulated|8504/2
C0334376|T191|PT|232313|MEDCIN|intracystic carcinoma of breast|8504/3
C0334376|T191|PN|NOCODE|MTH|Intracystic Papillary Breast Carcinoma|8504/3
C0334376|T191|SY|C7645|NCI|Intracystic Breast Carcinoma|8504/3
C0334376|T191|SY|C7645|NCI|Intracystic Papillary Adenocarcinoma|8504/3
C0334376|T191|PT|C7645|NCI|Intracystic Papillary Breast Carcinoma|8504/3
C0334376|T191|SY|C7645|NCI|Noninfiltrating Intracystic Breast Carcinoma|8504/3
C0334376|T191|PT|X77nv|RCD|Intracystic carcinoma|8504/3
C0334376|T191|AB|X77nv|RCD|Intracystic papillary adenoca|8504/3
C0334376|T191|SY|X77nv|RCD|Intracystic papillary adenocarcinoma|8504/3
C0334376|T191|OP|BB9M.|RCDSY|Intracystic carcinoma NOS|8504/3
C3838872|T191|PT|703547006|SNOMEDCT_US|Encapsulated papillary carcinoma with invasion|8504/3
C3838872|T191|SY|703547006|SNOMEDCT_US|Encysted papillary carcinoma with invasion|8504/3
C0334376|T191|OAP|23746000|SNOMEDCT_US|Intracystic carcinoma|8504/3
C0334376|T191|IS|23746000|SNOMEDCT_US|Intracystic carcinoma, NOS|8504/3
C0334376|T191|OAS|23746000|SNOMEDCT_US|Intracystic papillary adenocarcinoma|8504/3
C3838872|T191|SY|703547006|SNOMEDCT_US|Intracystic papillary adenocarcinoma with invasion|8504/3
C3838872|T191|SY|703547006|SNOMEDCT_US|Intracystic papillary carcinoma with invasion|8504/3
C0334377|T191|PT|C7363|NCI|Intraductal Papillomatosis|8505/0
C0334377|T191|PT|Xa98v|RCD|Intraductal papillomatosis|8505/0
C0334377|T191|OA|BB99.|RCDSY|Intraduct.papillomatos.NOS|8505/0
C0334377|T191|OP|BB99.|RCDSY|Intraductal papillomatosis NOS|8505/0
C0334377|T191|PT|32296002|SNOMEDCT_US|Intraductal papillomatosis|8505/0
C0334377|T191|IS|32296002|SNOMEDCT_US|Intraductal papillomatosis, NOS|8505/0
C0334378|T191|SY|0000029967|CHV|adenoma of the nipple|8506/0
C0334378|T191|SY|0000029967|CHV|adenomas nipple|8506/0
C0334378|T191|PT|0000029967|CHV|nipple adenoma|8506/0
C0334378|T191|PT|MTHU003525|ICPC2ICD10ENG|adenoma; nipple|8506/0
C0334378|T191|PT|MTHU073741|ICPC2ICD10ENG|nipple; adenoma|8506/0
C0334378|T191|PCE|C000626393|MSH|Nipple Adenoma|8506/0
C0334378|T191|SY|C4192|NCI|Adenoma of Nipple|8506/0
C0334378|T191|SY|C4192|NCI|Adenoma of the Nipple|8506/0
C0334378|T191|PT|C4192|NCI|Nipple Adenoma|8506/0
C0334378|T191|SY|C4192|NCI|Papillomatosis, Subareolar Duct|8506/0
C0334378|T191|SY|C4192|NCI|Subareolar Duct Papillomatosis|8506/0
C0334378|T191|PT|Xa98w|RCD|Adenoma of nipple|8506/0
C0334378|T191|IS|BB9A.|RCD|Subareolar duct papillomatosis|8506/0
C0334378|T191|OA|BB9A.|RCDSY|Subareolar duct papillomat.|8506/0
C0334378|T191|PT|302829009|SNOMEDCT_US|Adenoma of nipple|8506/0
C0334378|T191|PT|65787003|SNOMEDCT_US|Adenoma of the nipple|8506/0
C0334378|T191|SY|65787003|SNOMEDCT_US|Subareolar duct papillomatosis|8506/0
C1334249|T191|PT|232266|MEDCIN|intraductal micropapillary carcinoma of breast|8507/2
C1266080|T191|PN|NOCODE|MTH|Intraductal micropapillary carcinoma|8507/2
C1334249|T191|PT|C5139|NCI|Intraductal Micropapillary Breast Carcinoma|8507/2
C1334249|T191|SY|TCGA|NCI|Intraductal Micropapillary Breast Carcinoma|8507/2
C1334249|T191|SY|C5139|NCI|Micropapillary DCIS of Breast|8507/2
C1334249|T191|SY|C5139|NCI|Micropapillary DCIS of the Breast|8507/2
C1334249|T191|SY|C5139|NCI|Micropapillary Ductal Breast Carcinoma in situ|8507/2
C1334249|T191|SY|C5139|NCI|Micropapillary Ductal Carcinoma in situ of Breast|8507/2
C1334249|T191|SY|C5139|NCI|Micropapillary Ductal Carcinoma in situ of the Breast|8507/2
C1334249|T191|SY|C5139|NCI|Non-Infiltrating Micropapillary Breast Carcinoma|8507/2
C1334249|T191|SY|C5139|NCI|Non-Infiltrating Micropapillary Carcinoma of Breast|8507/2
C1334249|T191|SY|C5139|NCI|Non-Infiltrating Micropapillary Carcinoma of the Breast|8507/2
C1334249|T191|SY|C5139|NCI|Non-Infiltrating Micropapillary Ductal Breast Carcinoma|8507/2
C1334249|T191|SY|C5139|NCI|Non-Infiltrating Micropapillary Ductal Carcinoma of Breast|8507/2
C1334249|T191|SY|C5139|NCI|Non-Infiltrating Micropapillary Ductal Carcinoma of the Breast|8507/2
C1334249|T191|SY|C5139|NCI|Non-Invasive Micropapillary Breast Carcinoma|8507/2
C1334249|T191|SY|C5139|NCI|Non-Invasive Micropapillary Carcinoma of Breast|8507/2
C1334249|T191|SY|C5139|NCI|Non-Invasive Micropapillary Carcinoma of the Breast|8507/2
C1334249|T191|SY|C5139|NCI|Non-Invasive Micropapillary Ductal Breast Carcinoma|8507/2
C1334249|T191|SY|C5139|NCI|Non-Invasive Micropapillary Ductal Carcinoma of Breast|8507/2
C1334249|T191|SY|C5139|NCI|Non-Invasive Micropapillary Ductal Carcinoma of the Breast|8507/2
C1266080|T191|SY|128696009|SNOMEDCT_US|Ductal carcinoma in situ, micropapillary|8507/2
C1266080|T191|IS|128696009|SNOMEDCT_US|Intraductal carcinoma, clinging|8507/2
C1266080|T191|SY|128696009|SNOMEDCT_US|Intraductal carcinoma, clinging, high grade|8507/2
C1266080|T191|PT|128696009|SNOMEDCT_US|Intraductal micropapillary carcinoma|8507/2
C1334280|T191|LLT|10073098|MDR|Invasive papillary breast carcinoma|8507/3
C1334280|T191|PT|10073098|MDR|Invasive papillary breast carcinoma|8507/3
C3838947|T191|SY|C36084|NCI|Infiltrating Micropapillary Breast Carcinoma|8507/3
C1334280|T191|SY|C36085|NCI|Infiltrating Papillary Breast Carcinoma|8507/3
C3838947|T191|PT|C36084|NCI|Invasive Micropapillary Breast Carcinoma|8507/3
C1334280|T191|PT|C36085|NCI|Invasive Papillary Breast Carcinoma|8507/3
C3838947|T191|PT|703578005|SNOMEDCT_US|Invasive micropapillary carcinoma of breast|8507/3
C3839300|T191|PT|703573001|SNOMEDCT_US|Cystic hypersecretory carcinoma, intraductal|8508/2
C0334371|T191|PT|232314|MEDCIN|hypersecretory cystic carcinoma of breast|8508/3
C0334371|T191|PT|232312|MEDCIN|secretory carcinoma of breast|8508/3
C0334371|T191|NM|C537535|MSH|Secretory breast carcinoma|8508/3
C0334371|T191|SY|C4189|NCI|Cystic Hypersecretory Breast Carcinoma|8508/3
C0334371|T191|SY|C4189|NCI|Cystic Hypersecretory Carcinoma of Breast|8508/3
C0334371|T191|SY|C4189|NCI|Cystic Hypersecretory Carcinoma of the Breast|8508/3
C0334371|T191|SY|C4189|NCI|Infiltrating Cystic Hypersecretory Duct Breast Carcinoma|8508/3
C0334371|T191|SY|C4189|NCI|Invasive Cystic Hypersecretory Duct Breast Carcinoma|8508/3
C0334371|T191|SY|C4189|NCI|Juvenile Breast Carcinoma|8508/3
C0334371|T191|SY|C4189|NCI|Juvenile Carcinoma of Breast|8508/3
C0334371|T191|SY|C4189|NCI|Juvenile Carcinoma of the Breast|8508/3
C0334371|T191|SY|C4189|NCI|Juvenile Secretory Breast Carcinoma|8508/3
C0334371|T191|SY|C4189|NCI|Juvenile Secretory Carcinoma of Breast|8508/3
C0334371|T191|SY|C4189|NCI|Juvenile Secretory Carcinoma of the Breast|8508/3
C0334371|T191|PT|C4189|NCI|Secretory Breast Carcinoma|8508/3
C0334371|T191|SY|C4189|NCI|Secretory Carcinoma|8508/3
C0334371|T191|SY|C4189|NCI|Secretory Carcinoma of Breast|8508/3
C0334371|T191|SY|C4189|NCI|Secretory Carcinoma of the Breast|8508/3
C0334371|T191|AB|BB94.|RCD|Juvenile carcinoma of breast|8508/3
C0334371|T191|PT|BB94.|RCD|Juvenile carcinoma of the breast|8508/3
C0334371|T191|AB|BB94.|RCD|Secretory carcinoma of breast|8508/3
C0334371|T191|SY|BB94.|RCD|Secretory carcinoma of the breast|8508/3
C1266081|T191|PT|128697000|SNOMEDCT_US|Cystic hypersecretory carcinoma|8508/3
C0334371|T191|PT|41919003|SNOMEDCT_US|Juvenile carcinoma of the breast|8508/3
C0334371|T191|SY|41919003|SNOMEDCT_US|Secretory carcinoma of the breast|8508/3
C3839648|T191|PT|703546002|SNOMEDCT_US|Solid papillary carcinoma in situ|8509/2
C3839652|T191|PT|703594003|SNOMEDCT_US|Solid papillary carcinoma with invasion|8509/3
C0206693|T191|PT|0000021025|CHV|medullary carcinoma|8510/3
C0206693|T191|LA|LA26495-4|LNC|Medullary carcinoma, NOS|8510/3
C0206693|T191|PT|271442|MEDCIN|medullary carcinoma|8510/3
C0206693|T191|MH|D018276|MSH|Carcinoma, Medullary|8510/3
C0206693|T191|PM|D018276|MSH|Carcinomas, Medullary|8510/3
C0206693|T191|PM|D018276|MSH|Medullary Carcinoma|8510/3
C0206693|T191|PM|D018276|MSH|Medullary Carcinomas|8510/3
C0206693|T191|PN|NOCODE|MTH|Medullary carcinoma|8510/3
C0206693|T191|OP|C66718|NCI|Medullary Carcinoma, NOS|8510/3
C0206693|T191|OP|C66718|NCI|Medullary Carcinoma, Not Otherwise Specified|8510/3
C0206693|T191|PT|C66718|NCI|Medullary Carcinoma, Not Otherwise Specified|8510/3
C0206693|T191|SY|Xa98x|RCD|Medullary adenocarcinoma|8510/3
C0206693|T191|PT|Xa98x|RCD|Medullary carcinoma|8510/3
C0206693|T191|OP|BB9B.|RCDSY|Medullary carcinoma NOS|8510/3
C0206693|T191|SY|32913002|SNOMEDCT_US|Medullary adenocarcinoma|8510/3
C0206693|T191|PT|32913002|SNOMEDCT_US|Medullary carcinoma|8510/3
C0206693|T191|IS|32913002|SNOMEDCT_US|Medullary carcinoma, NOS|8510/3
C3839099|T191|PT|703595002|SNOMEDCT_US|Medullary-like carcinoma|8510/3
C0860580|T191|SY|0000050759|CHV|breast carcinoma medullary|8512/3
C0860580|T191|SY|0000050759|CHV|medullary breast carcinoma|8512/3
C0860580|T191|SY|0000050759|CHV|medullary carcinoma breast|8512/3
C0860580|T191|PT|0000050759|CHV|medullary carcinoma of breast|8512/3
C0334380|T191|PT|MTHU014794|ICPC2ICD10ENG|carcinoma; medullary with lymphoid stroma, unspecified site|8512/3
C0334380|T191|PT|MTHU048009|ICPC2ICD10ENG|medullary; carcinoma with lymphoid stroma, unspecified site|8512/3
C0860580|T191|LLT|10027095|MDR|Medullary carcinoma of breast|8512/3
C0860580|T191|PT|10027095|MDR|Medullary carcinoma of breast|8512/3
C0860580|T191|PT|232315|MEDCIN|medullary carcinoma of breast|8512/3
C0860580|T191|PN|NOCODE|MTH|Medullary carcinoma of breast|8512/3
C0860580|T191|SY|C9119|NCI|Infiltrating Medullary Carcinoma of Breast|8512/3
C0860580|T191|SY|C9119|NCI|Infiltrating Medullary Carcinoma of the Breast|8512/3
C0860580|T191|SY|C9119|NCI|Invasive Medullary Breast Carcinoma|8512/3
C0860580|T191|SY|C9119|NCI|Invasive Medullary Carcinoma of Breast|8512/3
C0860580|T191|SY|C9119|NCI|Invasive Medullary Carcinoma of the Breast|8512/3
C0860580|T191|PT|C9119|NCI|Medullary Breast Carcinoma|8512/3
C0860580|T191|SY|C9119|NCI|Medullary Breast Carcinoma with Lymphoid Stroma|8512/3
C0860580|T191|SY|C9119|NCI|Medullary Carcinoma of Breast|8512/3
C0860580|T191|SY|C9119|NCI|Medullary Carcinoma of the Breast|8512/3
C0860580|T191|DN|C9119|NCI_CTRP|Medullary Breast Cancer|8512/3
C0860580|T191|PT|CDR0000044532|NCI_NCI-GLOSS|medullary breast carcinoma|8512/3
C0334380|T191|AB|BB9D.|RCD|Medullary ca + lymphoid stroma|8512/3
C0334380|T191|PT|BB9D.|RCD|Medullary carcinoma with lymphoid stroma|8512/3
C0334380|T191|PT|85654004|SNOMEDCT_US|Medullary carcinoma with lymphoid stroma|8512/3
C1879758|T191|PT|232317|MEDCIN|atypical medullary carcinoma of breast|8513/3
C1879758|T191|PT|C66719|NCI|Atypical Medullary Breast Carcinoma|8513/3
C1879758|T191|SY|C66719|NCI|Infiltrating Ductal Breast Carcinoma with Medullary Features|8513/3
C1266082|T191|PT|128698005|SNOMEDCT_US|Atypical medullary carcinoma|8513/3
C0346151|T191|SY|31657|MEDCIN|breast malignant carcinoma scirrhous|8514/3
C0346151|T191|PT|31657|MEDCIN|scirrhous carcinoma of breast|8514/3
C0346151|T191|SY|C7362|NCI|Infiltrating Carcinoma of Breast with Fibrotic Stroma|8514/3
C0346151|T191|SY|C7362|NCI|Infiltrating Carcinoma of the Breast with Fibrotic Stroma|8514/3
C0346151|T191|PT|C7362|NCI|Scirrhous Breast Carcinoma|8514/3
C0346151|T191|SY|C7362|NCI|Scirrhous Carcinoma of Breast|8514/3
C0346151|T191|SY|C7362|NCI|Scirrhous Carcinoma of the Breast|8514/3
C0346151|T191|PT|X78WO|RCD|Scirrhous carcinoma of breast|8514/3
C1266083|T191|PT|128699002|SNOMEDCT_US|Duct carcinoma, desmoplastic type|8514/3
C0346151|T191|PT|254839007|SNOMEDCT_US|Scirrhous carcinoma of breast|8514/3
C2919327|T191|SY|444591006|SNOMEDCT_US|LCIS, pleomorphic|8519/2
C2919327|T191|PT|444591006|SNOMEDCT_US|Pleomorphic lobular carcinoma in situ|8519/2
C0279563|T191|SY|0000027266|CHV|breast cancer lobular in situ|8520/2
C0279563|T191|SY|0000027266|CHV|breast carcinoma lobular situ|8520/2
C0279563|T191|SY|0000027266|CHV|breast lobular cancer in situ|8520/2
C0334381|T191|SY|0000029968|CHV|lcis|8520/2
C0279563|T191|SY|0000027266|CHV|lobular breast cancer in situ|8520/2
C0279563|T191|SY|0000027266|CHV|lobular breast carcinoma in situ|8520/2
C0279563|T191|PT|0000027266|CHV|lobular carcinoma in situ|8520/2
C0334381|T191|PT|0000029968|CHV|lobular carcinoma in situ|8520/2
C0334381|T191|SY|0000029968|CHV|lobular carcinoma in-situ|8520/2
C0279563|T191|PT|HP:0030076|HPO|Lobular carcinoma in situ|8520/2
C0334381|T191|PT|D05.0|ICD10|Lobular carcinoma in situ|8520/2
C0279563|T191|AB|D05.0|ICD10CM|Lobular carcinoma in situ of breast|8520/2
C0279563|T191|HT|D05.0|ICD10CM|Lobular carcinoma in situ of breast|8520/2
C0279563|T191|PT|MTHU047382|ICPC2ICD10ENG|breast; carcinoma in situ, lobular|8520/2
C0279563|T191|PT|MTHU047387|ICPC2ICD10ENG|breast; carcinoma, lobular, noninfiltrating|8520/2
C0279563|T191|PT|MTHU047437|ICPC2ICD10ENG|breast; lobular, noninfiltrating carcinoma|8520/2
C0279563|T191|PT|MTHU047453|ICPC2ICD10ENG|breast; noninfiltrating lobular carcinoma|8520/2
C0279563|T191|PT|MTHU014716|ICPC2ICD10ENG|carcinoma in situ; lobular, breast|8520/2
C0279563|T191|PT|MTHU014791|ICPC2ICD10ENG|carcinoma; lobular, noninfiltrating, breast|8520/2
C0279563|T191|PT|MTHU045799|ICPC2ICD10ENG|lobular; carcinoma in situ, breast|8520/2
C0279563|T191|PT|MTHU045807|ICPC2ICD10ENG|lobular; carcinoma, noninfiltrating, breast|8520/2
C0334381|T191|CN|MTHU056197|LNC|Lobular carcinoma in situ|8520/2
C0334381|T191|LPN|LP247941-0|LNC|Lobular carcinoma in situ|8520/2
C0279563|T191|LLT|10073099|MDR|Lobular breast carcinoma in situ|8520/2
C0279563|T191|PT|10073099|MDR|Lobular breast carcinoma in situ|8520/2
C0279563|T191|PT|232268|MEDCIN|lobular carcinoma in situ of breast|8520/2
C0334381|T191|ET|D000071960|MSH|LCIS, Lobular Carcinoma In Situ|8520/2
C0334381|T191|PEP|D000071960|MSH|Lobular Carcinoma In Situ|8520/2
C0279563|T191|PN|NOCODE|MTH|Lobular carcinoma in situ of breast|8520/2
C0334381|T191|PN|NOCODE|MTH|Non-infiltrating lobular carcinoma|8520/2
C0279563|T191|SY|C4018|NCI|LCIS|8520/2
C0279563|T191|PT|C4018|NCI|Lobular Breast Carcinoma In Situ|8520/2
C0279563|T191|SY|TCGA|NCI|Lobular Breast Carcinoma In Situ|8520/2
C0279563|T191|SY|C4018|NCI|Lobular Ca in situ of Breast|8520/2
C0279563|T191|SY|C4018|NCI|Lobular Ca in situ of the Breast|8520/2
C0279563|T191|SY|C4018|NCI|Lobular Carcinoma in situ|8520/2
C0279563|T191|SY|C4018|NCI|Lobular Carcinoma in situ of Breast|8520/2
C0279563|T191|SY|C4018|NCI|Lobular Carcinoma In Situ of the Breast|8520/2
C0279563|T191|SY|C4018|NCI|Non-Infiltrating Lobular Breast Carcinoma|8520/2
C0279563|T191|SY|C4018|NCI|Non-Infiltrating Lobular Carcinoma|8520/2
C0279563|T191|SY|C4018|NCI|Non-Infiltrating Lobular Carcinoma of Breast|8520/2
C0279563|T191|SY|C4018|NCI|Non-Infiltrating Lobular Carcinoma of the Breast|8520/2
C0279563|T191|SY|C4018|NCI|Non-Invasive Lobular Breast Carcinoma|8520/2
C0279563|T191|SY|C4018|NCI|Non-Invasive Lobular Carcinoma of Breast|8520/2
C0279563|T191|SY|C4018|NCI|Non-Invasive Lobular Carcinoma of the Breast|8520/2
C0279563|T191|PT|10024744|NCI_CTEP-SDC|Lobular carcinoma in situ|8520/2
C0279563|T191|PT|CDR0000044433|NCI_NCI-GLOSS|LCIS|8520/2
C0279563|T191|PT|CDR0000046315|NCI_NCI-GLOSS|lobular carcinoma in situ|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|in situ lobular breast carcinoma|8520/2
C0334381|T191|SY|CDR0000039848|PDQ|LCIS|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|LCIS of the breast|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|lobular breast cancer in situ|8520/2
C0279563|T191|PT|CDR0000039848|PDQ|lobular breast carcinoma in situ|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|lobular breast carcinoma, in situ|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Lobular Ca in situ of Breast|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Lobular Ca in situ of the Breast|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|lobular cancer in situ of the breast|8520/2
C0334381|T191|SY|CDR0000039848|PDQ|lobular carcinoma in situ|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Lobular Carcinoma in situ of Breast|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Lobular Carcinoma In Situ of the Breast|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|lobular in situ breast carcinoma|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Non-Infiltrating Lobular Breast Carcinoma|8520/2
C0334381|T191|SY|CDR0000039848|PDQ|Non-Infiltrating Lobular Carcinoma|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Non-Infiltrating Lobular Carcinoma of Breast|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Non-Infiltrating Lobular Carcinoma of the Breast|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Non-Invasive Lobular Breast Carcinoma|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Non-Invasive Lobular Carcinoma of Breast|8520/2
C0279563|T191|SY|CDR0000039848|PDQ|Non-Invasive Lobular Carcinoma of the Breast|8520/2
C0334381|T191|AB|BB9E.|RCD|LCIS - Lobular carc in situ|8520/2
C0334381|T191|SY|BB9E.|RCD|LCIS - Lobular carcinoma in situ|8520/2
C0279563|T191|AB|X78WV|RCD|Lobular ca in situ of breast|8520/2
C0334381|T191|PT|BB9E.|RCD|Lobular carcinoma in situ|8520/2
C0279563|T191|PT|X78WV|RCD|Lobular carcinoma in situ of breast|8520/2
C0334381|T191|AB|BB9E.|RCD|Non-infiltrating lobular ca|8520/2
C0334381|T191|SY|BB9E.|RCD|Non-infiltrating lobular carcinoma|8520/2
C2919427|T191|PT|444739008|SNOMEDCT_US|Classic lobular carcinoma in situ|8520/2
C0334381|T191|SY|77284006|SNOMEDCT_US|LCIS|8520/2
C0334381|T191|SY|77284006|SNOMEDCT_US|LCIS - Lobular carcinoma in situ|8520/2
C0334381|T191|PT|77284006|SNOMEDCT_US|Lobular carcinoma in situ|8520/2
C0279563|T191|PT|109888004|SNOMEDCT_US|Lobular carcinoma in situ of breast|8520/2
C0279563|T191|OAP|189337009|SNOMEDCT_US|Lobular carcinoma in situ of breast|8520/2
C0279563|T191|OF|189337009|SNOMEDCT_US|Lobular carcinoma in situ of breast|8520/2
C0334381|T191|SY|77284006|SNOMEDCT_US|Lobular carcinoma, noninfiltrating|8520/2
C0334381|T191|SY|77284006|SNOMEDCT_US|Non-infiltrating lobular carcinoma|8520/2
C0206692|T191|SY|0000021024|CHV|breast carcinoma lobular|8520/3
C0206692|T191|SY|0000021024|CHV|carcinoma infiltrated lobular|8520/3
C0206692|T191|SY|0000021024|CHV|carcinoma lobular|8520/3
C0206692|T191|SY|0000021024|CHV|infiltrating lobular carcinoma|8520/3
C0206692|T191|SY|0000021024|CHV|lobular breast carcinoma|8520/3
C0206692|T191|PT|0000021024|CHV|lobular carcinoma|8520/3
C0206692|T191|SY|0000021024|CHV|lobular carcinoma breast|8520/3
C0206692|T191|SY|0000021024|CHV|lobular carcinoma of breast|8520/3
C0206692|T191|SY|0000021024|CHV|lobular carcinomas|8520/3
C0206692|T191|LLT|10024750|MDR|Lobular carcinoma of breast|8520/3
C0206692|T191|PT|232319|MEDCIN|lobular carcinoma of breast|8520/3
C0206692|T191|MH|D018275|MSH|Carcinoma, Lobular|8520/3
C0206692|T191|PM|D018275|MSH|Carcinomas, Lobular|8520/3
C0206692|T191|PM|D018275|MSH|Lobular Carcinoma|8520/3
C0206692|T191|PM|D018275|MSH|Lobular Carcinomas|8520/3
C0206692|T191|PN|NOCODE|MTH|Carcinoma, Lobular|8520/3
C0206692|T191|SY|C3771|NCI|Lobular Adenocarcinoma|8520/3
C0206692|T191|PT|C3771|NCI|Lobular Breast Carcinoma|8520/3
C0206692|T191|SY|C3771|NCI|Lobular Carcinoma|8520/3
C0206692|T191|SY|C3771|NCI|Lobular Carcinoma of Breast|8520/3
C0206692|T191|SY|C3771|NCI|Lobular Carcinoma of the Breast|8520/3
C0206692|T191|DN|C3771|NCI_CTRP|Lobular Breast Carcinoma|8520/3
C0206692|T191|PT|CDR0000426416|NCI_NCI-GLOSS|lobular carcinoma|8520/3
C0206692|T191|SY|CDR0000039847|PDQ|lobular adenocarcinoma|8520/3
C0206692|T191|PT|CDR0000039847|PDQ|lobular breast carcinoma|8520/3
C0206692|T191|SY|CDR0000039847|PDQ|lobular carcinoma|8520/3
C0206692|T191|SY|CDR0000039847|PDQ|lobular carcinoma of breast|8520/3
C0206692|T191|SY|CDR0000039847|PDQ|lobular carcinoma of the breast|8520/3
C0206692|T191|SY|Xa98y|RCD|Infiltrating lobular carcinoma|8520/3
C0206692|T191|SY|Xa98y|RCD|Lobular adenocarcinoma|8520/3
C0206692|T191|PT|Xa98y|RCD|Lobular carcinoma|8520/3
C0206692|T191|PT|Xa0bU|RCD|Lobular carcinoma of breast|8520/3
C0206692|T191|OP|BB9F.|RCDSY|Lobular carcinoma NOS|8520/3
C0206692|T191|SY|89740008|SNOMEDCT_US|Infiltrating lobular carcinoma|8520/3
C0206692|T191|PT|278054005|SNOMEDCT_US|Infiltrating lobular carcinoma of breast|8520/3
C0206692|T191|SY|89740008|SNOMEDCT_US|Lobular adenocarcinoma|8520/3
C0206692|T191|PT|89740008|SNOMEDCT_US|Lobular carcinoma|8520/3
C0206692|T191|SY|278054005|SNOMEDCT_US|Lobular carcinoma of breast|8520/3
C0206692|T191|IS|89740008|SNOMEDCT_US|Lobular carcinoma, NOS|8520/3
C3838879|T191|PT|703596001|SNOMEDCT_US|Tubulolobular carcinoma|8520/3
C1134719|T191|PT|0042764|CCPSS|BREAST CANCER DUCTAL INFILTRATING|8521/3
C1134719|T191|SY|0000050852|CHV|breast cancer invasive ductal|8521/3
C1134719|T191|SY|0000056504|CHV|breast carcinoma ductal invasive|8521/3
C1134719|T191|SY|0000050852|CHV|cancer breast invasive ductal|8521/3
C1134719|T191|SY|0000054856|CHV|carcinoma ductal infiltrate|8521/3
C1134719|T191|SY|0000054856|CHV|carcinoma ductal infiltrated|8521/3
C1134719|T191|SY|0000056504|CHV|carcinoma infiltrating duct|8521/3
C1134719|T191|SY|0000054856|CHV|carcinomas ductal infiltrating|8521/3
C1134719|T191|SY|0000054856|CHV|ductal infiltrating carcinoma|8521/3
C1134719|T191|SY|0000050852|CHV|ductal invasive breast cancer|8521/3
C1134719|T191|PT|0000054856|CHV|infiltrating ductal carcinoma|8521/3
C1134719|T191|PT|0000050852|CHV|invasive ductal breast cancer|8521/3
C1134719|T191|PT|0000056504|CHV|invasive ductal breast carcinoma|8521/3
C1134719|T191|SY|0000056504|CHV|invasive ductal carcinoma breast|8521/3
C1134719|T191|PT|MTHU014743|ICPC2ICD10ENG|carcinoma; ductal, infiltrating, unspecified site|8521/3
C1134719|T191|PT|MTHU014744|ICPC2ICD10ENG|carcinoma; ductular, infiltrating, unspecified site|8521/3
C1134719|T191|PT|MTHU014770|ICPC2ICD10ENG|carcinoma; infiltrating duct, unspecified site|8521/3
C1134719|T191|PT|MTHU014771|ICPC2ICD10ENG|carcinoma; infiltrating ductular, unspecified site|8521/3
C1134719|T191|PT|MTHU024095|ICPC2ICD10ENG|ductal; carcinoma, infiltrating, unspecified site|8521/3
C1134719|T191|PT|MTHU024097|ICPC2ICD10ENG|ductular; carcinoma, infiltrating, unspecified site|8521/3
C1134719|T191|PT|MTHU039173|ICPC2ICD10ENG|infiltrating; ductal adenocarcinoma, unspecified site|8521/3
C1134719|T191|PT|MTHU039175|ICPC2ICD10ENG|infiltrating; ductal carcinoma, unspecified site|8521/3
C1134719|T191|PT|MTHU039176|ICPC2ICD10ENG|infiltrating; ductular carcinoma, unspecified site|8521/3
C1134719|T191|LLT|10006235|MDR|Breast ductal cancer infiltrating|8521/3
C1134719|T191|LLT|10006236|MDR|Breast ductal cancer invasive|8521/3
C1134719|T191|LLT|10021944|MDR|Infiltrating ductal breast cancer|8521/3
C1134719|T191|LLT|10022882|MDR|Invasive ductal breast cancer|8521/3
C1134719|T191|LLT|10073095|MDR|Invasive ductal breast carcinoma|8521/3
C1134719|T191|PT|10073095|MDR|Invasive ductal breast carcinoma|8521/3
C1134719|T191|PT|232310|MEDCIN|infiltrating ductal carcinoma of breast|8521/3
C1134719|T191|MH|D018270|MSH|Carcinoma, Ductal, Breast|8521/3
C1134719|T191|ET|D018270|MSH|Carcinoma, Infiltrating Duct|8521/3
C1134719|T191|ET|D018270|MSH|Carcinoma, Invasive Ductal, Breast|8521/3
C1134719|T191|PM|D018270|MSH|Carcinomas, Infiltrating Duct|8521/3
C1134719|T191|ET|D018270|MSH|Invasive Ductal Carcinoma, Breast|8521/3
C1134719|T191|PN|NOCODE|MTH|Invasive Ductal Breast Carcinoma|8521/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Adenocarcinoma|8521/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Breast Carcinoma|8521/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Carcinoma|8521/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Carcinoma of Breast|8521/3
C1134719|T191|SY|C4194|NCI|Infiltrating Ductal Carcinoma of the Breast|8521/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Adenocarcinoma|8521/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Breast Carcinoma|8521/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma|8521/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma of Breast|8521/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma of the Breast|8521/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma, No Specific Type|8521/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma, NOS|8521/3
C1134719|T191|SY|TCGA|NCI|Invasive Ductal Carcinoma, Not Otherwise Specified|8521/3
C1134719|T191|PT|C4194|NCI|Invasive Ductal Carcinoma, Not Otherwise Specified|8521/3
C1134719|T191|SY|C4194|NCI|Invasive Ductal Carcinoma, NST|8521/3
C1134719|T191|DN|C4194|NCI_CTRP|Invasive Ductal Carcinoma, NOS|8521/3
C1134719|T191|PT|CDR0000045099|NCI_NCI-GLOSS|infiltrating ductal carcinoma|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|ductal invasive breast carcinoma|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Adenocarcinoma|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Breast Carcinoma|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Carcinoma|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Carcinoma of Breast|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Infiltrating Ductal Carcinoma of the Breast|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Adenocarcinoma|8521/3
C1134719|T191|PT|CDR0000039843|PDQ|invasive ductal breast carcinoma|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma of Breast|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma of the Breast|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma, No Specific Type|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma, NOS|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma, Not Otherwise Specified|8521/3
C1134719|T191|SY|CDR0000039843|PDQ|Invasive Ductal Carcinoma, NST|8521/3
C1134719|T191|AB|BB9G.|RCD|Infiltrating ductular ca|8521/3
C1134719|T191|PT|BB9G.|RCD|Infiltrating ductular carcinoma|8521/3
C1134719|T191|PT|408643008|SNOMEDCT_US|Infiltrating duct carcinoma of breast|8521/3
C1134719|T191|SY|408643008|SNOMEDCT_US|Infiltrating ductal carcinoma of breast|8521/3
C1134719|T191|PT|58477004|SNOMEDCT_US|Infiltrating ductular carcinoma|8521/3
C1134719|T191|SY|408643008|SNOMEDCT_US|Invasive duct carcinoma of breast|8521/3
C1134719|T191|SY|408643008|SNOMEDCT_US|Invasive ductal carcinoma of breast|8521/3
C0334383|T191|PT|MTHU047384|ICPC2ICD10ENG|breast; carcinoma in situ, lobular with intraductal|8522/2
C0334383|T191|PT|MTHU014714|ICPC2ICD10ENG|carcinoma in situ; lobular with intraductal, breast|8522/2
C0334383|T191|PT|MTHU045802|ICPC2ICD10ENG|lobular; carcinoma in situ, with intraductal, breast|8522/2
C0334383|T191|PT|232269|MEDCIN|intraductal and lobular carcinoma in situ of breast|8522/2
C0334383|T191|SY|C4195|NCI|DCIS and LCIS of Breast|8522/2
C0334383|T191|SY|C4195|NCI|DCIS and LCIS of the Breast|8522/2
C0334383|T191|SY|C4195|NCI|Ductal and Lobular Breast Carcinoma in situ|8522/2
C0334383|T191|SY|C4195|NCI|Ductal and Lobular Carcinoma in situ of Breast|8522/2
C0334383|T191|SY|C4195|NCI|Ductal and Lobular Carcinoma in situ of the Breast|8522/2
C0334383|T191|PT|C4195|NCI|Ductal Breast Carcinoma In Situ and Lobular Carcinoma In Situ|8522/2
C0334383|T191|SY|TCGA|NCI|Ductal Breast Carcinoma In Situ and Lobular Carcinoma In Situ|8522/2
C0334383|T191|SY|C4195|NCI|Ductal Carcinoma in situ with Lobular Carcinoma in situ of Breast|8522/2
C0334383|T191|SY|C4195|NCI|Ductal Carcinoma in situ with Lobular Carcinoma in situ of the Breast|8522/2
C0334383|T191|SY|C4195|NCI|Intraductal and Lobular Breast Carcinoma in situ|8522/2
C0334383|T191|SY|C4195|NCI|Intraductal and Lobular Carcinoma in situ of Breast|8522/2
C0334383|T191|SY|C4195|NCI|Intraductal and Lobular Carcinoma in situ of the Breast|8522/2
C0334383|T191|SY|C4195|NCI|Intraductal Carcinoma and Lobular Carcinoma in situ|8522/2
C0334383|T191|SY|C4195|NCI|Non-Infiltrating Ductal and Non-Infiltrating Lobular Breast Carcinoma|8522/2
C0334383|T191|SY|C4195|NCI|Non-Infiltrating Ductal with Non-Infiltrating Lobular Carcinoma of Breast|8522/2
C0334383|T191|SY|C4195|NCI|Non-Infiltrating Ductal with Non-Infiltrating Lobular Carcinoma of the Breast|8522/2
C0334383|T191|SY|C4195|NCI|Non-Invasive Ductal and Non-Invasive Lobular Breast Carcinoma|8522/2
C0334383|T191|SY|C4195|NCI|Non-Invasive Ductal and Non-Invasive Lobular Carcinoma|8522/2
C0334383|T191|SY|C4195|NCI|Non-Invasive Ductal Breast Carcinoma with Non-Invasive Lobular Breast Carcinoma|8522/2
C0334383|T191|SY|C4195|NCI|Non-Invasive Ductal Carcinoma with Non-Invasive Lobular Carcinoma of Breast|8522/2
C0334383|T191|SY|C4195|NCI|Non-Invasive Ductal Carcinoma with Non-Invasive Lobular Carcinoma of the Breast|8522/2
C0334383|T191|SY|C4195|NCI|Non-Invasive Ductal with Non-Invasive Lobular Breast Carcinoma|8522/2
C0334383|T191|AB|X77o0|RCD|Intraduct ca+lobul ca in situ|8522/2
C0334383|T191|PT|X77o0|RCD|Intraductal carcinoma and lobular carcinoma in situ|8522/2
C0334383|T191|OA|BB9E0|RCDSY|Intrad carc+lobul carc situ|8522/2
C0334383|T191|OP|BB9E0|RCDSY|Intraductal carcinoma and lobular carcinoma in situ|8522/2
C0334383|T191|PT|18680006|SNOMEDCT_US|Intraductal carcinoma and lobular carcinoma in situ|8522/2
C0334384|T191|PT|MTHU014769|ICPC2ICD10ENG|carcinoma; infiltrating duct with lobular ca, unspecified site|8522/3
C0334384|T191|LLT|10073983|MDR|Mixed ductal lobular breast carcinoma|8522/3
C0334384|T191|SY|355752|MEDCIN|breast neoplasm malignant carcinoma with ductal and lobular features|8522/3
C0334384|T191|PT|355752|MEDCIN|Carcinoma of breast with ductal and lobular features|8522/3
C0334384|T191|SY|C6939|NCI|DCIS and ILC|8522/3
C0334384|T191|SY|C6939|NCI|DCIS and Infiltrating Lobular Carcinoma|8522/3
C0334384|T191|SY|C5160|NCI|Ductal and Lobular Carcinoma|8522/3
C0334384|T191|PT|C6939|NCI|Ductal Breast Carcinoma In Situ and Invasive Lobular Carcinoma|8522/3
C0334384|T191|SY|C6939|NCI|Ductal Carcinoma in situ and Infiltrating Lobular Carcinoma|8522/3
C1334277|T191|SY|C7688|NCI|Infiltrating Ductal and Lobular Carcinoma|8522/3
C0334384|T191|SY|C7689|NCI|Infiltrating Ductal and Lobular Carcinoma in situ|8522/3
C0334384|T191|PT|C7690|NCI|Intraductal and Lobular Carcinoma|8522/3
C1334277|T191|SY|C7688|NCI|Invasive Duct and Lobular Carcinoma|8522/3
C1334277|T191|PT|C7688|NCI|Invasive Ductal and Lobular Carcinoma|8522/3
C0334384|T191|PT|C7689|NCI|Invasive Ductal and Lobular Carcinoma In Situ|8522/3
C0334384|T191|SY|C7689|NCI|LCIS and Infiltrating Ductal Carcinoma|8522/3
C0334384|T191|SY|C7689|NCI|Lobular Carcinoma in situ and Infiltrating Ductal Carcinoma|8522/3
C0334384|T191|SY|C7689|NCI|Lobular Carcinoma in situ and Invasive Ductal Carcinoma|8522/3
C0334384|T191|SY|C5160|NCI|Mixed Ductal and Lobular Breast Carcinoma|8522/3
C0334384|T191|SY|C5160|NCI|Mixed Ductal and Lobular Carcinoma of Breast|8522/3
C0334384|T191|SY|C5160|NCI|Mixed Ductal and Lobular Carcinoma of the Breast|8522/3
C0334384|T191|PT|C5160|NCI|Mixed Lobular and Ductal Breast Carcinoma|8522/3
C0334384|T191|SY|C5160|NCI|Mixed Lobular and Ductal Carcinoma|8522/3
C0334384|T191|SY|C5160|NCI|Mixed Lobular and Ductal Carcinoma of Breast|8522/3
C0334384|T191|SY|C5160|NCI|Mixed Lobular and Ductal Carcinoma of the Breast|8522/3
C0334384|T191|SY|C6939|NCI|Non-Infiltrating Ductal Carcinoma and ILC|8522/3
C0334384|T191|SY|C6939|NCI|Non-Infiltrating Ductal Carcinoma and Infiltrating Lobular Carcinoma|8522/3
C0334384|T191|AB|X77nw|RCD|Infilt duct+lobular ca in situ|8522/3
C0334384|T191|AB|X77nw|RCD|Infiltrating duct + lobular ca|8522/3
C0334384|T191|PT|X77nw|RCD|Infiltrating duct and lobular carcinoma|8522/3
C0334384|T191|SY|X77nw|RCD|Infiltrating duct and lobular carcinoma in situ|8522/3
C0334384|T191|AB|X77nw|RCD|Intraductal and lobular ca|8522/3
C0334384|T191|SY|X77nw|RCD|Intraductal and lobular carcinoma|8522/3
C0334384|T191|SY|X77nw|RCD|Lobular and ductal carcinoma|8522/3
C0334384|T191|AB|X77nw|RCDSY|Infiltr duct+lobul carcinom|8522/3
C0334384|T191|SY|444604002|SNOMEDCT_US|Carcinoma of breast with ductal and lobular features|8522/3
C2732747|T191|PT|444057000|SNOMEDCT_US|Infiltrating carcinoma with ductal and lobular features|8522/3
C0334384|T191|PT|35232005|SNOMEDCT_US|Infiltrating duct and lobular carcinoma|8522/3
C0334384|T191|OAP|189707003|SNOMEDCT_US|Infiltrating duct and lobular carcinoma|8522/3
C0334384|T191|OF|189707003|SNOMEDCT_US|Infiltrating duct and lobular carcinoma|8522/3
C0334384|T191|SY|35232005|SNOMEDCT_US|Infiltrating duct and lobular carcinoma in situ|8522/3
C0334384|T191|SY|35232005|SNOMEDCT_US|Infiltrating lobular carcinoma and ductal carcinoma in situ|8522/3
C0334384|T191|SY|35232005|SNOMEDCT_US|Intraductal and lobular carcinoma|8522/3
C0334384|T191|SY|35232005|SNOMEDCT_US|Lobular and ductal carcinoma|8522/3
C0334384|T191|PT|444604002|SNOMEDCT_US|Mixed ductal and lobular carcinoma of breast|8522/3
C1517577|T191|SY|C40347|NCI|Infiltrating Mixed Breast Carcinoma|8523/3
C1517577|T191|PT|C40347|NCI|Invasive Mixed Breast Carcinoma|8523/3
C1266084|T191|SY|128700001|SNOMEDCT_US|Infiltrating duct and colloid carcinoma|8523/3
C1266084|T191|SY|128700001|SNOMEDCT_US|Infiltrating duct and cribriform carcinoma|8523/3
C1266084|T191|SY|128700001|SNOMEDCT_US|Infiltrating duct and mucinous carcinoma|8523/3
C1266084|T191|SY|128700001|SNOMEDCT_US|Infiltrating duct and tubular carcinoma|8523/3
C1266084|T191|PT|128700001|SNOMEDCT_US|Infiltrating duct mixed with other types of carcinoma|8523/3
C1517577|T191|SY|C40347|NCI|Infiltrating Mixed Breast Carcinoma|8524/3
C1517577|T191|PT|C40347|NCI|Invasive Mixed Breast Carcinoma|8524/3
C1266085|T191|PT|128701002|SNOMEDCT_US|Infiltrating lobular mixed with other types of carcinoma|8524/3
C1335907|T191|PT|39574|MEDCIN|polymorphous low grade adenocarcinoma of salivary gland|8525/3
C1335907|T191|PT|355370|MEDCIN|polymorphous low-grade adenocarcinoma of salivary gland|8525/3
C1335907|T191|PT|82865|MEDCIN|Salivary gland biopsy: polymorphous low-grade adenocarcinoma of salivary gland|8525/3
C1335907|T191|SY|355370|MEDCIN|salivary gland carcinoma polymorphous low-grade adenocarcinoma|8525/3
C1266086|T191|PN|NOCODE|MTH|Polymorphous low grade adenocarcinoma|8525/3
C1335907|T191|PN|NOCODE|MTH|Polymorphous low grade adenocarcinoma of salivary gland|8525/3
C1335907|T191|SY|C35702|NCI|Polymorphous adenocarcinoma, classic|8525/3
C1335907|T191|SY|C35702|NCI|Salivary Gland Polymorphous Adenocarcinoma, Classical Variant|8525/3
C1335907|T191|PT|C35702|NCI|Salivary Gland Polymorphous Low Grade Adenocarcinoma|8525/3
C1335907|T191|SY|C35702|NCI|Salivary Gland Terminal Duct Adenocarcinoma|8525/3
C1266086|T191|PT|128702009|SNOMEDCT_US|Polymorphous low grade adenocarcinoma|8525/3
C1335907|T191|PT|423038006|SNOMEDCT_US|Polymorphous low grade adenocarcinoma of salivary gland|8525/3
C1266086|T191|SY|128702009|SNOMEDCT_US|Terminal duct adenocarcinoma|8525/3
C0278601|T191|SY|0000027199|CHV|breast cancer inflammatory|8530/3
C0278601|T191|SY|0000027199|CHV|breast inflammatory cancer|8530/3
C0278601|T191|SY|0000027199|CHV|breast inflammatory carcinoma|8530/3
C0278601|T191|PT|0000027199|CHV|inflammatory breast cancer|8530/3
C0278601|T191|SY|0000027199|CHV|inflammatory breast carcinoma|8530/3
C0278601|T191|SY|0000027199|CHV|inflammatory cancer breast|8530/3
C0334385|T191|PT|0000029969|CHV|inflammatory carcinoma|8530/3
C0278601|T191|SY|0000027199|CHV|inflammatory carcinoma breast|8530/3
C0334385|T191|PT|MTHU014773|ICPC2ICD10ENG|carcinoma; inflammatory, unspecified site|8530/3
C0334385|T191|PT|MTHU039180|ICPC2ICD10ENG|inflammatory; carcinoma, unspecified site|8530/3
C0278601|T191|LLT|10006205|MDR|Breast carcinoma inflammatory|8530/3
C0278601|T191|LLT|10021974|MDR|Inflammatory breast cancer|8530/3
C0278601|T191|LLT|10021980|MDR|Inflammatory carcinoma of the breast|8530/3
C0278601|T191|PT|10021980|MDR|Inflammatory carcinoma of the breast|8530/3
C0278601|T191|PT|232324|MEDCIN|inflammatory carcinoma of breast|8530/3
C0278601|T191|PM|D058922|MSH|Breast Cancer, Inflammatory|8530/3
C0278601|T191|PM|D058922|MSH|Breast Cancers, Inflammatory|8530/3
C0278601|T191|PM|D058922|MSH|Breast Carcinoma, Inflammatory|8530/3
C0278601|T191|PM|D058922|MSH|Breast Carcinomas, Inflammatory|8530/3
C0278601|T191|PM|D058922|MSH|Breast Neoplasm, Inflammatory|8530/3
C0278601|T191|PM|D058922|MSH|Breast Neoplasms, Inflammatory|8530/3
C0278601|T191|PM|D058922|MSH|Cancer, Inflammatory Breast|8530/3
C0278601|T191|PM|D058922|MSH|Cancers, Inflammatory Breast|8530/3
C0278601|T191|PM|D058922|MSH|Carcinoma, Inflammatory Breast|8530/3
C0278601|T191|PM|D058922|MSH|Carcinomas, Inflammatory Breast|8530/3
C0278601|T191|ET|D058922|MSH|Inflammatory Breast Cancer|8530/3
C0278601|T191|PM|D058922|MSH|Inflammatory Breast Cancers|8530/3
C0278601|T191|ET|D058922|MSH|Inflammatory Breast Carcinoma|8530/3
C0278601|T191|PM|D058922|MSH|Inflammatory Breast Carcinomas|8530/3
C0278601|T191|PM|D058922|MSH|Inflammatory Breast Neoplasm|8530/3
C0278601|T191|MH|D058922|MSH|Inflammatory Breast Neoplasms|8530/3
C0278601|T191|PM|D058922|MSH|Neoplasm, Inflammatory Breast|8530/3
C0278601|T191|PM|D058922|MSH|Neoplasms, Inflammatory Breast|8530/3
C0278601|T191|PN|NOCODE|MTH|Inflammatory Breast Carcinoma|8530/3
C0334385|T191|PN|NOCODE|MTH|Inflammatory carcinoma|8530/3
C0278601|T191|SY|C4001|NCI|Inflammatory Breast Cancer|8530/3
C0278601|T191|PT|C4001|NCI|Inflammatory Breast Carcinoma|8530/3
C0278601|T191|SY|C4001|NCI|Inflammatory Carcinoma of Breast|8530/3
C0278601|T191|SY|C4001|NCI|Inflammatory Carcinoma of the Breast|8530/3
C0278601|T191|SY|C4001|NCI|Mastitis Carcinomatosa|8530/3
C0278601|T191|PT|10021980|NCI_CTEP-SDC|Inflammatory breast carcinoma|8530/3
C0278601|T191|DN|C4001|NCI_CTRP|Inflammatory Breast Cancer|8530/3
C0278601|T191|PT|CDR0000045313|NCI_NCI-GLOSS|inflammatory breast cancer|8530/3
C0278601|T191|SY|CDR0000040816|PDQ|breast cancer, inflammatory|8530/3
C0278601|T191|SY|CDR0000040816|PDQ|carcinoma of the breast, inflammatory|8530/3
C0278601|T191|PSC|CDR0000040816|PDQ|inflammatory breast cancer|8530/3
C0334385|T191|SY|BB9H.|RCD|Inflammatory adenocarcinoma|8530/3
C0334385|T191|PT|BB9H.|RCD|Inflammatory carcinoma|8530/3
C0278601|T191|AB|X78WP|RCD|Inflammatory carcinoma breast|8530/3
C0278601|T191|PT|X78WP|RCD|Inflammatory carcinoma of breast|8530/3
C0278601|T191|SY|X78WP|RCD|Mastitis carcinomatosa|8530/3
C0334385|T191|SY|32968003|SNOMEDCT_US|Inflammatory adenocarcinoma|8530/3
C0334385|T191|PT|32968003|SNOMEDCT_US|Inflammatory carcinoma|8530/3
C0278601|T191|PT|254840009|SNOMEDCT_US|Inflammatory carcinoma of breast|8530/3
C0278601|T191|SY|254840009|SNOMEDCT_US|Mastitis carcinomatosa|8530/3
C0030185|T191|PT|0024219|CCPSS|PAGET DISEASE MAMMARY|8540/3
C0030185|T191|SY|0000009182|CHV|breast disease paget|8540/3
C0030185|T191|SY|0000009182|CHV|breast disease paget's|8540/3
C0030185|T191|SY|0000009182|CHV|breast disease pagets|8540/3
C0030185|T191|SY|0000009182|CHV|breast diseases paget|8540/3
C0030185|T191|SY|0000009182|CHV|breast diseases pagets|8540/3
C0030185|T191|SY|0000009182|CHV|breast paget disease|8540/3
C0030185|T191|SY|0000009182|CHV|breast paget's disease|8540/3
C0030185|T191|SY|0000009182|CHV|breast pagets disease|8540/3
C0030185|T191|SY|0000009182|CHV|disease nipple paget|8540/3
C0030185|T191|SY|0000009182|CHV|disease nipple pagets|8540/3
C0030185|T191|SY|0000009182|CHV|disease nipples paget|8540/3
C0030185|T191|SY|0000009182|CHV|disease nipples paget's|8540/3
C0030185|T191|SY|0000009182|CHV|mammary paget disease|8540/3
C0030185|T191|SY|0000009182|CHV|mammary paget's disease|8540/3
C0030185|T191|SY|0000009182|CHV|paget disease breast|8540/3
C0030185|T191|SY|0000009182|CHV|paget disease of breast|8540/3
C0030185|T191|SY|0000009182|CHV|paget's breast disease|8540/3
C0030185|T191|SY|0000009182|CHV|paget's disease breast|8540/3
C0030185|T191|SY|0000009182|CHV|paget's disease mammary|8540/3
C0030185|T191|SY|0000009182|CHV|paget's disease of breast|8540/3
C0030185|T191|SY|0000009182|CHV|paget's disease of nipple|8540/3
C0030185|T191|PT|0000009182|CHV|paget's disease of the breast|8540/3
C0030185|T191|SY|0000009182|CHV|paget's disease of the nipple|8540/3
C0030185|T191|SY|0000009182|CHV|pagets breast disease|8540/3
C0030185|T191|SY|0000009182|CHV|pagets disease breast|8540/3
C0030185|T191|PT|NOCODE|COSTAR|Paget's Disease of Breast|8540/3
C0030185|T191|PT|2000-8560|CSP|Paget's disease of breast|8540/3
C0030185|T191|DI|U001377|DXP|PAGET DISEASE, BREAST|8540/3
C0030185|T191|ET|C50|ICD10CM|Paget's disease of breast|8540/3
C0030185|T191|PT|MTHU047359|ICPC2ICD10ENG|breast; disorder, Paget|8540/3
C0030185|T191|PT|MTHU047461|ICPC2ICD10ENG|breast; Paget|8540/3
C0030185|T191|PT|MTHU057029|ICPC2ICD10ENG|Paget; breast|8540/3
C0030185|T191|LLT|10033367|MDR|Paget's disease of the breast|8540/3
C0030185|T191|PT|31658|MEDCIN|Paget's disease of breast|8540/3
C0030185|T191|ET|3|MEDLINEPLUS|Paget's Disease of Breast|8540/3
C0030185|T191|PM|D010144|MSH|Disease, Mammary Paget|8540/3
C0030185|T191|PM|D010144|MSH|Disease, Mammary Paget's|8540/3
C0030185|T191|DEV|D010144|MSH|MAMMARY PAGET DIS|8540/3
C0030185|T191|ET|D010144|MSH|Mammary Paget Disease|8540/3
C0030185|T191|ET|D010144|MSH|Mammary Paget's Disease|8540/3
C0030185|T191|DEV|D010144|MSH|MAMMARY PAGETS DIS|8540/3
C0030185|T191|PM|D010144|MSH|Mammary Pagets Disease|8540/3
C0030185|T191|DEV|D010144|MSH|PAGET DIS BREAST|8540/3
C0030185|T191|DEV|D010144|MSH|PAGET DIS MAMMARY|8540/3
C0030185|T191|ET|D010144|MSH|Paget Disease of Breast|8540/3
C0030185|T191|PM|D010144|MSH|Paget Disease, Breast|8540/3
C0030185|T191|ET|D010144|MSH|Paget Disease, Mammary|8540/3
C0030185|T191|ET|D010144|MSH|Paget's Disease of Breast|8540/3
C0030185|T191|ET|D010144|MSH|Paget's Disease of the Breast|8540/3
C0030185|T191|ET|D010144|MSH|Paget's Disease of the Nipple|8540/3
C0030185|T191|ET|D010144|MSH|Paget's Disease of the Nipple and Areola|8540/3
C0030185|T191|MH|D010144|MSH|Paget's Disease, Mammary|8540/3
C0030185|T191|DEV|D010144|MSH|PAGETS DIS BREAST|8540/3
C0030185|T191|DEV|D010144|MSH|PAGETS DIS MAMMARY|8540/3
C0030185|T191|PM|D010144|MSH|Pagets Disease, Breast|8540/3
C0030185|T191|PM|D010144|MSH|Pagets Disease, Mammary|8540/3
C0030185|T191|ET|D010144|MSH|Pigmented Mammary Paget Disease|8540/3
C0030185|T191|PN|NOCODE|MTH|Paget's Disease, Mammary|8540/3
C0030185|T191|SY|C47857|NCI|Mammary Paget's Disease|8540/3
C0030185|T191|PT|C47857|NCI|Paget Disease of the Breast|8540/3
C0030185|T191|SY|C47857|NCI|Paget's Disease of Breast|8540/3
C0030185|T191|SY|C47857|NCI|Paget's Disease of the Breast|8540/3
C0030185|T191|DN|C47857|NCI_CTRP|Paget Disease of the Breast|8540/3
C0030185|T191|SY|CDR0000039851|PDQ|mammary paget's disease|8540/3
C0030185|T191|PT|CDR0000039851|PDQ|Paget disease of the breast|8540/3
C0030185|T191|SY|CDR0000039851|PDQ|Paget's disease of breast|8540/3
C0030185|T191|LV|CDR0000039851|PDQ|Paget's disease of the breast|8540/3
C0030185|T191|PT|BB9J.|RCD|Mammary Paget's disease|8540/3
C0030185|T191|SY|BB9J.|RCD|Paget's disease of breast|8540/3
C0030185|T191|SY|2985005|SNOMEDCT_US|Mammary Paget's disease|8540/3
C0030185|T191|SY|2985005|SNOMEDCT_US|Paget disease, mammary|8540/3
C0030185|T191|SY|2985005|SNOMEDCT_US|Paget's disease of breast|8540/3
C0030185|T191|PT|2985005|SNOMEDCT_US|Paget's disease, mammary|8540/3
C0334386|T191|PT|232389|MEDCIN|Paget's disease and infiltrating duct carcinoma of breast|8541/3
C0279567|T191|PT|C7951|NCI|Paget Disease of the Breast with Invasive Ductal Carcinoma|8541/3
C0279567|T191|SY|C7951|NCI|Paget's Disease and Infiltrating Ductal Carcinoma of Breast|8541/3
C0279567|T191|SY|C7951|NCI|Paget's Disease and Infiltrating Ductal Carcinoma of the Breast|8541/3
C0279567|T191|SY|C7951|NCI|Paget's Disease and Invasive Ductal Carcinoma of Breast|8541/3
C0279567|T191|SY|C7951|NCI|Paget's Disease and Invasive Ductal Carcinoma of the Breast|8541/3
C0279567|T191|SY|C7951|NCI|Paget's Disease of Breast with Infiltrating Ductal Carcinoma|8541/3
C0279567|T191|SY|C7951|NCI|Paget's Disease of Breast with Invasive Ductal Carcinoma|8541/3
C0279567|T191|SY|C7951|NCI|Paget's Disease of the Breast with Infiltrating Ductal Carcinoma|8541/3
C0279567|T191|SY|C7951|NCI|Paget's Disease of the Breast with Invasive Ductal Carcinoma|8541/3
C0279567|T191|DN|C7951|NCI_CTRP|Paget Disease of the Breast with Invasive Ductal Carcinoma|8541/3
C0279567|T191|PT|CDR0000039853|PDQ|Paget disease of the breast with invasive ductal carcinoma|8541/3
C0279567|T191|SY|CDR0000039853|PDQ|Paget's disease and infiltrating ductal carcinoma of breast|8541/3
C0279567|T191|SY|CDR0000039853|PDQ|Paget's disease and infiltrating ductal carcinoma of the breast|8541/3
C0279567|T191|SY|CDR0000039853|PDQ|Paget's disease and invasive ductal carcinoma of breast|8541/3
C0279567|T191|SY|CDR0000039853|PDQ|Paget's disease and invasive ductal carcinoma of the breast|8541/3
C0279567|T191|SY|CDR0000039853|PDQ|Paget's disease of breast with infiltrating ductal carcinoma|8541/3
C0279567|T191|SY|CDR0000039853|PDQ|Paget's disease of breast with invasive ductal carcinoma|8541/3
C0279567|T191|SY|CDR0000039853|PDQ|Paget's disease of the breast with infiltrating ductal carcinoma|8541/3
C0279567|T191|SY|CDR0000039853|PDQ|Paget's disease of the breast with invasive ductal carcinoma|8541/3
C0334386|T191|PT|BB9K.|RCD|Paget's disease and infiltrating duct carcinoma of breast|8541/3
C0334386|T191|AB|BB9K.|RCD|Paget's+infiltr duct ca breast|8541/3
C0334386|T191|SY|82591005|SNOMEDCT_US|Paget disease and infiltrating duct carcinoma of breast|8541/3
C0334386|T191|PT|82591005|SNOMEDCT_US|Paget's disease and infiltrating duct carcinoma of breast|8541/3
C0030186|T191|SY|0000032319|CHV|diseases paget's skin|8542/3
C0030186|T191|SY|0000009183|CHV|extra mammary paget's disease|8542/3
C0030186|T191|SY|0000009183|CHV|extra-mammary paget's disease|8542/3
C0030186|T191|SY|0000009183|CHV|extra-mammary pagets disease|8542/3
C0030186|T191|SY|0000009183|CHV|extramammary paget disease|8542/3
C0030186|T191|PT|0000009183|CHV|extramammary paget's disease|8542/3
C0030186|T191|SY|0000009183|CHV|extramammary pagets disease|8542/3
C0030186|T191|SY|0000009183|CHV|paget's disease extramammary|8542/3
C0030186|T191|SY|0000032319|CHV|paget's disease of skin|8542/3
C0030186|T191|PT|0000032319|CHV|paget's skin disease|8542/3
C0030186|T191|DI|U001378|DXP|PAGET DISEASE, EXTRAMAMMARY|8542/3
C0030186|T191|PT|10068223|MDR|Extramammary Paget's disease|8542/3
C0030186|T191|LLT|10068223|MDR|Extramammary Paget's disease|8542/3
C0030186|T191|LLT|10033366|MDR|Paget's disease of skin|8542/3
C0030186|T191|PT|31702|MEDCIN|extramammary Paget's disease|8542/3
C0030186|T191|DEV|D010145|MSH|EXTRA MAMMARY PAGET DIS|8542/3
C0030186|T191|PM|D010145|MSH|Extra Mammary Paget Disease|8542/3
C0030186|T191|PM|D010145|MSH|Extra Mammary Paget's Disease|8542/3
C0030186|T191|DEV|D010145|MSH|EXTRA MAMMARY PAGETS DIS|8542/3
C0030186|T191|ET|D010145|MSH|Extra-Mammary Paget Disease|8542/3
C0030186|T191|ET|D010145|MSH|Extra-Mammary Paget's Disease|8542/3
C0030186|T191|PM|D010145|MSH|Extra-Mammary Pagets Disease|8542/3
C0030186|T191|DEV|D010145|MSH|EXTRAMAMMARY PAGET DIS|8542/3
C0030186|T191|ET|D010145|MSH|Extramammary Paget Disease|8542/3
C0030186|T191|ET|D010145|MSH|Extramammary Paget's Disease|8542/3
C0030186|T191|DEV|D010145|MSH|EXTRAMAMMARY PAGETS DIS|8542/3
C0030186|T191|PM|D010145|MSH|Extramammary Pagets Disease|8542/3
C0030186|T191|PM|D010145|MSH|Extramammary, Paget Disease|8542/3
C0030186|T191|DEV|D010145|MSH|PAGET DIS EXTRA MAMMARY|8542/3
C0030186|T191|DEV|D010145|MSH|PAGET DIS EXTRAMAMMARY|8542/3
C0030186|T191|ET|D010145|MSH|Paget Disease Extramammary|8542/3
C0030186|T191|PM|D010145|MSH|Paget Disease, Extra Mammary|8542/3
C0030186|T191|ET|D010145|MSH|Paget Disease, Extra-Mammary|8542/3
C0030186|T191|MH|D010145|MSH|Paget Disease, Extramammary|8542/3
C0030186|T191|PM|D010145|MSH|Paget's Disease, Extra Mammary|8542/3
C0030186|T191|ET|D010145|MSH|Paget's Disease, Extra-Mammary|8542/3
C0030186|T191|ET|D010145|MSH|Paget's Disease, Extramammary|8542/3
C0030186|T191|DEV|D010145|MSH|PAGETS DIS EXTRA MAMMARY|8542/3
C0030186|T191|DEV|D010145|MSH|PAGETS DIS EXTRAMAMMARY|8542/3
C0030186|T191|PM|D010145|MSH|Pagets Disease, Extra-Mammary|8542/3
C0030186|T191|PM|D010145|MSH|Pagets Disease, Extramammary|8542/3
C0030186|T191|PN|NOCODE|MTH|Paget Disease Extramammary|8542/3
C0030186|T191|SY|C3302|NCI|Cutaneous Paget's Disease|8542/3
C0030186|T191|PT|C3302|NCI|Extramammary Paget Disease|8542/3
C0030186|T191|SY|C3302|NCI|Extramammary Paget's Disease|8542/3
C0030186|T191|SY|C3302|NCI|Paget Disease Extramammary|8542/3
C0030186|T191|SY|C3302|NCI|Paget's Disease of Skin|8542/3
C0030186|T191|SY|C3302|NCI|Paget's Disease of the Skin|8542/3
C0030186|T191|SY|C3302|NCI|Paget's Skin Disease|8542/3
C0030186|T191|PT|Xa98z|RCD|Extramammary Paget's disease|8542/3
C0030186|T191|PT|X00kl|RCD|Paget's disease of skin|8542/3
C0030186|T191|OA|BB9L.|RCDSY|Paget's dis ex-mamm ex bone|8542/3
C0030186|T191|OA|BB9L.|RCDSY|Paget's disease, extramammary, exc Paget's disease bone|8542/3
C0030186|T191|OP|BB9L.|RCDSY|Paget's disease, extramammary, excluding Paget's disease of bone|8542/3
C0030186|T191|OAP|302830004|SNOMEDCT_US|Extramammary Paget's disease|8542/3
C0030186|T191|SY|232336001|SNOMEDCT_US|Paget disease of skin|8542/3
C0030186|T191|PT|232336001|SNOMEDCT_US|Paget's disease of skin|8542/3
C0279566|T191|PT|232390|MEDCIN|Paget's disease and intraductal carcinoma of breast|8543/3
C0279566|T191|PT|C4019|NCI|Paget Disease and Intraductal Carcinoma of the Breast|8543/3
C0279566|T191|SY|C4019|NCI|Paget's Disease and Intraductal Carcinoma of Breast|8543/3
C0279566|T191|SY|C4019|NCI|Paget's Disease and Intraductal Carcinoma of the Breast|8543/3
C0279566|T191|SY|C4019|NCI|Paget's Disease of Breast with Intraductal Carcinoma|8543/3
C0279566|T191|SY|C4019|NCI|Paget's Disease of the Breast with Intraductal Carcinoma|8543/3
C0279566|T191|DN|C4019|NCI_CTRP|Paget Disease and Intraductal Carcinoma of the Breast|8543/3
C0279566|T191|SY|CDR0000039852|PDQ|Paget disease and intraductal carcinoma of the breast|8543/3
C0279566|T191|PT|CDR0000039852|PDQ|Paget disease of the breast with intraductal carcinoma|8543/3
C0279566|T191|SY|CDR0000039852|PDQ|Paget's disease and intraductal carcinoma of breast|8543/3
C0279566|T191|SY|CDR0000039852|PDQ|Paget's disease and intraductal carcinoma of the breast|8543/3
C0279566|T191|SY|CDR0000039852|PDQ|Paget's disease of breast with intraductal carcinoma|8543/3
C0279566|T191|LV|CDR0000039852|PDQ|Paget's Disease of the Breast with Intraductal Carcinoma|8543/3
C0279566|T191|PT|X77ny|RCD|Paget's disease and intraductal carcinoma of breast|8543/3
C0279566|T191|AB|X77ny|RCD|Paget's+intraductal ca breast|8543/3
C0279566|T191|AB|X77ny|RCDSY|Pagets+intradc carc breast|8543/3
C0279566|T191|SY|54666007|SNOMEDCT_US|Paget disease and intraductal carcinoma of breast|8543/3
C0279566|T191|PT|54666007|SNOMEDCT_US|Paget's disease and intraductal carcinoma of breast|8543/3
C0279566|T191|OAP|189714001|SNOMEDCT_US|Paget's disease and intraductal carcinoma of breast|8543/3
C0279566|T191|OF|189714001|SNOMEDCT_US|Paget's disease and intraductal carcinoma of breast|8543/3
C0334389|T191|PN|NOCODE|MTH|Acinar cell adenoma|8550/0
C0334389|T191|SY|C4196|NCI|Acinar Adenoma|8550/0
C0334389|T191|PT|C4196|NCI|Acinar Cell Adenoma|8550/0
C0334389|T191|SY|C4196|NCI|Acinic Cell Adenoma|8550/0
C0334389|T191|SY|C4196|NCI_CDISC|Acinar Adenoma|8550/0
C0334389|T191|SY|C4196|NCI_CDISC|Acinic Cell Adenoma|8550/0
C0334389|T191|PT|C4196|NCI_CDISC|ADENOMA, ACINAR CELL, BENIGN|8550/0
C0334389|T191|SY|BBA0.|RCD|Acinar adenoma|8550/0
C0334389|T191|PT|BBA0.|RCD|Acinar cell adenoma|8550/0
C0334389|T191|SY|BBA0.|RCD|Acinic cell adenoma|8550/0
C0334389|T191|SY|79041005|SNOMEDCT_US|Acinar adenoma|8550/0
C0334389|T191|PT|79041005|SNOMEDCT_US|Acinar cell adenoma|8550/0
C0334389|T191|SY|79041005|SNOMEDCT_US|Acinic cell adenoma|8550/0
C0334390|T191|PT|0000029970|CHV|acinar cell tumor|8550/1
C0334390|T191|SY|0000029970|CHV|acinic cell tumor|8550/1
C0334390|T191|PT|MTHU002964|ICPC2ICD10ENG|acinic cell; tumor|8550/1
C0334390|T191|PT|MTHU077008|ICPC2ICD10ENG|tumor; acinic cell|8550/1
C0334390|T191|PN|NOCODE|MTH|Acinar cell tumor|8550/1
C0334390|T191|PT|C4197|NCI|Acinar Cell Neoplasm|8550/1
C0334390|T191|SY|C4197|NCI|Acinar Cell Tumor|8550/1
C0334390|T191|PT|Xa990|RCD|Acinar cell tumour|8550/1
C0334390|T191|PT|Xa990|RCDAE|Acinar cell tumor|8550/1
C0334390|T191|OP|BBA1.|RCDSA|Acinar cell tumor|8550/1
C0334390|T191|OP|BBAz.|RCDSY|Acinar cell neoplasm NOS|8550/1
C0334390|T191|OP|BBA..|RCDSY|Acinar cell neoplasms|8550/1
C0334390|T191|OP|BBA1.|RCDSY|Acinar cell tumour|8550/1
C0334390|T191|PT|115219005|SNOMEDCT_US|Acinar cell neoplasm|8550/1
C0334390|T191|OAP|83472001|SNOMEDCT_US|Acinar cell tumor|8550/1
C0334390|T191|OAP|83472001|SNOMEDCT_US|Acinar cell tumour|8550/1
C0334390|T191|OAS|83472001|SNOMEDCT_US|Acinic cell tumor|8550/1
C0334390|T191|OAS|83472001|SNOMEDCT_US|Acinic cell tumour|8550/1
C0206685|T191|SY|0000021019|CHV|acinar adenocarcinoma|8550/3
C0206685|T191|PT|0000021019|CHV|acinar carcinoma|8550/3
C0206685|T191|SY|0000021019|CHV|acinar cell carcinoma|8550/3
C0206685|T191|LLT|10064646|MDR|Acinic cell carcinoma|8550/3
C0206685|T191|PT|271444|MEDCIN|acinar cell carcinoma|8550/3
C0206685|T191|ET|D018267|MSH|Acinar Carcinoma|8550/3
C0206685|T191|PM|D018267|MSH|Acinar Carcinomas|8550/3
C0206685|T191|ET|D018267|MSH|Acinar Cell Adenocarcinoma|8550/3
C0206685|T191|PM|D018267|MSH|Acinar Cell Adenocarcinomas|8550/3
C0206685|T191|PM|D018267|MSH|Acinar Cell Carcinoma|8550/3
C0206685|T191|PM|D018267|MSH|Acinar Cell Carcinomas|8550/3
C0206685|T191|ET|D018267|MSH|Acinic Cell Adenocarcinoma|8550/3
C0206685|T191|PM|D018267|MSH|Acinic Cell Adenocarcinomas|8550/3
C0206685|T191|ET|D018267|MSH|Acinic Cell Carcinoma|8550/3
C0206685|T191|PM|D018267|MSH|Acinic Cell Carcinomas|8550/3
C0206685|T191|ET|D018267|MSH|Acinic Cell Tumor|8550/3
C0206685|T191|PM|D018267|MSH|Acinic Cell Tumors|8550/3
C0206685|T191|PM|D018267|MSH|Adenocarcinoma, Acinar Cell|8550/3
C0206685|T191|PM|D018267|MSH|Adenocarcinoma, Acinic Cell|8550/3
C0206685|T191|PM|D018267|MSH|Adenocarcinomas, Acinar Cell|8550/3
C0206685|T191|PM|D018267|MSH|Adenocarcinomas, Acinic Cell|8550/3
C0206685|T191|PM|D018267|MSH|Carcinoma, Acinar|8550/3
C0206685|T191|MH|D018267|MSH|Carcinoma, Acinar Cell|8550/3
C0206685|T191|PM|D018267|MSH|Carcinoma, Acinic Cell|8550/3
C0206685|T191|PM|D018267|MSH|Carcinomas, Acinar|8550/3
C0206685|T191|PM|D018267|MSH|Carcinomas, Acinar Cell|8550/3
C0206685|T191|PM|D018267|MSH|Carcinomas, Acinic Cell|8550/3
C0206685|T191|PM|D018267|MSH|Tumor, Acinic Cell|8550/3
C0206685|T191|PM|D018267|MSH|Tumors, Acinic Cell|8550/3
C0206685|T191|PN|NOCODE|MTH|Acinar Cell Carcinoma|8550/3
C0206685|T191|SY|C3768|NCI|Acinar Adenocarcinoma|8550/3
C0206685|T191|SY|C3768|NCI|Acinar Carcinoma|8550/3
C0206685|T191|SY|C3768|NCI|Acinar Cell Adenocarcinoma|8550/3
C0206685|T191|SY|TCGA|NCI|Acinar Cell Carcinoma|8550/3
C0206685|T191|PT|C3768|NCI|Acinar Cell Carcinoma|8550/3
C0206685|T191|SY|C3768|NCI|Acinic Cell Adenocarcinoma|8550/3
C0206685|T191|SY|C3768|NCI|Acinic Cell Carcinoma|8550/3
C0206685|T191|SY|C3768|NCI_CDISC|Acinar Adenocarcinoma|8550/3
C0206685|T191|SY|C3768|NCI_CDISC|Acinar Carcinoma|8550/3
C0206685|T191|SY|C3768|NCI_CDISC|Acinar Cell Adenocarcinoma|8550/3
C0206685|T191|SY|C3768|NCI_CDISC|Acinic Cell Adenocarcinoma|8550/3
C0206685|T191|SY|C3768|NCI_CDISC|Acinic Cell Carcinoma|8550/3
C0206685|T191|PT|C3768|NCI_CDISC|CARCINOMA, ACINAR CELL, MALIGNANT|8550/3
C0206685|T191|SY|BBA2.|RCD|Acinar adenocarcinoma|8550/3
C0206685|T191|SY|BBA2.|RCD|Acinar carcinoma|8550/3
C0206685|T191|PT|BBA2.|RCD|Acinar cell carcinoma|8550/3
C0206685|T191|SY|BBA2.|RCD|Acinic cell adenocarcinoma|8550/3
C0206685|T191|SY|45410002|SNOMEDCT_US|Acinar adenocarcinoma|8550/3
C0206685|T191|SY|45410002|SNOMEDCT_US|Acinar carcinoma|8550/3
C0206685|T191|PT|45410002|SNOMEDCT_US|Acinar cell carcinoma|8550/3
C0206685|T191|SY|45410002|SNOMEDCT_US|Acinic cell adenocarcinoma|8550/3
C1266087|T191|PT|271445|MEDCIN|acinar cell cystadenocarcinoma|8551/3
C1266087|T191|PT|38723|MEDCIN|acinar cell cystadenocarcinoma of pancreas|8551/3
C1266087|T191|SY|C5727|NCI|Acinar Cell Cystadenocarcinoma|8551/3
C1266087|T191|SY|C3874|NCI|Acinar Cell Cystadenocarcinoma|8551/3
C1266087|T191|SY|C5727|NCI|Acinar Cell Cystadenocarcinoma of Pancreas|8551/3
C1266087|T191|SY|C5727|NCI|Acinar Cell Cystadenocarcinoma of the Pancreas|8551/3
C1266087|T191|PT|C5727|NCI|Pancreatic Acinar Cell Cystadenocarcinoma|8551/3
C1266087|T191|SY|TCGA|NCI|Pancreatic Acinar Cell Cystadenocarcinoma|8551/3
C1266087|T191|PT|128703004|SNOMEDCT_US|Acinar cell cystadenocarcinoma|8551/3
C4518208|T191|PT|733855008|SNOMEDCT_US|Acinar cell cystadenoma|8551/3
C2987160|T191|PT|C95458|NCI|Mixed Acinar-Ductal Carcinoma of the Pancreas|8552/3
C3472609|T191|PT|450897002|SNOMEDCT_US|Mixed acinar-ductal carcinoma|8552/3
C1314684|T191|PN|NOCODE|MTH|Mixed squamous cell and glandular papilloma|8560/0
C1708774|T191|SY|C45602|NCI|Lung Mixed Squamous and Glandular Papilloma|8560/0
C1708774|T191|PT|C45602|NCI|Lung Mixed Squamous Cell and Glandular Papilloma|8560/0
C1314684|T191|PT|107692003|SNOMEDCT_US|Mixed squamous cell and glandular papilloma|8560/0
C0206623|T191|PT|0034009|CCPSS|ADENOSQUAMOUS CARCINOMA|8560/3
C0206623|T191|LA|LA15446-0|LNC|Adenosquamous carcinoma|8560/3
C0206623|T191|PT|10068873|MDR|Adenosquamous cell carcinoma|8560/3
C0206623|T191|LLT|10068873|MDR|Adenosquamous cell carcinoma|8560/3
C0206623|T191|PT|271446|MEDCIN|adenosquamous carcinoma|8560/3
C0206623|T191|PM|D018196|MSH|Adenosquamous Carcinoma|8560/3
C0206623|T191|PM|D018196|MSH|Adenosquamous Carcinomas|8560/3
C0206623|T191|MH|D018196|MSH|Carcinoma, Adenosquamous|8560/3
C0206623|T191|PM|D018196|MSH|Carcinomas, Adenosquamous|8560/3
C0206623|T191|PN|NOCODE|MTH|Adenosquamous carcinoma|8560/3
C0206623|T191|SY|TCGA|NCI|Adenosquamous Carcinoma|8560/3
C0206623|T191|PT|C3727|NCI|Adenosquamous Carcinoma|8560/3
C0206623|T191|SY|C3727|NCI|Mixed Adenocarcinoma and Epidermoid Carcinoma|8560/3
C0206623|T191|SY|C3727|NCI|Mixed Adenocarcinoma and Epidermoid Cell Carcinoma|8560/3
C0206623|T191|SY|C3727|NCI|Mixed Adenocarcinoma and Squamous Carcinoma|8560/3
C0206623|T191|SY|C3727|NCI|Mixed Adenocarcinoma and Squamous Cell Carcinoma|8560/3
C0206623|T191|PT|C3727|NCI_CDISC|CARCINOMA, ADENOSQUAMOUS, MALIGNANT|8560/3
C0206623|T191|SY|C3727|NCI_CDISC|Mixed Adenocarcinoma and Epidermoid Carcinoma|8560/3
C0206623|T191|SY|C3727|NCI_CDISC|Mixed Adenocarcinoma and Epidermoid Cell Carcinoma|8560/3
C0206623|T191|SY|C3727|NCI_CDISC|Mixed Adenocarcinoma and Squamous Carcinoma|8560/3
C0206623|T191|SY|C3727|NCI_CDISC|Mixed Adenocarcinoma and Squamous Cell Carcinoma|8560/3
C0206623|T191|PT|C3727|NCI_CPTAC|Adenosquamous Carcinoma|8560/3
C0206623|T191|PT|CDR0000476766|NCI_NCI-GLOSS|adenosquamous carcinoma|8560/3
C0206623|T191|PT|BBB0.|RCD|Adenosquamous carcinoma|8560/3
C0206623|T191|AB|BBB0.|RCD|Mixed adenoca+epidermoid ca|8560/3
C0206623|T191|AB|BBB0.|RCD|Mixed adenoca+squamous cell ca|8560/3
C0206623|T191|SY|BBB0.|RCD|Mixed adenocarcinoma and epidermoid carcinoma|8560/3
C0206623|T191|SY|BBB0.|RCD|Mixed adenocarcinoma and squamous cell carcinoma|8560/3
C0206623|T191|SY|403902008|SNOMEDCT_US|Adenosquamous carcinoma|8560/3
C0206623|T191|PT|59367005|SNOMEDCT_US|Adenosquamous carcinoma|8560/3
C0206623|T191|PT|403902008|SNOMEDCT_US|Adenosquamous cell carcinoma|8560/3
C0206623|T191|SY|59367005|SNOMEDCT_US|Mixed adenocarcinoma and epidermoid carcinoma|8560/3
C0206623|T191|SY|59367005|SNOMEDCT_US|Mixed adenocarcinoma and squamous cell carcinoma|8560/3
C0001429|T191|SY|0000000715|CHV|adenolymphoma|8561/0
C0001429|T191|SY|0000031263|CHV|tumor warthin's|8561/0
C0001429|T191|SY|0000000715|CHV|tumor warthin's|8561/0
C0001429|T191|SY|0000000715|CHV|tumor warthins|8561/0
C0001429|T191|SY|0000031263|CHV|tumors warthin's|8561/0
C0001429|T191|SY|0000000715|CHV|tumors warthin's|8561/0
C0001429|T191|SY|0000000715|CHV|warthin tumor|8561/0
C0001429|T191|PT|0000000715|CHV|warthin's tumor|8561/0
C0001429|T191|PT|0000031263|CHV|warthin's tumor|8561/0
C0001429|T191|SY|0000031263|CHV|warthin's tumour|8561/0
C0001429|T191|SY|0000000715|CHV|warthin's tumour|8561/0
C0001429|T191|PT|U000066|LCH|Adenolymphoma|8561/0
C0001429|T191|PT|sh85000842|LCH_NW|Adenolymphoma|8561/0
C0001429|T191|PT|10070460|MDR|Adenolymphoma|8561/0
C0001429|T191|LLT|10070460|MDR|Adenolymphoma|8561/0
C0001429|T191|LLT|10074291|MDR|Papillary cystadenoma lymphomatosum|8561/0
C0001429|T191|PT|10074291|MDR|Papillary cystadenoma lymphomatosum|8561/0
C0001429|T191|LLT|10074288|MDR|Warthin's tumor|8561/0
C0001429|T191|LLT|10074292|MDR|Warthin's tumour|8561/0
C0001429|T191|MH|D000235|MSH|Adenolymphoma|8561/0
C0001429|T191|PM|D000235|MSH|Adenolymphomas|8561/0
C0001429|T191|ET|D000235|MSH|Cystadenoma Lymphomatosum, Papillary|8561/0
C0001429|T191|PM|D000235|MSH|Papillary Cystadenoma Lymphomatosum|8561/0
C0001429|T191|PM|D000235|MSH|Tumor, Warthin|8561/0
C0001429|T191|ET|D000235|MSH|Warthin Tumor|8561/0
C0001429|T191|PN|NOCODE|MTH|Adenolymphoma|8561/0
C0001429|T191|SY|C2854|NCI|Adenolymphoma|8561/0
C0001429|T191|SY|C2854|NCI|Papillary Cystadenoma Lymphomatosum|8561/0
C0001429|T191|PT|C2854|NCI|Warthin Tumor|8561/0
C0001429|T191|SY|C2854|NCI|Warthin's Tumor|8561/0
C0001429|T191|PT|BBB1.|RCD|Adenolymphoma|8561/0
C0001429|T191|AB|BBB1.|RCD|Papill cystadenoma lymphomatos|8561/0
C0001429|T191|SY|BBB1.|RCD|Papillary cystadenoma lymphomatosum|8561/0
C0001429|T191|PT|422470007|SNOMEDCT_US|Adenolymphoma|8561/0
C0001429|T191|PT|20776008|SNOMEDCT_US|Adenolymphoma|8561/0
C0001429|T191|SY|422470007|SNOMEDCT_US|Papillary cystadenoma lymphomatosum|8561/0
C0001429|T191|SY|20776008|SNOMEDCT_US|Papillary cystadenoma lymphomatosum|8561/0
C0001429|T191|SY|422470007|SNOMEDCT_US|Warthin's tumor|8561/0
C0001429|T191|SY|20776008|SNOMEDCT_US|Warthin's tumor|8561/0
C0001429|T191|SYGB|422470007|SNOMEDCT_US|Warthin's tumour|8561/0
C0001429|T191|SYGB|20776008|SNOMEDCT_US|Warthin's tumour|8561/0
C0334392|T191|PT|271447|MEDCIN|epithelial-myoepithelial carcinoma|8562/3
C0334392|T191|PT|C4199|NCI|Epithelial-Myoepithelial Carcinoma|8562/3
C0334392|T191|PT|C4199|NCI_CPTAC|Epithelial-Myoepithelial Carcinoma|8562/3
C0334392|T191|AB|X77o1|RCD|Epithelial-myoepithelial ca|8562/3
C0334392|T191|PT|X77o1|RCD|Epithelial-myoepithelial carcinoma|8562/3
C0334392|T191|AB|X77o1|RCDSY|Epith-myoepithel carcinoma|8562/3
C0334392|T191|OF|189722008|SNOMEDCT_US|Epithelial-myoepithelial carcinoma|8562/3
C0334392|T191|PT|9618003|SNOMEDCT_US|Epithelial-myoepithelial carcinoma|8562/3
C0334392|T191|OAP|189722008|SNOMEDCT_US|Epithelial-myoepithelial carcinoma|8562/3
C0334393|T191|PT|271467|MEDCIN|adenocarcinoma with squamous metaplasia|8570/3
C0334393|T191|PN|NOCODE|MTH|Adenocarcinoma with squamous metaplasia|8570/3
C0334393|T191|SY|C4200|NCI|Adenoacanthoma|8570/3
C0334393|T191|PT|C4200|NCI|Adenocarcinoma with Squamous Metaplasia|8570/3
C0334393|T191|SY|TCGA|NCI|Adenocarcinoma with Squamous Metaplasia|8570/3
C0334393|T191|SY|C4200|NCI_CDISC|Adenoacanthoma|8570/3
C0334393|T191|PT|C4200|NCI_CDISC|ADENOACANTHOMA, MALIGNANT|8570/3
C0334393|T191|SY|BBB2.|RCD|Adenoacanthoma|8570/3
C0334393|T191|AB|BBB2.|RCD|Adenoca + squamous metaplasia|8570/3
C0334393|T191|PT|BBB2.|RCD|Adenocarcinoma with squamous metaplasia|8570/3
C0334393|T191|SY|15176003|SNOMEDCT_US|Adenoacanthoma|8570/3
C0334393|T191|PT|15176003|SNOMEDCT_US|Adenocarcinoma with squamous metaplasia|8570/3
C0334394|T191|PT|271468|MEDCIN|adenocarcinoma with cartilaginous and osseous metaplasia|8571/3
C0334394|T191|PT|C7683|NCI|Adenocarcinoma with Cartilaginous and Osseous Metaplasia|8571/3
C0334394|T191|SY|TCGA|NCI|Adenocarcinoma with Cartilaginous and Osseous Metaplasia|8571/3
C0334394|T191|AB|BBB3.|RCD|Adenoca+cartil+osseous metapl|8571/3
C0334394|T191|PT|BBB3.|RCD|Adenocarcinoma with cartilaginous and osseous metaplasia|8571/3
C0334394|T191|PT|56484001|SNOMEDCT_US|Adenocarcinoma with cartilaginous and osseous metaplasia|8571/3
C0334395|T191|PT|271469|MEDCIN|adenocarcinoma with spindle cell metaplasia|8572/3
C0334395|T191|PT|C4201|NCI|Adenocarcinoma with Spindle Cell Metaplasia|8572/3
C0334395|T191|SY|TCGA|NCI|Adenocarcinoma with Spindle Cell Metaplasia|8572/3
C0334395|T191|AB|BBB4.|RCD|Adenoca+spindle cell metaplas|8572/3
C0334395|T191|PT|BBB4.|RCD|Adenocarcinoma with spindle cell metaplasia|8572/3
C0334395|T191|PT|68358000|SNOMEDCT_US|Adenocarcinoma with spindle cell metaplasia|8572/3
C4518223|T191|PT|733875004|SNOMEDCT_US|Fibromatosis-like metaplastic carcinoma|8572/3
C0334396|T191|PT|271470|MEDCIN|adenocarcinoma with apocrine metaplasia|8573/3
C0334396|T191|PT|C4202|NCI|Adenocarcinoma with Apocrine Metaplasia|8573/3
C0334396|T191|AB|BBB5.|RCD|Adenoca + apocrine metaplasia|8573/3
C0334396|T191|PT|BBB5.|RCD|Adenocarcinoma with apocrine metaplasia|8573/3
C0334396|T191|SY|BBB5.|RCD|Carcinoma with apocrine metaplasia|8573/3
C0334396|T191|AB|BBB5.|RCD|Carcinoma+apocrine metaplasia|8573/3
C0334396|T191|PT|22694002|SNOMEDCT_US|Adenocarcinoma with apocrine metaplasia|8573/3
C0334396|T191|SY|22694002|SNOMEDCT_US|Carcinoma with apocrine metaplasia|8573/3
C1266088|T191|PT|271471|MEDCIN|adenocarcinoma with neuroendocrine differentiation|8574/3
C1266088|T191|PT|C66745|NCI|Adenocarcinoma with Neuroendocrine Differentiation|8574/3
C1266088|T191|PT|128704005|SNOMEDCT_US|Adenocarcinoma with neuroendocrine differentiation|8574/3
C1266088|T191|SY|128704005|SNOMEDCT_US|Carcinoma with neuroendocrine differentiation|8574/3
C1266089|T191|PT|0000056682|CHV|metaplastic carcinoma|8575/3
C1266089|T191|PT|C27949|NCI|Metaplastic Carcinoma|8575/3
C1266089|T191|SY|TCGA|NCI|Metaplastic Carcinoma|8575/3
C1266089|T191|PT|C27949|NCI_CPTAC|Metaplastic Carcinoma|8575/3
C1266089|T191|PT|CDR0000044243|NCI_NCI-GLOSS|metaplastic carcinoma|8575/3
C1266089|T191|PT|128705006|SNOMEDCT_US|Metaplastic carcinoma|8575/3
C1266090|T191|LA|LA26097-8|LNC|Hepatoid adenocarcinoma|8576/3
C1266090|T191|PT|C66950|NCI|Hepatoid Adenocarcinoma|8576/3
C1266090|T191|SY|C66950|NCI|Hepatoid Carcinoma|8576/3
C1266090|T191|PT|128706007|SNOMEDCT_US|Hepatoid adenocarcinoma|8576/3
C1266090|T191|SY|128706007|SNOMEDCT_US|Hepatoid carcinoma|8576/3
C0040101|T191|PT|0007269|CCPSS|THYMOMA BENIGN|8580/0
C0040101|T191|PT|0000012247|CHV|benign thymoma|8580/0
C0040101|T191|SY|0000012247|CHV|thymoma benign|8580/0
C0040101|T191|PN|U000312|MTH|Benign Thymoma|8580/0
C0040101|T191|PT|C66746|NCI|Benign Thymoma|8580/0
C0040101|T191|OP|C66746|NCI|Benign Thymoma|8580/0
C0040101|T191|PT|BBB60|RCD|Benign thymoma|8580/0
C0040101|T191|PT|784307009|SNOMEDCT_US|Benign thymoma|8580/0
C0040101|T191|SY|21181001|SNOMEDCT_US|Benign thymoma|8580/0
C0040101|T191|OAP|134159004|SNOMEDCT_US|Benign thymoma|8580/0
C0040101|T191|PT|21181001|SNOMEDCT_US|Thymoma, benign|8580/0
C0040101|T191|IS|21181001|SNOMEDCT_US|Thymoma, NOS|8580/0
C0040100|T191|PT|0000012246|CHV|thymoma|8580/1
C0040100|T191|SY|0000012246|CHV|thymomas|8580/1
C0040100|T191|DI|U001857|DXP|THYMOMA|8580/1
C0040100|T191|PT|HP:0100522|HPO|Thymoma|8580/1
C0040100|T191|PT|MTHU074105|ICPC2ICD10ENG|thymoma|8580/1
C0040100|T191|PT|10043670|MDR|Thymoma|8580/1
C0040100|T191|LLT|10043670|MDR|Thymoma|8580/1
C0040100|T191|LLT|10043675|MDR|Thymoma NOS|8580/1
C0040100|T191|SY|1245|MEDLINEPLUS|Thymoma|8580/1
C0040100|T191|MH|D013945|MSH|Thymoma|8580/1
C0040100|T191|PM|D013945|MSH|Thymomas|8580/1
C0040100|T191|PN|NOCODE|MTH|Thymoma|8580/1
C1709024|T191|SY|C45706|NCI|Micronodular Thymoma|8580/1
C1709024|T191|SY|C45706|NCI|Micronodular Thymoma with Lymphoid B-Cell Hyperplasia|8580/1
C1709024|T191|PT|C45706|NCI|Micronodular Thymoma with Lymphoid Stroma|8580/1
C0040100|T191|PT|C3411|NCI|Thymoma|8580/1
C0040100|T191|PT|C3411|NCI_CPTAC|Thymoma|8580/1
C0040100|T191|PT|10043673|NCI_CTEP-SDC|Thymoma|8580/1
C0040100|T191|DN|C3411|NCI_CTRP|Thymoma|8580/1
C0040100|T191|PT|C3411|NCI_CTRP|Thymoma|8580/1
C0040100|T191|PT|CDR0000046002|NCI_NCI-GLOSS|thymoma|8580/1
C0040100|T191|PT|BBB6.|RCD|Thymoma|8580/1
C0040100|T191|OP|BBB6z|RCDSY|Thymoma NOS|8580/1
C1709024|T191|PT|726423000|SNOMEDCT_US|Micronodular thymoma with lymphoid stroma|8580/1
C0040100|T191|PT|444231005|SNOMEDCT_US|Thymoma|8580/1
C0040100|T191|PT|128856005|SNOMEDCT_US|Thymoma|8580/1
C0040100|T191|SY|128856005|SNOMEDCT_US|Thymoma, no ICD-O subtype|8580/1
C0040100|T191|SY|128856005|SNOMEDCT_US|Thymoma, no International Classification of Diseases for Oncology subtype|8580/1
C1322286|T191|PT|0025239|CCPSS|THYMOMA MALIGNANT|8580/3
C1322286|T191|SY|0000020761|CHV|malignant thymoma|8580/3
C1322286|T191|PT|MTHU047313|ICPC2ICD10ENG|malignant; thymoma|8580/3
C1322286|T191|PT|MTHU074106|ICPC2ICD10ENG|thymoma; malignant|8580/3
C1322286|T191|LLT|10061031|MDR|Thymoma malignant|8580/3
C1322286|T191|PT|10061031|MDR|Thymoma malignant|8580/3
C1322286|T191|LLT|10043673|MDR|Thymoma malignant NOS|8580/3
C1322286|T191|SY|230402|MEDCIN|malignant thymoma|8580/3
C1322286|T191|PT|230402|MEDCIN|malignant thymoma of thymus|8580/3
C1322286|T191|PN|NOCODE|MTH|Malignant Thymoma|8580/3
C1710027|T191|SY|C45709|NCI|Ancient Thymoma|8580/3
C1708993|T191|SY|C45707|NCI|Biphasic Thymoma|8580/3
C1708557|T191|PT|C45638|NCI|Intrapulmonary Thymoma|8580/3
C1708993|T191|SY|C45707|NCI|Low Grade Thymic Metaplastic Carcinoma|8580/3
C1322286|T191|PT|C7612|NCI|Malignant Thymoma|8580/3
C1708993|T191|PT|C45707|NCI|Metaplastic Thymoma|8580/3
C1708993|T191|SY|C45707|NCI|Mixed Polygonal and Spindle Cell Type Thymoma|8580/3
C1710027|T191|PT|C45709|NCI|Sclerosing Thymoma|8580/3
C1708993|T191|SY|C45707|NCI|Thymoma with Pseudosarcomatous Stroma|8580/3
C1322286|T191|PT|C7612|NCI_CDISC|THYMOMA, MALIGNANT|8580/3
C1322286|T191|DN|C7612|NCI_CTRP|Malignant Thymoma|8580/3
C1708557|T191|PT|734038002|SNOMEDCT_US|Intrapulmonary thymoma|8580/3
C1322286|T191|PT|444596001|SNOMEDCT_US|Malignant thymoma|8580/3
C1322286|T191|SY|15949004|SNOMEDCT_US|Malignant thymoma|8580/3
C1708993|T191|PT|726421003|SNOMEDCT_US|Metaplastic thymoma|8580/3
C1710027|T191|PT|733075000|SNOMEDCT_US|Sclerosing thymoma|8580/3
C1322286|T191|IS|15949004|SNOMEDCT_US|Thymic carcinoma|8580/3
C1322286|T191|PT|15949004|SNOMEDCT_US|Thymoma, malignant|8580/3
C1266091|T191|SY|C6454|NCI|Medullary Thymoma|8581/1
C1266091|T191|SY|C6454|NCI|Spindle Cell Thymoma|8581/1
C1266091|T191|PT|C6454|NCI|Thymoma Type A|8581/1
C1266091|T191|DN|C6454|NCI_CTRP|Thymoma Type A|8581/1
C1266091|T191|SY|CDR0000040002|PDQ|medullary thymoma|8581/1
C1266091|T191|SY|CDR0000040002|PDQ|spindle cell thymoma|8581/1
C1266091|T191|SY|CDR0000040002|PDQ|Thymoma Type A|8581/1
C1266091|T191|PT|CDR0000040002|PDQ|type A thymoma|8581/1
C1266091|T191|SY|128707003|SNOMEDCT_US|Thymoma, medullary|8581/1
C1266091|T191|SY|128707003|SNOMEDCT_US|Thymoma, spindle cell|8581/1
C1266091|T191|PT|128707003|SNOMEDCT_US|Thymoma, type A|8581/1
C0279707|T191|LLT|10041607|MDR|Spindle cell malignant thymoma|8581/3
C0279707|T191|PT|230403|MEDCIN|malignant type A thymoma|8581/3
C0279707|T191|PT|C7999|NCI|Malignant Type A Thymoma|8581/3
C0279707|T191|DN|C7999|NCI_CTRP|Malignant Type A Thymoma|8581/3
C0279707|T191|SY|128708008|SNOMEDCT_US|Thymoma, medullary, malignant|8581/3
C0279707|T191|SY|128708008|SNOMEDCT_US|Thymoma, spindle cell, malignant|8581/3
C0279707|T191|PT|128708008|SNOMEDCT_US|Thymoma, type A, malignant|8581/3
C1266092|T191|SY|C6885|NCI|Mixed Type Thymoma|8582/1
C1266092|T191|PT|C6885|NCI|Thymoma Type AB|8582/1
C1266092|T191|DN|C6885|NCI_CTRP|Thymoma Type AB|8582/1
C1266092|T191|SY|CDR0000331488|PDQ|mixed thymoma|8582/1
C1266092|T191|SY|CDR0000331488|PDQ|Mixed Type Thymoma|8582/1
C1266092|T191|SY|CDR0000331488|PDQ|Thymoma Type AB|8582/1
C1266092|T191|PT|CDR0000331488|PDQ|type AB thymoma|8582/1
C1266092|T191|SY|128709000|SNOMEDCT_US|Thymoma, mixed type|8582/1
C1266092|T191|PT|128709000|SNOMEDCT_US|Thymoma, type AB|8582/1
C1266093|T191|PT|230404|MEDCIN|malignant type AB thymoma|8582/3
C1266093|T191|PT|C6886|NCI|Malignant Type AB Thymoma|8582/3
C1266093|T191|DN|C6886|NCI_CTRP|Malignant Type AB Thymoma|8582/3
C1266093|T191|SY|128710005|SNOMEDCT_US|Thymoma, mixed type, malignant|8582/3
C1266093|T191|PT|128710005|SNOMEDCT_US|Thymoma, type AB, malignant|8582/3
C1266094|T191|PT|0000056683|CHV|lymphocytic thymoma|8583/1
C1266094|T191|SY|0000056683|CHV|type b1 thymoma|8583/1
C1266094|T191|SY|C6887|NCI|Lymphocyte-Predominant Thymoma|8583/1
C1266094|T191|SY|C6887|NCI|Lymphocyte-Rich Thymoma|8583/1
C1266094|T191|SY|C6887|NCI|Organoid Thymoma|8583/1
C1266094|T191|SY|C6887|NCI|Predominantly Cortical Thymoma|8583/1
C1266094|T191|PT|C6887|NCI|Thymoma Type B1|8583/1
C1266094|T191|DN|C6887|NCI_CTRP|Thymoma Type B1|8583/1
C1266094|T191|SY|CDR0000039999|PDQ|Lymphocyte-Predominant Thymoma|8583/1
C1266094|T191|SY|CDR0000039999|PDQ|lymphocyte-rich thymoma|8583/1
C1266094|T191|SY|CDR0000039999|PDQ|lymphocytic thymoma|8583/1
C1266094|T191|SY|CDR0000039999|PDQ|organoid thymoma|8583/1
C1266094|T191|SY|CDR0000039999|PDQ|predominantly cortical thymoma|8583/1
C1266094|T191|SY|CDR0000039999|PDQ|Thymoma Type B1|8583/1
C1266094|T191|PT|CDR0000039999|PDQ|type B1 thymoma|8583/1
C1266094|T191|SY|128711009|SNOMEDCT_US|Thymoma, lymphocyte-rich|8583/1
C1266094|T191|SY|128711009|SNOMEDCT_US|Thymoma, lymphocytic|8583/1
C1266094|T191|SY|128711009|SNOMEDCT_US|Thymoma, organoid|8583/1
C1266094|T191|SY|128711009|SNOMEDCT_US|Thymoma, predominantly cortical|8583/1
C1266094|T191|PT|128711009|SNOMEDCT_US|Thymoma, type B1|8583/1
C0279704|T191|LLT|10025272|MDR|Lymphocytic malignant thymoma|8583/3
C0279704|T191|PT|230405|MEDCIN|malignant type B1 thymoma|8583/3
C0279704|T191|PT|C7996|NCI|Malignant Type B1 Thymoma|8583/3
C0279704|T191|DN|C7996|NCI_CTRP|Malignant Type B1 Thymoma|8583/3
C0279704|T191|SY|128712002|SNOMEDCT_US|Thymoma, lymphocyte-rich, malignant|8583/3
C0279704|T191|SY|128712002|SNOMEDCT_US|Thymoma, lymphocytic, malignant|8583/3
C0279704|T191|SY|128712002|SNOMEDCT_US|Thymoma, organoid, malignant|8583/3
C0279704|T191|SY|128712002|SNOMEDCT_US|Thymoma, predominantly cortical, malignant|8583/3
C0279704|T191|PT|128712002|SNOMEDCT_US|Thymoma, type B1, malignant|8583/3
C1266095|T191|SY|C6888|NCI|Cortical Thymoma|8584/1
C1266095|T191|SY|C6888|NCI|Polygonal Cell Thymoma|8584/1
C1266095|T191|PT|C6888|NCI|Thymoma Type B2|8584/1
C1266095|T191|DN|C6888|NCI_CTRP|Thymoma Type B2|8584/1
C1266095|T191|SY|CDR0000331683|PDQ|cortical thymoma|8584/1
C1266095|T191|SY|CDR0000331683|PDQ|polygonal cell thymoma|8584/1
C1266095|T191|SY|CDR0000331683|PDQ|Thymoma Type B2|8584/1
C1266095|T191|PT|CDR0000331683|PDQ|type B2 thymoma|8584/1
C1266095|T191|SY|128713007|SNOMEDCT_US|Thymoma, cortical|8584/1
C1266095|T191|PT|128713007|SNOMEDCT_US|Thymoma, type B2|8584/1
C1266096|T191|PT|230406|MEDCIN|malignant type B2 thymoma|8584/3
C1266096|T191|PT|C6889|NCI|Malignant Type B2 Thymoma|8584/3
C1266096|T191|DN|C6889|NCI_CTRP|Malignant Type B2 Thymoma|8584/3
C1266096|T191|SY|128714001|SNOMEDCT_US|Thymoma, cortical, malignant|8584/3
C1266096|T191|PT|128714001|SNOMEDCT_US|Thymoma, type B2, malignant|8584/3
C0279705|T191|LLT|10015094|MDR|Epithelial malignant thymoma|8585/1
C0279705|T191|PT|230407|MEDCIN|malignant type B3 thymoma|8585/1
C0279705|T191|SY|C7997|NCI|Atypical Thymoma|8585/1
C0279705|T191|SY|C7997|NCI|Epithelial Malignant Thymoma|8585/1
C0279705|T191|SY|C7997|NCI|Epithelial Thymoma|8585/1
C0279705|T191|SY|C7997|NCI|Malignant Thymoma Type B3|8585/1
C0279705|T191|SY|C7997|NCI|Squamoid Thymoma|8585/1
C0279705|T191|PT|C7997|NCI|Thymoma Type B3|8585/1
C0279705|T191|SY|C7997|NCI|Well Differentiated Thymic Carcinoma|8585/1
C0279705|T191|SY|C7997|NCI|Well-Differentiated Thymic Carcinoma|8585/1
C0279705|T191|DN|C7997|NCI_CTRP|Thymoma Type B3|8585/1
C0279705|T191|SY|CDR0000040000|PDQ|atypical thymoma|8585/1
C0279705|T191|SY|CDR0000040000|PDQ|Epithelial Malignant Thymoma|8585/1
C0279705|T191|SY|CDR0000040000|PDQ|epithelial thymoma|8585/1
C0279705|T191|SY|CDR0000040000|PDQ|Malignant Thymoma Type B3|8585/1
C0279705|T191|SY|CDR0000040000|PDQ|squamoid thymoma|8585/1
C0279705|T191|SY|CDR0000040000|PDQ|Thymoma Type B3|8585/1
C0279705|T191|PT|CDR0000040000|PDQ|type B3 thymoma|8585/1
C0279705|T191|SY|CDR0000040000|PDQ|Well Differentiated Thymic Carcinoma|8585/1
C0279705|T191|SY|CDR0000040000|PDQ|well-differentiated thymic carcinoma|8585/1
C0279705|T191|SY|128715000|SNOMEDCT_US|Thymoma, atypical|8585/1
C0279705|T191|SY|128716004|SNOMEDCT_US|Thymoma, atypical, malignant|8585/1
C0279705|T191|SY|128715000|SNOMEDCT_US|Thymoma, epithelial|8585/1
C0279705|T191|SY|128716004|SNOMEDCT_US|Thymoma, epithelial, malignant|8585/1
C0279705|T191|PT|128715000|SNOMEDCT_US|Thymoma, type B3|8585/1
C0279705|T191|PT|128716004|SNOMEDCT_US|Thymoma, type B3, malignant|8585/1
C0279705|T191|SY|128716004|SNOMEDCT_US|Well differentiated thymic carcinoma|8585/1
C0279705|T191|LLT|10015094|MDR|Epithelial malignant thymoma|8585/3
C0279705|T191|PT|230407|MEDCIN|malignant type B3 thymoma|8585/3
C0279705|T191|SY|C7997|NCI|Atypical Thymoma|8585/3
C0279705|T191|SY|C7997|NCI|Epithelial Malignant Thymoma|8585/3
C0279705|T191|SY|C7997|NCI|Epithelial Thymoma|8585/3
C0279705|T191|SY|C7997|NCI|Malignant Thymoma Type B3|8585/3
C0279705|T191|SY|C7997|NCI|Squamoid Thymoma|8585/3
C0279705|T191|PT|C7997|NCI|Thymoma Type B3|8585/3
C0279705|T191|SY|C7997|NCI|Well Differentiated Thymic Carcinoma|8585/3
C0279705|T191|SY|C7997|NCI|Well-Differentiated Thymic Carcinoma|8585/3
C0279705|T191|DN|C7997|NCI_CTRP|Thymoma Type B3|8585/3
C0279705|T191|SY|CDR0000040000|PDQ|atypical thymoma|8585/3
C0279705|T191|SY|CDR0000040000|PDQ|Epithelial Malignant Thymoma|8585/3
C0279705|T191|SY|CDR0000040000|PDQ|epithelial thymoma|8585/3
C0279705|T191|SY|CDR0000040000|PDQ|Malignant Thymoma Type B3|8585/3
C0279705|T191|SY|CDR0000040000|PDQ|squamoid thymoma|8585/3
C0279705|T191|SY|CDR0000040000|PDQ|Thymoma Type B3|8585/3
C0279705|T191|PT|CDR0000040000|PDQ|type B3 thymoma|8585/3
C0279705|T191|SY|CDR0000040000|PDQ|Well Differentiated Thymic Carcinoma|8585/3
C0279705|T191|SY|CDR0000040000|PDQ|well-differentiated thymic carcinoma|8585/3
C0279705|T191|SY|128715000|SNOMEDCT_US|Thymoma, atypical|8585/3
C0279705|T191|SY|128716004|SNOMEDCT_US|Thymoma, atypical, malignant|8585/3
C0279705|T191|SY|128715000|SNOMEDCT_US|Thymoma, epithelial|8585/3
C0279705|T191|SY|128716004|SNOMEDCT_US|Thymoma, epithelial, malignant|8585/3
C0279705|T191|PT|128715000|SNOMEDCT_US|Thymoma, type B3|8585/3
C0279705|T191|PT|128716004|SNOMEDCT_US|Thymoma, type B3, malignant|8585/3
C0279705|T191|SY|128716004|SNOMEDCT_US|Well differentiated thymic carcinoma|8585/3
C0205969|T191|PT|0000020761|CHV|thymic carcinoma|8586/3
C0205969|T191|SY|0000020761|CHV|thymic carcinomas|8586/3
C0205969|T191|PT|MTHU014826|ICPC2ICD10ENG|carcinoma; thymic|8586/3
C0205969|T191|PT|MTHU074116|ICPC2ICD10ENG|thymic; carcinoma|8586/3
C0205969|T191|PEP|D013945|MSH|Carcinoma, Thymic|8586/3
C0205969|T191|PM|D013945|MSH|Carcinomas, Thymic|8586/3
C0205969|T191|PM|D013945|MSH|Thymic Carcinoma|8586/3
C0205969|T191|PM|D013945|MSH|Thymic Carcinomas|8586/3
C0205969|T191|PN|NOCODE|MTH|Thymic Carcinoma|8586/3
C0205969|T191|PT|C7569|NCI|Thymic Carcinoma|8586/3
C0205969|T191|SY|C7569|NCI|Thymic Carcinoma Excluding Well Differentiated Thymic Carcinoma|8586/3
C0205969|T191|OP|C7569|NCI|Thymoma Type C|8586/3
C0205969|T191|PT|C7569|NCI_CPTAC|Thymic Carcinoma|8586/3
C0205969|T191|PT|C7569|NCI_CTRP|Thymic Carcinoma|8586/3
C0205969|T191|DN|C7569|NCI_CTRP|Thymic Carcinoma|8586/3
C0205969|T191|PT|CDR0000455462|NCI_NCI-GLOSS|thymic carcinoma|8586/3
C0205969|T191|PT|CDR0000467224|NCI_NCI-GLOSS|type C thymoma|8586/3
C0205969|T191|ET|CDR0000331691|PDQ|thymic carcinoma|8586/3
C0205969|T191|PT|CDR0000331691|PDQ|thymic carcinoma|8586/3
C0205969|T191|SY|CDR0000331691|PDQ|Thymic Carcinoma Excluding Well Differentiated Thymic Carcinoma|8586/3
C0205969|T191|ET|CDR0000038797|PDQ|Thymoma and thymic carcinoma|8586/3
C0205969|T191|PSC|CDR0000038797|PDQ|thymoma and thymic carcinoma|8586/3
C0205969|T191|IS|CDR0000331691|PDQ|Thymoma Type C|8586/3
C0205969|T191|SY|CDR0000331691|PDQ|type C thymoma|8586/3
C0205969|T191|PT|BBB61|RCD|Malignant thymoma|8586/3
C0205969|T191|SY|BBB61|RCD|Thymic carcinoma|8586/3
C0205969|T191|SY|128717008|SNOMEDCT_US|Thymic carcinoma|8586/3
C0205969|T191|PT|128717008|SNOMEDCT_US|Thymoma, type C|8586/3
C0205969|T191|PT|444374006|SNOMEDCT_US|Type C thymoma|8586/3
C1266098|T191|SY|C53595|NCI|Branchial Anlage Mixed Tumor|8587/0
C1266098|T191|PT|C53595|NCI|Ectopic Hamartomatous Thymoma|8587/0
C1266098|T191|PT|128718003|SNOMEDCT_US|Ectopic hamartomatous thymoma|8587/0
C1266099|T191|PT|0000056684|CHV|settle|8588/3
C1266099|T191|SY|0000056684|CHV|settles|8588/3
C1266099|T191|PT|230409|MEDCIN|spindle epithelial tumor with thymus-like element|8588/3
C1266099|T191|PN|NOCODE|MTH|Thyroid Gland Spindle Cell Tumor with Thymus-Like Differentiation|8588/3
C1266099|T191|AB|C46105|NCI|SETTLE|8588/3
C1266099|T191|PT|C46105|NCI|Thyroid Gland Spindle Cell Tumor with Thymus-Like Differentiation|8588/3
C1266099|T191|SY|128719006|SNOMEDCT_US|SETTLE|8588/3
C1266099|T191|SY|128719006|SNOMEDCT_US|Spindle epithelial tumor with thymus-like differentiation|8588/3
C1266099|T191|PT|128719006|SNOMEDCT_US|Spindle epithelial tumor with thymus-like element|8588/3
C1266099|T191|SYGB|128719006|SNOMEDCT_US|Spindle epithelial tumour with thymus-like differentiation|8588/3
C1266099|T191|PTGB|128719006|SNOMEDCT_US|Spindle epithelial tumour with thymus-like element|8588/3
C1266100|T191|PT|0000056685|CHV|carcinoma showing thymus-like element|8589/3
C1266100|T191|SY|0000056685|CHV|castle|8589/3
C1266100|T191|SY|0000056685|CHV|castles|8589/3
C1266100|T191|PT|230410|MEDCIN|carcinoma showing thymus-like element|8589/3
C1266100|T191|PN|NOCODE|MTH|Carcinoma showing thymus-like element|8589/3
C1704613|T191|PN|NOCODE|MTH|Thyroid Gland Carcinoma Showing Thymus-Like Differentiation|8589/3
C1704613|T191|AB|C46106|NCI|CASTLE|8589/3
C1704613|T191|PT|C46106|NCI|Intrathyroid Thymic Carcinoma|8589/3
C1704613|T191|SY|C46106|NCI|Thyroid Gland Carcinoma Showing Thymus-Like Differentiation|8589/3
C1266100|T191|SY|128720000|SNOMEDCT_US|Carcinoma showing thymus-like differentiation|8589/3
C1266100|T191|PT|128720000|SNOMEDCT_US|Carcinoma showing thymus-like element|8589/3
C1266100|T191|SY|128720000|SNOMEDCT_US|CASTLE|8589/3
C3838965|T191|PT|703599008|SNOMEDCT_US|Microcystic stromal tumor|8590/0
C3838965|T191|PTGB|703599008|SNOMEDCT_US|Microcystic stromal tumour|8590/0
C3839428|T191|PT|703597005|SNOMEDCT_US|Sex cord-stromal tumor, benign|8590/0
C3839428|T191|PTGB|703597005|SNOMEDCT_US|Sex cord-stromal tumour, benign|8590/0
C3839205|T191|PT|703598000|SNOMEDCT_US|Signet-ring stromal tumor|8590/0
C3839205|T191|PTGB|703598000|SNOMEDCT_US|Signet-ring stromal tumour|8590/0
C0206724|T191|SY|0000021048|CHV|cord sex stromal tumors|8590/1
C0206724|T191|SY|0000021048|CHV|cord sex tumors|8590/1
C0206724|T191|SY|0000021048|CHV|gonadal stromal tumor|8590/1
C0206724|T191|PT|0000021048|CHV|sex cord stromal tumor|8590/1
C0206724|T191|SY|0000021048|CHV|sex cord tumor|8590/1
C0206724|T191|PM|D018312|MSH|Sex Cord Stromal Tumor|8590/1
C0206724|T191|MH|D018312|MSH|Sex Cord-Gonadal Stromal Tumors|8590/1
C0206724|T191|ET|D018312|MSH|Sex Cord-Stromal Tumor|8590/1
C0206724|T191|PM|D018312|MSH|Sex Cord-Stromal Tumors|8590/1
C0206724|T191|PM|D018312|MSH|Tumor, Sex Cord-Stromal|8590/1
C0206724|T191|PM|D018312|MSH|Tumors, Sex Cord-Stromal|8590/1
C0206724|T191|PN|NOCODE|MTH|Sex Cord-Stromal Tumor|8590/1
C0206724|T191|SY|C3794|NCI|Sex Cord-Stromal Neoplasm|8590/1
C0206724|T191|PT|C3794|NCI|Sex Cord-Stromal Tumor|8590/1
C0206724|T191|PT|CDR0000642163|NCI_NCI-GLOSS|sex cord tumor|8590/1
C0206724|T191|PT|CDR0000642165|NCI_NCI-GLOSS|sex cord-gonadal stromal tumor|8590/1
C0206724|T191|PT|CDR0000642164|NCI_NCI-GLOSS|sex cord-stromal tumor|8590/1
C0206724|T191|PT|C3794|NCI_NICHD|Sex Cord-Stromal Tumor|8590/1
C0206724|T191|IS|X77o4|RCD|Gonadal stromal tumour|8590/1
C0206724|T191|IS|X77o4|RCD|Sex cord stromal tumour|8590/1
C0206724|T191|IS|X77o4|RCD|Sex cord tumour|8590/1
C0206724|T191|PT|Xa99B|RCD|Specialised gonadal tumour|8590/1
C0206724|T191|IS|X77o4|RCDAE|Gonadal stromal tumor|8590/1
C0206724|T191|IS|X77o4|RCDAE|Sex cord stromal tumor|8590/1
C0206724|T191|IS|X77o4|RCDAE|Sex cord tumor|8590/1
C0206724|T191|PT|Xa99B|RCDAE|Specialized gonadal tumor|8590/1
C0206724|T191|OA|BBC..|RCDSA|Specialized gonadal neopl.|8590/1
C0206724|T191|OP|BBCz.|RCDSA|Specialized gonadal neoplasm NOS|8590/1
C0206724|T191|OP|BBC..|RCDSA|Specialized gonadal neoplasms|8590/1
C0206724|T191|OA|BBCz.|RCDSY|Special gonadal neopl.NOS|8590/1
C0206724|T191|OA|BBC..|RCDSY|Specialised gonadal neopl.|8590/1
C0206724|T191|OP|BBCz.|RCDSY|Specialised gonadal neoplasm NOS|8590/1
C0206724|T191|OP|BBC..|RCDSY|Specialised gonadal neoplasms|8590/1
C0206724|T191|SY|71440001|SNOMEDCT_US|Gonadal stromal tumor|8590/1
C0206724|T191|SYGB|71440001|SNOMEDCT_US|Gonadal stromal tumour|8590/1
C0206724|T191|OAS|253028001|SNOMEDCT_US|Sex cord stromal tumor|8590/1
C0206724|T191|OAS|253028001|SNOMEDCT_US|Sex cord stromal tumour|8590/1
C0206724|T191|SY|71440001|SNOMEDCT_US|Sex cord tumor|8590/1
C0206724|T191|IS|71440001|SNOMEDCT_US|Sex cord tumor, NOS|8590/1
C0206724|T191|SYGB|71440001|SNOMEDCT_US|Sex cord tumour|8590/1
C0206724|T191|PT|71440001|SNOMEDCT_US|Sex cord-stromal tumor|8590/1
C0206724|T191|SY|71440001|SNOMEDCT_US|Sex cord-stromal tumor, no ICD-O subtype|8590/1
C0206724|T191|SY|71440001|SNOMEDCT_US|Sex cord-stromal tumor, no International Classification of Diseases for Oncology subtype|8590/1
C0206724|T191|PTGB|71440001|SNOMEDCT_US|Sex cord-stromal tumour|8590/1
C0206724|T191|SYGB|71440001|SNOMEDCT_US|Sex cord-stromal tumour, no ICD-O subtype|8590/1
C0206724|T191|PTGB|115221000|SNOMEDCT_US|Specialised gonadal neoplasm|8590/1
C0206724|T191|OAP|134323003|SNOMEDCT_US|Specialised gonadal tumour|8590/1
C0206724|T191|PT|115221000|SNOMEDCT_US|Specialized gonadal neoplasm|8590/1
C0206724|T191|OAP|134323003|SNOMEDCT_US|Specialized gonadal tumor|8590/1
C3839747|T191|PT|703600006|SNOMEDCT_US|Uterine tumor resembling ovarian sex cord tumor|8590/1
C3839747|T191|PTGB|703600006|SNOMEDCT_US|Uterine tumour resembling ovarian sex cord tumour|8590/1
C1848186|T191|PT|C67561|NCI|Malignant Sex Cord-Stromal Tumor|8590/3
C1848186|T191|SY|C67561|NCI_CDISC|Sex Cord Stromal Tumor, Malignant|8590/3
C1848186|T191|PT|C67561|NCI_CDISC|STROMAL TUMOR, GONADAL, MALIGNANT|8590/3
C1266102|T191|PN|NOCODE|MTH|Testicular Sex Cord-Gonadal Stromal Tumor, Incompletely Differentiated|8591/1
C1266102|T191|SY|C66748|NCI|Sex Cord-Gonadal Stromal Tumor, Incompletely Differentiated|8591/1
C1266102|T191|SY|C66748|NCI|Testicular Sex Cord-Gonadal Stromal Tumor with Indeterminate Differentiation|8591/1
C1266102|T191|SY|C66748|NCI|Testicular Sex Cord-Gonadal Stromal Tumor, Incompletely Differentiated|8591/1
C1266102|T191|SY|C66748|NCI|Unclassified Testicular Sex Cord-Gonadal Stromal Tumor|8591/1
C1266102|T191|PT|C66748|NCI|Unclassified Testicular Sex Cord-Stromal Tumor|8591/1
C1266102|T191|PT|128721001|SNOMEDCT_US|Sex cord-gonadal stromal tumor, incompletely differentiated|8591/1
C1266102|T191|PTGB|128721001|SNOMEDCT_US|Sex cord-gonadal stromal tumour, incompletely differentiated|8591/1
C1266103|T191|PN|NOCODE|MTH|Testicular Sex Cord-Gonadal Stromal Tumor, Mixed Forms|8592/1
C1321220|T191|SY|C5241|NCI|Mixed Germ Cell-Sex Cord Neoplasm|8592/1
C1321220|T191|SY|C5241|NCI|Mixed Germ Cell-Sex Cord Tumor|8592/1
C1321220|T191|SY|C5241|NCI|Mixed Germ Cell-Sex Cord-Stromal Neoplasm|8592/1
C1321220|T191|PT|C5241|NCI|Mixed Germ Cell-Sex Cord-Stromal Tumor|8592/1
C1266103|T191|SY|C66991|NCI|Mixed Testicular Sex Cord-Gonadal Stromal Tumor|8592/1
C1266103|T191|PT|C66991|NCI|Mixed Testicular Sex Cord-Stromal Tumor|8592/1
C1266103|T191|SY|C66991|NCI|Sex Cord-Gonadal Stromal Tumor, Mixed Forms|8592/1
C1266103|T191|SY|C66991|NCI|Testicular Sex Cord-Gonadal Stromal Tumor, Mixed Forms|8592/1
C1321220|T191|PT|C5241|NCI_NICHD|Mixed Germ Cell-Sex Cord-Stromal Tumor|8592/1
C1321220|T191|OP|703601005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumor|8592/1
C1321220|T191|PT|406096006|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumor|8592/1
C1321220|T191|PT|703601005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumor, no International Classification of Diseases for Oncology subtype|8592/1
C1321220|T191|OP|703601005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumour|8592/1
C1321220|T191|PTGB|406096006|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumour|8592/1
C1321220|T191|PTGB|703601005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumour, no International Classification of Diseases for Oncology subtype|8592/1
C1266103|T191|PT|128722008|SNOMEDCT_US|Sex cord-gonadal stromal tumor, mixed forms|8592/1
C1266103|T191|PTGB|128722008|SNOMEDCT_US|Sex cord-gonadal stromal tumour, mixed forms|8592/1
C1883177|T191|PN|NOCODE|MTH|Ovarian Stromal Tumor with Minor Sex Cord Elements|8593/1
C1266104|T191|PN|NOCODE|MTH|Stromal tumor with minor sex cord elements|8593/1
C1883177|T191|PT|C66749|NCI|Ovarian Stromal Tumor with Minor Sex Cord Elements|8593/1
C1883177|T191|SY|C66749|NCI|Stromal Tumor with Minor Sex Cord Elements|8593/1
C1266104|T191|PT|128723003|SNOMEDCT_US|Stromal tumor with minor sex cord elements|8593/1
C1266104|T191|PTGB|128723003|SNOMEDCT_US|Stromal tumour with minor sex cord elements|8593/1
C1321220|T191|SY|C5241|NCI|Mixed Germ Cell-Sex Cord Neoplasm|8594/1
C1321220|T191|SY|C5241|NCI|Mixed Germ Cell-Sex Cord Tumor|8594/1
C1321220|T191|SY|C5241|NCI|Mixed Germ Cell-Sex Cord-Stromal Neoplasm|8594/1
C1321220|T191|PT|C5241|NCI|Mixed Germ Cell-Sex Cord-Stromal Tumor|8594/1
C1321220|T191|PT|C5241|NCI_NICHD|Mixed Germ Cell-Sex Cord-Stromal Tumor|8594/1
C1321220|T191|OP|703601005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumor|8594/1
C1321220|T191|PT|406096006|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumor|8594/1
C1321220|T191|PT|703601005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumor, no International Classification of Diseases for Oncology subtype|8594/1
C3839834|T191|PT|703602003|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumor, unclassified|8594/1
C1321220|T191|OP|703601005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumour|8594/1
C1321220|T191|PTGB|406096006|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumour|8594/1
C1321220|T191|PTGB|703601005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumour, no International Classification of Diseases for Oncology subtype|8594/1
C3839834|T191|PTGB|703602003|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumour, unclassified|8594/1
C0039747|T191|SY|0000012152|CHV|theca cell tumor|8600/0
C0039747|T191|PT|0000012152|CHV|thecoma|8600/0
C0039747|T191|SY|0000012152|CHV|thecomas|8600/0
C0039747|T191|SY|NOCODE|DXP|THECOMA|8600/0
C0039747|T191|PT|MTHU073984|ICPC2ICD10ENG|theca cell; tumor|8600/0
C0039747|T191|PT|MTHU073986|ICPC2ICD10ENG|thecoma|8600/0
C0039747|T191|PT|MTHU077162|ICPC2ICD10ENG|tumor; theca cell|8600/0
C0039747|T191|LLT|10062594|MDR|Thecoma|8600/0
C0039747|T191|PN|NOCODE|MTH|Thecoma|8600/0
C0039747|T191|PT|C3405|NCI|Thecoma|8600/0
C0039747|T191|SY|X77o6|RCD|Theca cell tumour|8600/0
C0039747|T191|PT|X77o6|RCD|Thecoma|8600/0
C0039747|T191|SY|X77o6|RCDAE|Theca cell tumor|8600/0
C0039747|T191|OP|BBC1z|RCDSY|Thecal cell neoplasm NOS|8600/0
C0039747|T191|OP|BBC1.|RCDSY|Thecal cell neoplasms|8600/0
C0039747|T191|OP|BBC10|RCDSY|Thecoma NOS|8600/0
C0039747|T191|IS|52490000|SNOMEDCT_US|Fibrothecoma|8600/0
C0039747|T191|SY|52490000|SNOMEDCT_US|Theca cell tumor|8600/0
C0039747|T191|SYGB|52490000|SNOMEDCT_US|Theca cell tumour|8600/0
C0039747|T191|PT|52490000|SNOMEDCT_US|Thecoma|8600/0
C0039747|T191|SY|52490000|SNOMEDCT_US|Thecoma, no ICD-O subtype|8600/0
C0039747|T191|SY|52490000|SNOMEDCT_US|Thecoma, no International Classification of Diseases for Oncology subtype|8600/0
C0039747|T191|IS|52490000|SNOMEDCT_US|Thecoma, NOS|8600/0
C0334398|T191|SY|NOCODE|DXP|OVARIAN CANCER, THECA CELL|8600/3
C0334398|T191|PT|MTHU047312|ICPC2ICD10ENG|malignant; thecoma|8600/3
C0334398|T191|PT|MTHU073988|ICPC2ICD10ENG|thecoma; malignant|8600/3
C0334398|T191|PT|233140|MEDCIN|malignant thecoma of ovary|8600/3
C0334398|T191|PN|NOCODE|MTH|Malignant Ovarian Thecoma|8600/3
C0334398|T191|SY|C6929|NCI|Malignant Ovarian Thecal Cell Neoplasm|8600/3
C0334398|T191|SY|C6929|NCI|Malignant Ovarian Thecal Cell Tumor|8600/3
C0334398|T191|PT|C6929|NCI|Malignant Ovarian Thecoma|8600/3
C0334398|T191|SY|C6929|NCI|Malignant Thecal Cell Neoplasm of Ovary|8600/3
C0334398|T191|SY|C6929|NCI|Malignant Thecal Cell Neoplasm of the Ovary|8600/3
C0334398|T191|SY|C6929|NCI|Malignant Thecal Cell Tumor of Ovary|8600/3
C0334398|T191|SY|C6929|NCI|Malignant Thecal Cell Tumor of the Ovary|8600/3
C0334398|T191|SY|C6929|NCI|Malignant Thecoma of Ovary|8600/3
C0334398|T191|SY|C6929|NCI|Malignant Thecoma of the Ovary|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Malignant Ovarian Thecal Cell Neoplasm|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Malignant Ovarian Thecal Cell Tumor|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Malignant Thecal Cell Neoplasm of Ovary|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Malignant Thecal Cell Neoplasm of the Ovary|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Malignant Thecal Cell Tumor of Ovary|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Malignant Thecal Cell Tumor of the Ovary|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Malignant Thecoma of Ovary|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Malignant Thecoma of the Ovary|8600/3
C0334398|T191|SY|C6929|NCI_CDISC|Thecoma, Malignant|8600/3
C0334398|T191|PT|C6929|NCI_CDISC|THECOMA, OVARIAN, MALIGNANT|8600/3
C0334398|T191|PT|X77o7|RCD|Malignant thecoma|8600/3
C0334398|T191|SY|57622002|SNOMEDCT_US|Malignant thecoma|8600/3
C0334398|T191|PT|57622002|SNOMEDCT_US|Thecoma, malignant|8600/3
C0334399|T191|PT|MTHU031190|ICPC2ICD10ENG|luteinized; thecoma|8601/0
C0334399|T191|PT|MTHU073987|ICPC2ICD10ENG|thecoma; luteinized|8601/0
C0334399|T191|SY|C4203|NCI|Luteinized Ovarian Thecoma|8601/0
C0334399|T191|SY|C4203|NCI|Luteinized Thecoma of Ovary|8601/0
C0334399|T191|SY|C4203|NCI|Luteinized Thecoma of the Ovary|8601/0
C0334399|T191|PT|C4203|NCI|Ovarian Luteinized Thecoma|8601/0
C0334399|T191|PT|X77o8|RCD|Luteinised thecoma|8601/0
C0334399|T191|PT|X77o8|RCDAE|Luteinized thecoma|8601/0
C0334399|T191|OAP|189730009|SNOMEDCT_US|Luteinised thecoma|8601/0
C0334399|T191|OF|189730009|SNOMEDCT_US|Luteinised thecoma|8601/0
C0334399|T191|OAP|189730009|SNOMEDCT_US|Luteinized thecoma|8601/0
C0334399|T191|PTGB|54482004|SNOMEDCT_US|Thecoma, luteinised|8601/0
C0334399|T191|PT|54482004|SNOMEDCT_US|Thecoma, luteinized|8601/0
C0334400|T191|PT|MTHU066710|ICPC2ICD10ENG|sclerosing; stromal tumor|8602/0
C0334400|T191|PT|MTHU077148|ICPC2ICD10ENG|tumor; sclerosing stromal|8602/0
C1368821|T191|SY|C4204|NCI|Ovarian Sclerosing Stromal Neoplasm|8602/0
C1368821|T191|PT|C4204|NCI|Ovarian Sclerosing Stromal Tumor|8602/0
C1368821|T191|SY|C4204|NCI|Sclerosing Stromal Neoplasm of Ovary|8602/0
C1368821|T191|SY|C4204|NCI|Sclerosing Stromal Neoplasm of the Ovary|8602/0
C1368821|T191|SY|C4204|NCI|Sclerosing Stromal Tumor of Ovary|8602/0
C1368821|T191|SY|C4204|NCI|Sclerosing Stromal Tumor of the Ovary|8602/0
C0334400|T191|PT|X77o5|RCD|Sclerosing stromal tumour|8602/0
C0334400|T191|PT|X77o5|RCDAE|Sclerosing stromal tumor|8602/0
C0334400|T191|OAP|189740007|SNOMEDCT_US|Sclerosing stromal tumor|8602/0
C0334400|T191|PT|64512009|SNOMEDCT_US|Sclerosing stromal tumor|8602/0
C0334400|T191|OF|189740007|SNOMEDCT_US|Sclerosing stromal tumour|8602/0
C0334400|T191|PTGB|64512009|SNOMEDCT_US|Sclerosing stromal tumour|8602/0
C0334400|T191|OAP|189740007|SNOMEDCT_US|Sclerosing stromal tumour|8602/0
C0024167|T191|SY|0000007582|CHV|luteinoma|8610/0
C0024167|T191|PT|0000007582|CHV|luteoma|8610/0
C0024167|T191|ET|2016-1387|CSP|luteoma|8610/0
C0024167|T191|PT|MTHU046318|ICPC2ICD10ENG|luteinoma|8610/0
C0024167|T191|PT|MTHU046320|ICPC2ICD10ENG|luteoma|8610/0
C0024167|T191|ET|D018311|MSH|Luteinoma|8610/0
C0024167|T191|MH|D018311|MSH|Luteoma|8610/0
C0024167|T191|PM|D018311|MSH|Luteomas|8610/0
C0024167|T191|SY|C3202|NCI|Luteal Cell Neoplasm|8610/0
C0024167|T191|SY|C3202|NCI|Luteal Cell Tumor|8610/0
C0024167|T191|SY|C3202|NCI|Luteinoma|8610/0
C0024167|T191|SY|C3202|NCI|Luteoma|8610/0
C0024167|T191|PT|C3202|NCI|Ovarian Stromal Luteoma|8610/0
C0024167|T191|SY|C3202|NCI_CDISC|Luteal Cell Neoplasm|8610/0
C0024167|T191|SY|C3202|NCI_CDISC|Luteal Cell Tumor|8610/0
C0024167|T191|SY|C3202|NCI_CDISC|Luteinoma|8610/0
C0024167|T191|SY|C3202|NCI_CDISC|Luteoma|8610/0
C0024167|T191|PT|C3202|NCI_CDISC|LUTEOMA, BENIGN|8610/0
C0024167|T191|SY|C3202|NCI_CDISC|Ovarian Stroma Luteoma|8610/0
C0024167|T191|SY|Xa99E|RCD|Luteinoma|8610/0
C0024167|T191|PT|Xa99E|RCD|Luteoma|8610/0
C0024167|T191|OP|BBC2.|RCDSY|Luteoma NOS|8610/0
C0024167|T191|SY|26372004|SNOMEDCT_US|Luteal cell tumor|8610/0
C0024167|T191|SYGB|26372004|SNOMEDCT_US|Luteal cell tumour|8610/0
C0024167|T191|SY|26372004|SNOMEDCT_US|Luteinoma|8610/0
C0024167|T191|PT|26372004|SNOMEDCT_US|Luteoma|8610/0
C0024167|T191|IS|26372004|SNOMEDCT_US|Luteoma, NOS|8610/0
C0018206|T191|SY|0000005693|CHV|cell granulosa tumor|8620/1
C0018206|T191|SY|0000005693|CHV|cells granulosa tumor|8620/1
C0018206|T191|PT|0000005693|CHV|granulosa cell tumor|8620/1
C0018206|T191|SY|0000005693|CHV|granulosa cell tumors|8620/1
C0018206|T191|SY|0000005693|CHV|granulosa cell tumour|8620/1
C0018206|T191|SY|0000005693|CHV|tumor cell granulosa|8620/1
C0018206|T191|PT|MTHU032840|ICPC2ICD10ENG|granulosa cell; tumor|8620/1
C0018206|T191|PT|MTHU077068|ICPC2ICD10ENG|tumor; granulosa cell|8620/1
C0018206|T191|MH|D006106|MSH|Granulosa Cell Tumor|8620/1
C0018206|T191|PM|D006106|MSH|Granulosa Cell Tumors|8620/1
C0018206|T191|PM|D006106|MSH|Tumor, Granulosa Cell|8620/1
C0018206|T191|PM|D006106|MSH|Tumors, Granulosa Cell|8620/1
C0018206|T191|PN|NOCODE|MTH|granulosa cell tumor|8620/1
C1879643|T191|PT|C66750|NCI|Adult Type Granulosa Cell Tumor|8620/1
C0018206|T191|SY|C3070|NCI|Granulosa Cell Neoplasm|8620/1
C0018206|T191|PT|C3070|NCI|Granulosa Cell Tumor|8620/1
C0018206|T191|PT|CDR0000044780|NCI_NCI-GLOSS|granulosa cell tumor|8620/1
C0018206|T191|PT|C3070|NCI_NICHD|Granulosa Cell Tumor|8620/1
C0018206|T191|PT|Xa99G|RCD|Granulosa cell tumour|8620/1
C0018206|T191|PT|Xa99G|RCDAE|Granulosa cell tumor|8620/1
C0018206|T191|OP|BBC3.|RCDSA|Granulosa cell tumor NOS|8620/1
C0018206|T191|OP|BBC3.|RCDSY|Granulosa cell tumour NOS|8620/1
C4542861|T191|PT|734274003|SNOMEDCT_US|Adult type granulosa cell tumor of testis|8620/1
C4542861|T191|PTGB|734274003|SNOMEDCT_US|Adult type granulosa cell tumour of testis|8620/1
C0018206|T191|PT|46585005|SNOMEDCT_US|Granulosa cell tumor|8620/1
C0018206|T191|SY|46585005|SNOMEDCT_US|Granulosa cell tumor, adult type|8620/1
C0018206|T191|IS|46585005|SNOMEDCT_US|Granulosa cell tumor, NOS|8620/1
C0018206|T191|PTGB|46585005|SNOMEDCT_US|Granulosa cell tumour|8620/1
C0018206|T191|SYGB|46585005|SNOMEDCT_US|Granulosa cell tumour, adult type|8620/1
C0018206|T191|SY|0000005693|CHV|cell granulosa tumor|8620/3
C0018206|T191|SY|0000005693|CHV|cells granulosa tumor|8620/3
C0018206|T191|PT|0000005693|CHV|granulosa cell tumor|8620/3
C0018206|T191|SY|0000005693|CHV|granulosa cell tumors|8620/3
C0018206|T191|SY|0000005693|CHV|granulosa cell tumour|8620/3
C0018206|T191|SY|0000005693|CHV|tumor cell granulosa|8620/3
C0334401|T191|PT|MTHU014761|ICPC2ICD10ENG|carcinoma; granulosa cell|8620/3
C0334401|T191|PT|MTHU032839|ICPC2ICD10ENG|granulosa cell; carcinoma|8620/3
C0018206|T191|PT|MTHU032840|ICPC2ICD10ENG|granulosa cell; tumor|8620/3
C0334401|T191|PT|MTHU032842|ICPC2ICD10ENG|granulosa cell; tumor, malignant|8620/3
C0018206|T191|PT|MTHU077068|ICPC2ICD10ENG|tumor; granulosa cell|8620/3
C0334401|T191|PT|MTHU077070|ICPC2ICD10ENG|tumor; granulosa cell, malignant|8620/3
C0018206|T191|MH|D006106|MSH|Granulosa Cell Tumor|8620/3
C0018206|T191|PM|D006106|MSH|Granulosa Cell Tumors|8620/3
C0018206|T191|PM|D006106|MSH|Tumor, Granulosa Cell|8620/3
C0018206|T191|PM|D006106|MSH|Tumors, Granulosa Cell|8620/3
C0018206|T191|PN|NOCODE|MTH|granulosa cell tumor|8620/3
C0334401|T191|PN|NOCODE|MTH|Malignant Granulosa Cell Tumor|8620/3
C0018206|T191|SY|C3070|NCI|Granulosa Cell Neoplasm|8620/3
C0018206|T191|PT|C3070|NCI|Granulosa Cell Tumor|8620/3
C0334401|T191|SY|C4205|NCI|Malignant Granulosa Cell Neoplasm|8620/3
C0334401|T191|PT|C4205|NCI|Malignant Granulosa Cell Tumor|8620/3
C0334401|T191|PT|C4205|NCI_CDISC|GRANULOSA CELL TUMOR, MALIGNANT|8620/3
C0334401|T191|SY|C4205|NCI_CDISC|Malignant Granulosa Cell Tumor|8620/3
C0018206|T191|PT|CDR0000044780|NCI_NCI-GLOSS|granulosa cell tumor|8620/3
C0018206|T191|PT|C3070|NCI_NICHD|Granulosa Cell Tumor|8620/3
C0334401|T191|SY|BBC4.|RCD|Granulosa cell carcinoma|8620/3
C0018206|T191|PT|Xa99G|RCD|Granulosa cell tumour|8620/3
C0334401|T191|AB|BBC4.|RCD|Malign granulosa cell tumour|8620/3
C0334401|T191|PT|BBC4.|RCD|Malignant granulosa cell tumour|8620/3
C0018206|T191|PT|Xa99G|RCDAE|Granulosa cell tumor|8620/3
C0334401|T191|AB|BBC4.|RCDAE|Malign granulosa cell tumor|8620/3
C0334401|T191|PT|BBC4.|RCDAE|Malignant granulosa cell tumor|8620/3
C0018206|T191|OP|BBC3.|RCDSA|Granulosa cell tumor NOS|8620/3
C0018206|T191|OP|BBC3.|RCDSY|Granulosa cell tumour NOS|8620/3
C0334401|T191|SY|18861007|SNOMEDCT_US|Granulosa cell carcinoma|8620/3
C0018206|T191|PT|46585005|SNOMEDCT_US|Granulosa cell tumor|8620/3
C0018206|T191|SY|46585005|SNOMEDCT_US|Granulosa cell tumor, adult type|8620/3
C0334401|T191|PT|18861007|SNOMEDCT_US|Granulosa cell tumor, malignant|8620/3
C0018206|T191|IS|46585005|SNOMEDCT_US|Granulosa cell tumor, NOS|8620/3
C0334401|T191|SY|18861007|SNOMEDCT_US|Granulosa cell tumor, sarcomatoid|8620/3
C0018206|T191|PTGB|46585005|SNOMEDCT_US|Granulosa cell tumour|8620/3
C0018206|T191|SYGB|46585005|SNOMEDCT_US|Granulosa cell tumour, adult type|8620/3
C0334401|T191|PTGB|18861007|SNOMEDCT_US|Granulosa cell tumour, malignant|8620/3
C0334401|T191|SYGB|18861007|SNOMEDCT_US|Granulosa cell tumour, sarcomatoid|8620/3
C0334401|T191|SY|18861007|SNOMEDCT_US|Malignant granulosa cell tumor|8620/3
C0334401|T191|SYGB|18861007|SNOMEDCT_US|Malignant granulosa cell tumour|8620/3
C0334402|T191|SY|0000029971|CHV|cell granulosa theca tumor|8621/1
C0334402|T191|SY|0000029971|CHV|cell granulosa theca tumors|8621/1
C0334402|T191|PT|0000029971|CHV|granulosa cell-theca cell tumor|8621/1
C0334402|T191|PT|MTHU032843|ICPC2ICD10ENG|granulosa cell-theca cell; tumor|8621/1
C0334402|T191|PT|MTHU073985|ICPC2ICD10ENG|theca cell-granulosa cell; tumor|8621/1
C0334402|T191|PT|MTHU077071|ICPC2ICD10ENG|tumor; granulosa cell-theca cell|8621/1
C0334402|T191|PT|MTHU077163|ICPC2ICD10ENG|tumor; theca cell-granulosa cell|8621/1
C0334402|T191|OP|C66751|NCI|Granulosa Cell-Theca Cell Tumor|8621/1
C0334402|T191|PT|C66751|NCI|Granulosa Cell-Theca Cell Tumor|8621/1
C0334402|T191|PT|BBC5.|RCD|Granulosa cell - theca cell tumour|8621/1
C0334402|T191|AB|BBC5.|RCD|Granulosa cell-theca cell tum|8621/1
C0334402|T191|SY|BBC5.|RCD|Theca cell - granulosa cell tumour|8621/1
C0334402|T191|AB|BBC5.|RCD|Theca cell-granulosa cell tum|8621/1
C0334402|T191|PT|BBC5.|RCDAE|Granulosa cell - theca cell tumor|8621/1
C0334402|T191|SY|BBC5.|RCDAE|Theca cell - granulosa cell tumor|8621/1
C0334402|T191|SY|31296004|SNOMEDCT_US|Granulosa cell - theca cell tumor|8621/1
C0334402|T191|SYGB|31296004|SNOMEDCT_US|Granulosa cell - theca cell tumour|8621/1
C0334402|T191|PT|31296004|SNOMEDCT_US|Granulosa cell-theca cell tumor|8621/1
C0334402|T191|PTGB|31296004|SNOMEDCT_US|Granulosa cell-theca cell tumour|8621/1
C0334402|T191|SY|31296004|SNOMEDCT_US|Theca cell - granulosa cell tumor|8621/1
C0334402|T191|SYGB|31296004|SNOMEDCT_US|Theca cell - granulosa cell tumour|8621/1
C0334402|T191|SY|31296004|SNOMEDCT_US|Theca cell-granulosa cell tumor|8621/1
C0334402|T191|SYGB|31296004|SNOMEDCT_US|Theca cell-granulosa cell tumour|8621/1
C0334403|T191|PT|0000029972|CHV|juvenile granulosa cell tumor|8622/1
C0334403|T191|PT|MTHU032841|ICPC2ICD10ENG|granulosa cell; tumor, juvenile|8622/1
C0334403|T191|PT|MTHU040684|ICPC2ICD10ENG|juvenile; granulosa cell tumor|8622/1
C0334403|T191|PT|MTHU077069|ICPC2ICD10ENG|tumor; granulosa cell, juvenile|8622/1
C0334403|T191|SY|C4207|NCI|Juvenile Type Granulosa Cell Neoplasm|8622/1
C0334403|T191|PT|C4207|NCI|Juvenile Type Granulosa Cell Tumor|8622/1
C0334403|T191|PT|C4207|NCI_NICHD|Juvenile Type Granulosa Cell Tumor|8622/1
C0334403|T191|PT|X77o9|RCD|Juvenile granulosa cell tumour|8622/1
C0334403|T191|PT|X77o9|RCDAE|Juvenile granulosa cell tumor|8622/1
C0334403|T191|AB|X77o9|RCDSY|Juvenil granulos cell tumur|8622/1
C0334403|T191|OAP|189735004|SNOMEDCT_US|Juvenile granulosa cell tumor|8622/1
C0334403|T191|PT|77029009|SNOMEDCT_US|Juvenile granulosa cell tumor|8622/1
C0334403|T191|OAP|189735004|SNOMEDCT_US|Juvenile granulosa cell tumour|8622/1
C0334403|T191|OF|189735004|SNOMEDCT_US|Juvenile granulosa cell tumour|8622/1
C0334403|T191|PTGB|77029009|SNOMEDCT_US|Juvenile granulosa cell tumour|8622/1
C0334404|T191|PT|MTHU067627|ICPC2ICD10ENG|sex cord; tumor, with annular tubules|8623/1
C0334404|T191|PT|MTHU077156|ICPC2ICD10ENG|tumor; sex cord, with annular tubules|8623/1
C1519276|T191|SY|C4208|NCI|Ovarian Sertoli Cell Tumor, Annular Tubular Variant|8623/1
C1519276|T191|SY|C4208|NCI|Ovarian Sex Cord Neoplasm with Annular Tubules|8623/1
C1519276|T191|PT|C4208|NCI|Ovarian Sex Cord Tumor with Annular Tubules|8623/1
C0334404|T191|AB|X77oA|RCD|Sex cord tum + annular tubules|8623/1
C0334404|T191|PT|X77oA|RCD|Sex cord tumour with annular tubules|8623/1
C0334404|T191|PT|X77oA|RCDAE|Sex cord tumor with annular tubules|8623/1
C0334404|T191|AB|X77oA|RCDSY|Sex cord tum+annular tubule|8623/1
C0334404|T191|OAP|189726006|SNOMEDCT_US|Sex cord tumor with annular tubules|8623/1
C0334404|T191|PT|72457004|SNOMEDCT_US|Sex cord tumor with annular tubules|8623/1
C0334404|T191|OAP|189726006|SNOMEDCT_US|Sex cord tumour with annular tubules|8623/1
C0334404|T191|OF|189726006|SNOMEDCT_US|Sex cord tumour with annular tubules|8623/1
C0334404|T191|PTGB|72457004|SNOMEDCT_US|Sex cord tumour with annular tubules|8623/1
C1879826|T191|PN|NOCODE|MTH|Benign Sertoli Cell Tumor|8630/0
C0334405|T191|PN|NOCODE|MTH|Well Differentiated Ovarian Sertoli-Leydig Cell Tumor|8630/0
C1879826|T191|PT|C67012|NCI|Benign Sertoli Cell Tumor|8630/0
C0334405|T191|PT|C4209|NCI|Well Differentiated Ovarian Sertoli-Leydig Cell Tumor|8630/0
C1879826|T191|SY|C67012|NCI_CDISC|Benign Androblastoma|8630/0
C1879826|T191|PT|C67012|NCI_CDISC|SERTOLI CELL TUMOR, BENIGN|8630/0
C0334405|T191|PT|BBC60|RCD|Benign androblastoma|8630/0
C0334405|T191|SY|BBC60|RCD|Benign arrhenoblastoma|8630/0
C0334405|T191|PT|83802009|SNOMEDCT_US|Androblastoma, benign|8630/0
C0334405|T191|SY|83802009|SNOMEDCT_US|Arrhenoblastoma, benign|8630/0
C0334405|T191|SY|83802009|SNOMEDCT_US|Benign androblastoma|8630/0
C0334405|T191|SY|83802009|SNOMEDCT_US|Benign arrhenoblastoma|8630/0
C0003810|T191|SY|0000001439|CHV|androblastoma|8630/1
C0003810|T191|SY|0000001439|CHV|androblastomas|8630/1
C0003810|T191|PT|0000001439|CHV|arrhenoblastoma|8630/1
C0003810|T191|PT|0000031051|CHV|arrhenoblastoma of ovary|8630/1
C0003810|T191|SY|0000001439|CHV|arrhenoblastomas|8630/1
C0003810|T191|SY|0000031051|CHV|cell ovary sertoli-leydig tumor|8630/1
C0036769|T191|SY|0000011228|CHV|cell sertoli tumors|8630/1
C0036769|T191|PT|0000011228|CHV|sertoli cell tumor|8630/1
C0036769|T191|SY|0000011228|CHV|sertoli cell tumour|8630/1
C0036769|T191|ET|2016-2999|CSP|Sertoli cell tumor|8630/1
C0003810|T191|LLT|10073278|MDR|Ovarian Sertoli-Leydig cell tumor|8630/1
C0003810|T191|MTH_PT|10073270|MDR|Ovarian Sertoli-Leydig cell tumor|8630/1
C0003810|T191|LLT|10073270|MDR|Ovarian Sertoli-Leydig cell tumour|8630/1
C0003810|T191|PT|10073270|MDR|Ovarian Sertoli-Leydig cell tumour|8630/1
C0036769|T191|PT|31526|MEDCIN|adenoma of testis|8630/1
C0003810|T191|PT|31609|MEDCIN|malignant arrhenoblastoma of ovary|8630/1
C0003810|T191|SY|351076|MEDCIN|ovarian malignant neoplasm sertoli-leydig tumor|8630/1
C0003810|T191|PT|351076|MEDCIN|Sertoli-Leydig cell tumor of ovary|8630/1
C0036769|T191|SY|31526|MEDCIN|testicular adenoma|8630/1
C0003810|T191|NM|C537588|MSH|Androblastoma of ovary|8630/1
C0036769|T191|MH|D012707|MSH|Sertoli Cell Tumor|8630/1
C0003810|T191|CE|C537588|MSH|Sertoli-leydig cell tumor of the ovary|8630/1
C0036769|T191|PM|D012707|MSH|Tumor, Sertoli Cell|8630/1
C0036769|T191|PN|NOCODE|MTH|Sertoli Cell Tumor|8630/1
C0003810|T191|PN|NOCODE|MTH|Sertoli-Leydig cell tumor of ovary|8630/1
C0003810|T191|SY|C2880|NCI|Androblastoma|8630/1
C0003810|T191|SY|C2880|NCI|Arrhenoblastoma|8630/1
C0003810|T191|SY|C2880|NCI|Ovarian Sertoli-Leydig Cell Neoplasm|8630/1
C0003810|T191|PT|C2880|NCI|Ovarian Sertoli-Leydig Cell Tumor|8630/1
C0036769|T191|PT|C39976|NCI|Sertoli Cell Tumor|8630/1
C0003810|T191|SY|C2880|NCI|Sertoli-Leydig Cell Tumor of Ovary|8630/1
C0003810|T191|SY|C2880|NCI|Sertoli-Leydig Cell Tumor of the Ovary|8630/1
C0003810|T191|SY|C2880|NCI|Sertoli-Leydig Neoplasm of Ovary|8630/1
C0003810|T191|SY|C2880|NCI|Sertoli-Leydig Neoplasm of the Ovary|8630/1
C0003810|T191|PT|CDR0000407749|NCI_NCI-GLOSS|androblastoma|8630/1
C0003810|T191|PT|CDR0000407750|NCI_NCI-GLOSS|arrhenoblastoma|8630/1
C0003810|T191|PT|CDR0000407748|NCI_NCI-GLOSS|Sertoli-Leydig cell tumor of the ovary|8630/1
C0003810|T191|PT|C2880|NCI_NICHD|Ovarian Sertoli-Leydig Cell Tumor|8630/1
C0036769|T191|PT|C39976|NCI_NICHD|Sertoli Cell Tumor|8630/1
C0003810|T191|PT|BBC6.|RCD|Androblastoma|8630/1
C0003810|T191|SY|BBC6.|RCD|Arrhenoblastoma|8630/1
C0003810|T191|SY|X78X4|RCD|Arrhenoblastoma of ovary|8630/1
C0036769|T191|SY|Xa99J|RCD|Pick's tubular adenoma|8630/1
C0036769|T191|SY|Xa99J|RCD|Sertoli cell adenoma|8630/1
C0036769|T191|PT|Xa99J|RCD|Sertoli cell tumour|8630/1
C0003810|T191|AB|X78X4|RCD|Sertoli-Leydig cell tum ovary|8630/1
C0003810|T191|PT|X78X4|RCD|Sertoli-Leydig cell tumour of ovary|8630/1
C0036769|T191|SY|Xa99J|RCD|Testicular adenoma|8630/1
C0036769|T191|SY|Xa99J|RCD|Tubular androblastoma|8630/1
C0036769|T191|PT|Xa99J|RCDAE|Sertoli cell tumor|8630/1
C0003810|T191|PT|X78X4|RCDAE|Sertoli-Leydig cell tumor of ovary|8630/1
C0003810|T191|OP|BBC6z|RCDSY|Androblastoma NOS|8630/1
C0036769|T191|OP|BBC9.|RCDSY|Tubular androblastoma NOS|8630/1
C0003810|T191|PT|62283005|SNOMEDCT_US|Androblastoma|8630/1
C0003810|T191|SY|62283005|SNOMEDCT_US|Androblastoma, no ICD-O subtype|8630/1
C0003810|T191|SY|62283005|SNOMEDCT_US|Androblastoma, no International Classification of Diseases for Oncology subtype|8630/1
C0003810|T191|IS|62283005|SNOMEDCT_US|Androblastoma, NOS|8630/1
C0003810|T191|SY|62283005|SNOMEDCT_US|Arrhenoblastoma|8630/1
C0003810|T191|SY|254866007|SNOMEDCT_US|Arrhenoblastoma of ovary|8630/1
C0003810|T191|IS|62283005|SNOMEDCT_US|Arrhenoblastoma, NOS|8630/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Pick tubular adenoma|8630/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Pick's tubular adenoma|8630/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sertoli cell adenoma|8630/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Sertoli cell adenoma|8630/1
C0036769|T191|OAP|89089007|SNOMEDCT_US|Sertoli cell tumor|8630/1
C0036769|T191|PT|128857001|SNOMEDCT_US|Sertoli cell tumor|8630/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sertoli cell tumor -RETIRED-|8630/1
C0036769|T191|OF|89089007|SNOMEDCT_US|Sertoli cell tumor -RETIRED-|8630/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Sertoli cell tumor, no ICD-O subtype|8630/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Sertoli cell tumor, no International Classification of Diseases for Oncology subtype|8630/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sertoli cell tumor, NOS|8630/1
C0036769|T191|OAP|89089007|SNOMEDCT_US|Sertoli cell tumour|8630/1
C0036769|T191|PTGB|128857001|SNOMEDCT_US|Sertoli cell tumour|8630/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sertoli cell tumour -RETIRED-|8630/1
C0036769|T191|SYGB|128857001|SNOMEDCT_US|Sertoli cell tumour, no ICD-O subtype|8630/1
C0003810|T191|PT|254866007|SNOMEDCT_US|Sertoli-Leydig cell tumor of ovary|8630/1
C0003810|T191|PTGB|254866007|SNOMEDCT_US|Sertoli-Leydig cell tumour of ovary|8630/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sustentacular cell tumor|8630/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Testicular adenoma|8630/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Testicular adenoma|8630/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Tubular androblastoma|8630/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Tubular androblastoma, NOS|8630/1
C0334406|T191|PT|271488|MEDCIN|malignant androblastoma|8630/3
C0334406|T191|PN|NOCODE|MTH|Malignant Sertoli Cell Tumor|8630/3
C0334406|T191|PT|C67006|NCI|Malignant Sertoli Cell Tumor|8630/3
C0334406|T191|SY|C67006|NCI_CDISC|Malignant Androblastoma|8630/3
C0334406|T191|PT|C67006|NCI_CDISC|SERTOLI CELL TUMOR, MALIGNANT|8630/3
C0334406|T191|PT|BBC61|RCD|Malignant androblastoma|8630/3
C0334406|T191|SY|BBC61|RCD|Malignant arrhenoblastoma|8630/3
C0334406|T191|PT|12323008|SNOMEDCT_US|Androblastoma, malignant|8630/3
C0334406|T191|SY|12323008|SNOMEDCT_US|Arrhenoblastoma, malignant|8630/3
C0334406|T191|SY|12323008|SNOMEDCT_US|Malignant androblastoma|8630/3
C0334406|T191|SY|12323008|SNOMEDCT_US|Malignant arrhenoblastoma|8630/3
C0334405|T191|PN|NOCODE|MTH|Well Differentiated Ovarian Sertoli-Leydig Cell Tumor|8631/0
C0334405|T191|PT|C4209|NCI|Well Differentiated Ovarian Sertoli-Leydig Cell Tumor|8631/0
C0334405|T191|PT|BBC60|RCD|Benign androblastoma|8631/0
C0334405|T191|SY|BBC60|RCD|Benign arrhenoblastoma|8631/0
C0334405|T191|PT|83802009|SNOMEDCT_US|Androblastoma, benign|8631/0
C0334405|T191|SY|83802009|SNOMEDCT_US|Arrhenoblastoma, benign|8631/0
C0334405|T191|SY|83802009|SNOMEDCT_US|Benign androblastoma|8631/0
C0334405|T191|SY|83802009|SNOMEDCT_US|Benign arrhenoblastoma|8631/0
C1314745|T191|PT|34110004|SNOMEDCT_US|Sertoli-Leydig cell tumor, well differentiated|8631/0
C1314745|T191|PTGB|34110004|SNOMEDCT_US|Sertoli-Leydig cell tumour, well differentiated|8631/0
C1318541|T191|PN|NOCODE|MTH|Sertoli-Leydig cell tumor of intermediate differentiation|8631/1
C1512860|T191|SY|C39968|NCI|Intermediate Differentiated Ovarian Sertoli-Leydig Cell Tumor|8631/1
C1512860|T191|PT|C39968|NCI|Moderately Differentiated Ovarian Sertoli-Leydig Cell Tumor|8631/1
C1318541|T191|SY|128905000|SNOMEDCT_US|Sertoli-Leydig cell tumor|8631/1
C1318541|T191|PT|128905000|SNOMEDCT_US|Sertoli-Leydig cell tumor of intermediate differentiation|8631/1
C1318541|T191|SY|128905000|SNOMEDCT_US|Sertoli-Leydig cell tumor, moderately differentiated|8631/1
C1318541|T191|SYGB|128905000|SNOMEDCT_US|Sertoli-Leydig cell tumour|8631/1
C1318541|T191|PTGB|128905000|SNOMEDCT_US|Sertoli-Leydig cell tumour of intermediate differentiation|8631/1
C1318541|T191|SYGB|128905000|SNOMEDCT_US|Sertoli-Leydig cell tumour, moderately differentiated|8631/1
C1879314|T191|PT|233163|MEDCIN|poorly differentiated Sertoli-Leydig cell tumor of ovary|8631/3
C1879314|T191|PN|NOCODE|MTH|Poorly Differentiated Ovarian Sertoli-Leydig Cell Tumor|8631/3
C1879314|T191|PT|C4210|NCI|Poorly Differentiated Ovarian Sertoli-Leydig Cell Tumor|8631/3
C1266105|T191|PT|128906004|SNOMEDCT_US|Sertoli-Leydig cell tumor, poorly differentiated|8631/3
C1266105|T191|SY|128906004|SNOMEDCT_US|Sertoli-Leydig cell tumor, sarcomatoid|8631/3
C1266105|T191|PTGB|128906004|SNOMEDCT_US|Sertoli-Leydig cell tumour, poorly differentiated|8631/3
C1266105|T191|SYGB|128906004|SNOMEDCT_US|Sertoli-Leydig cell tumour, sarcomatoid|8631/3
C0018413|T191|PEP|D018312|MSH|Gynandroblastoma|8632/1
C0018413|T191|PM|D018312|MSH|Gynandroblastomas|8632/1
C0346178|T191|NM|C538459|MSH|Ovarian gynandroblastoma|8632/1
C0018413|T191|PN|NOCODE|MTH|Gynandroblastoma|8632/1
C0346178|T191|PN|NOCODE|MTH|Ovarian gynandroblastoma|8632/1
C0346178|T191|SY|C3072|NCI|Gynandroblastoma|8632/1
C0346178|T191|SY|C3072|NCI|Gynandroblastoma of Ovary|8632/1
C0346178|T191|SY|C3072|NCI|Gynandroblastoma of the Ovary|8632/1
C0346178|T191|PT|C3072|NCI|Ovarian Gynandroblastoma|8632/1
C0018413|T191|PT|BBC8.|RCD|Gynandroblastoma|8632/1
C0346178|T191|PT|X78X5|RCD|Gynandroblastoma of ovary|8632/1
C0018413|T191|PT|26735007|SNOMEDCT_US|Gynandroblastoma|8632/1
C0346178|T191|PT|254867003|SNOMEDCT_US|Gynandroblastoma of ovary|8632/1
C1518728|T191|PT|C39971|NCI|Ovarian Retiform Sertoli-Leydig Cell Tumor|8633/1
C1266106|T191|PT|128724009|SNOMEDCT_US|Sertoli-Leydig cell tumor, retiform|8633/1
C1266106|T191|PTGB|128724009|SNOMEDCT_US|Sertoli-Leydig cell tumour, retiform|8633/1
C1512861|T191|SY|C39972|NCI|Intermediate Differentiated Ovarian Sertoli-Leydig Cell Tumor, Variant with Heterologous Elements|8634/1
C1512861|T191|PT|C39972|NCI|Moderately Differentiated Ovarian Sertoli-Leydig Cell Tumor, Variant with Heterologous Elements|8634/1
C1266107|T191|PT|128725005|SNOMEDCT_US|Sertoli-Leydig cell tumor, intermediate differentiation, with heterologous elements|8634/1
C1266107|T191|SY|128725005|SNOMEDCT_US|Sertoli-Leydig cell tumor, moderately differentiated, with heterologous elements|8634/1
C1266107|T191|SY|128725005|SNOMEDCT_US|Sertoli-Leydig cell tumor, retiform, with heterologous elements|8634/1
C1266107|T191|PTGB|128725005|SNOMEDCT_US|Sertoli-Leydig cell tumour, intermediate differentiation, with heterologous elements|8634/1
C1266107|T191|SYGB|128725005|SNOMEDCT_US|Sertoli-Leydig cell tumour, moderately differentiated, with heterologous elements|8634/1
C1266107|T191|SYGB|128725005|SNOMEDCT_US|Sertoli-Leydig cell tumour, retiform, with heterologous elements|8634/1
C1514226|T191|PT|C39973|NCI|Poorly Differentiated Ovarian Sertoli-Leydig Cell Tumor, Variant with Heterologous Elements|8634/3
C1266108|T191|PT|128727002|SNOMEDCT_US|Sertoli-Leydig cell tumor, poorly differentiated, with heterologous elements|8634/3
C1266108|T191|PTGB|128727002|SNOMEDCT_US|Sertoli-Leydig cell tumour, poorly differentiated, with heterologous elements|8634/3
C0036769|T191|SY|0000011228|CHV|cell sertoli tumors|8640/1
C0036769|T191|PT|0000011228|CHV|sertoli cell tumor|8640/1
C0036769|T191|SY|0000011228|CHV|sertoli cell tumour|8640/1
C0036769|T191|ET|2016-2999|CSP|Sertoli cell tumor|8640/1
C0036769|T191|PT|31526|MEDCIN|adenoma of testis|8640/1
C0036769|T191|SY|31526|MEDCIN|testicular adenoma|8640/1
C0036769|T191|MH|D012707|MSH|Sertoli Cell Tumor|8640/1
C0036769|T191|PM|D012707|MSH|Tumor, Sertoli Cell|8640/1
C0036769|T191|PN|NOCODE|MTH|Sertoli Cell Tumor|8640/1
C0036769|T191|PT|C39976|NCI|Sertoli Cell Tumor|8640/1
C0036769|T191|PT|C39976|NCI_NICHD|Sertoli Cell Tumor|8640/1
C0036769|T191|SY|Xa99J|RCD|Pick's tubular adenoma|8640/1
C0036769|T191|SY|Xa99J|RCD|Sertoli cell adenoma|8640/1
C0036769|T191|PT|Xa99J|RCD|Sertoli cell tumour|8640/1
C0036769|T191|SY|Xa99J|RCD|Testicular adenoma|8640/1
C0036769|T191|SY|Xa99J|RCD|Tubular androblastoma|8640/1
C0036769|T191|PT|Xa99J|RCDAE|Sertoli cell tumor|8640/1
C0036769|T191|OP|BBC9.|RCDSY|Tubular androblastoma NOS|8640/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Pick tubular adenoma|8640/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Pick's tubular adenoma|8640/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Sertoli cell adenoma|8640/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sertoli cell adenoma|8640/1
C0036769|T191|PT|128857001|SNOMEDCT_US|Sertoli cell tumor|8640/1
C0036769|T191|OAP|89089007|SNOMEDCT_US|Sertoli cell tumor|8640/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sertoli cell tumor -RETIRED-|8640/1
C0036769|T191|OF|89089007|SNOMEDCT_US|Sertoli cell tumor -RETIRED-|8640/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Sertoli cell tumor, no ICD-O subtype|8640/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Sertoli cell tumor, no International Classification of Diseases for Oncology subtype|8640/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sertoli cell tumor, NOS|8640/1
C0036769|T191|OAP|89089007|SNOMEDCT_US|Sertoli cell tumour|8640/1
C0036769|T191|PTGB|128857001|SNOMEDCT_US|Sertoli cell tumour|8640/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sertoli cell tumour -RETIRED-|8640/1
C0036769|T191|SYGB|128857001|SNOMEDCT_US|Sertoli cell tumour, no ICD-O subtype|8640/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Sustentacular cell tumor|8640/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Testicular adenoma|8640/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Testicular adenoma|8640/1
C0036769|T191|SY|128857001|SNOMEDCT_US|Tubular androblastoma|8640/1
C0036769|T191|IS|89089007|SNOMEDCT_US|Tubular androblastoma, NOS|8640/1
C0334406|T191|PT|271488|MEDCIN|malignant androblastoma|8640/3
C0334406|T191|PN|NOCODE|MTH|Malignant Sertoli Cell Tumor|8640/3
C0334406|T191|PT|C67006|NCI|Malignant Sertoli Cell Tumor|8640/3
C0334406|T191|SY|C67006|NCI_CDISC|Malignant Androblastoma|8640/3
C0334406|T191|PT|C67006|NCI_CDISC|SERTOLI CELL TUMOR, MALIGNANT|8640/3
C0334406|T191|PT|BBC61|RCD|Malignant androblastoma|8640/3
C0334406|T191|SY|BBC61|RCD|Malignant arrhenoblastoma|8640/3
C0334407|T191|PT|BBCA.|RCD|Sertoli cell carcinoma|8640/3
C0334406|T191|PT|12323008|SNOMEDCT_US|Androblastoma, malignant|8640/3
C0334406|T191|SY|12323008|SNOMEDCT_US|Arrhenoblastoma, malignant|8640/3
C0334406|T191|SY|12323008|SNOMEDCT_US|Malignant androblastoma|8640/3
C0334406|T191|SY|12323008|SNOMEDCT_US|Malignant arrhenoblastoma|8640/3
C0334407|T191|PT|80091008|SNOMEDCT_US|Sertoli cell carcinoma|8640/3
C1515296|T191|PT|C39943|NCI|Testicular Sertoli Cell Tumor, Lipid Rich Variant|8641/0
C0334408|T191|SY|BBCB.|RCD|Folliculome lipidique|8641/0
C0334408|T191|AB|BBCB.|RCD|Sertoli cell tum+lipid storage|8641/0
C0334408|T191|PT|BBCB.|RCD|Sertoli cell tumour with lipid storage|8641/0
C0334408|T191|AB|BBCB.|RCD|Tubul androblastoma+lipid stor|8641/0
C0334408|T191|SY|BBCB.|RCD|Tubular androblastoma with lipid storage|8641/0
C0334408|T191|PT|BBCB.|RCDAE|Sertoli cell tumor with lipid storage|8641/0
C0334408|T191|SY|24815001|SNOMEDCT_US|Folliculome lipidique|8641/0
C0334408|T191|SY|24815001|SNOMEDCT_US|Lipid-rich Sertoli cell tumor|8641/0
C0334408|T191|SYGB|24815001|SNOMEDCT_US|Lipid-rich Sertoli cell tumour|8641/0
C0334408|T191|PT|24815001|SNOMEDCT_US|Sertoli cell tumor with lipid storage|8641/0
C0334408|T191|PTGB|24815001|SNOMEDCT_US|Sertoli cell tumour with lipid storage|8641/0
C0334408|T191|SY|24815001|SNOMEDCT_US|Tubular androblastoma with lipid storage|8641/0
C1515287|T191|PT|C39944|NCI|Testicular Large Cell Calcifying Sertoli Cell Tumor|8642/1
C1266109|T191|PT|128728007|SNOMEDCT_US|Large cell calcifying Sertoli cell tumor|8642/1
C1266109|T191|PTGB|128728007|SNOMEDCT_US|Large cell calcifying Sertoli cell tumour|8642/1
C0334409|T191|PN|NOCODE|MTH|Leydig cell tumor, benign|8650/0
C0334409|T191|SY|C4212|NCI|Benign Interstitial Cell Neoplasm|8650/0
C0334409|T191|SY|C4212|NCI|Benign Interstitial Cell Tumor|8650/0
C0334409|T191|SY|C4212|NCI|Benign Leydig Cell Neoplasm|8650/0
C0334409|T191|PT|C4212|NCI|Benign Leydig Cell Tumor|8650/0
C0334409|T191|SY|C4212|NCI_CDISC|Adenoma, Interstitial|8650/0
C0334409|T191|SY|C4212|NCI_CDISC|Adenoma, Leydig Cell|8650/0
C0334409|T191|SY|C4212|NCI_CDISC|Benign Interstitial Cell Neoplasm|8650/0
C0334409|T191|SY|C4212|NCI_CDISC|Benign Interstitial Cell Tumor|8650/0
C0334409|T191|SY|C4212|NCI_CDISC|Benign Leydig Cell Neoplasm|8650/0
C0334409|T191|PT|C4212|NCI_CDISC|LEYDIG CELL TUMOR, BENIGN|8650/0
C0334409|T191|AB|BBCC0|RCD|Benign interstitial cell tum|8650/0
C0334409|T191|SY|BBCC0|RCD|Benign interstitial cell tumour|8650/0
C0334409|T191|PT|BBCC0|RCD|Benign Leydig cell tumour|8650/0
C0334409|T191|SY|BBCC0|RCDAE|Benign interstitial cell tumor|8650/0
C0334409|T191|PT|BBCC0|RCDAE|Benign Leydig cell tumor|8650/0
C0334409|T191|SY|5014008|SNOMEDCT_US|Benign interstitial cell tumor|8650/0
C0334409|T191|SYGB|5014008|SNOMEDCT_US|Benign interstitial cell tumour|8650/0
C0334409|T191|SY|5014008|SNOMEDCT_US|Benign Leydig cell tumor|8650/0
C0334409|T191|SYGB|5014008|SNOMEDCT_US|Benign Leydig cell tumour|8650/0
C0334409|T191|SY|5014008|SNOMEDCT_US|Interstitial cell tumor|8650/0
C0334409|T191|SY|5014008|SNOMEDCT_US|Interstitial cell tumor, benign|8650/0
C0334409|T191|SYGB|5014008|SNOMEDCT_US|Interstitial cell tumour|8650/0
C0334409|T191|SYGB|5014008|SNOMEDCT_US|Interstitial cell tumour, benign|8650/0
C0334409|T191|SY|5014008|SNOMEDCT_US|Leydig cell tumor|8650/0
C0334409|T191|PT|5014008|SNOMEDCT_US|Leydig cell tumor, benign|8650/0
C0334409|T191|SY|5014008|SNOMEDCT_US|Leydig cell tumor, no ICD-O subtype|8650/0
C0334409|T191|SYGB|5014008|SNOMEDCT_US|Leydig cell tumour|8650/0
C0334409|T191|PTGB|5014008|SNOMEDCT_US|Leydig cell tumour, benign|8650/0
C0334409|T191|SYGB|5014008|SNOMEDCT_US|Leydig cell tumour, no ICD-O subtype|8650/0
C0023601|T191|SY|0000007380|CHV|cell leydig tumors|8650/1
C0023601|T191|SY|0000007380|CHV|cell leydig tumour|8650/1
C0023601|T191|SY|0000007380|CHV|cells leydig tumor|8650/1
C0023601|T191|SY|0000007380|CHV|interstitial cell tumor|8650/1
C0023601|T191|PT|0000007380|CHV|leydig cell tumor|8650/1
C0023601|T191|SY|0000007380|CHV|leydig cell tumour|8650/1
C0023601|T191|ET|2016-2999|CSP|Leydig cell tumor|8650/1
C0023601|T191|SY|NOCODE|DXP|LEYDIG CELL TUMOR|8650/1
C0023601|T191|DI|U001833|DXP|TESTIS, INTERSTITIAL CELL TUMOR|8650/1
C0023601|T191|ET|D007984|MSH|Interstitial Cell Tumor|8650/1
C0023601|T191|PM|D007984|MSH|Interstitial Cell Tumors|8650/1
C0023601|T191|MH|D007984|MSH|Leydig Cell Tumor|8650/1
C0023601|T191|PM|D007984|MSH|Tumor, Interstitial Cell|8650/1
C0023601|T191|PM|D007984|MSH|Tumor, Leydig Cell|8650/1
C0023601|T191|PM|D007984|MSH|Tumors, Interstitial Cell|8650/1
C0023601|T191|PN|NOCODE|MTH|Leydig Cell Tumor|8650/1
C0023601|T191|SY|C3188|NCI|Interstitial Cell Neoplasm|8650/1
C0023601|T191|SY|C3188|NCI|Interstitial Cell Tumor|8650/1
C0023601|T191|SY|C3188|NCI|Leydig Cell Neoplasm|8650/1
C0023601|T191|PT|C3188|NCI|Leydig Cell Tumor|8650/1
C0023601|T191|DN|C3188|NCI_CTRP|Leydig Cell Tumor|8650/1
C0023601|T191|PT|C3188|NCI_NICHD|Leydig Cell Tumor|8650/1
C0023601|T191|SY|CDR0000686432|PDQ|interstitial cell neoplasm|8650/1
C0023601|T191|SY|CDR0000686432|PDQ|interstitial cell tumor|8650/1
C0023601|T191|SY|CDR0000686432|PDQ|leydig cell neoplasm|8650/1
C0023601|T191|PT|CDR0000686432|PDQ|Leydig cell tumor|8650/1
C0023601|T191|SY|BBCC.|RCD|Interstitial cell tumour|8650/1
C0023601|T191|PT|BBCC.|RCD|Leydig cell tumour|8650/1
C0023601|T191|SY|BBCC.|RCDAE|Interstitial cell tumor|8650/1
C0023601|T191|PT|BBCC.|RCDAE|Leydig cell tumor|8650/1
C0023601|T191|OP|BBCCz|RCDSA|Leydig cell tumor NOS|8650/1
C0023601|T191|OP|BBCCz|RCDSY|Leydig cell tumour NOS|8650/1
C0023601|T191|SY|45002009|SNOMEDCT_US|Interstitial cell tumor|8650/1
C0023601|T191|IS|45002009|SNOMEDCT_US|Interstitial cell tumor, NOS|8650/1
C0023601|T191|SYGB|45002009|SNOMEDCT_US|Interstitial cell tumour|8650/1
C0023601|T191|PT|45002009|SNOMEDCT_US|Leydig cell tumor|8650/1
C0023601|T191|SY|45002009|SNOMEDCT_US|Leydig cell tumor, no ICD-O subtype|8650/1
C0023601|T191|SY|45002009|SNOMEDCT_US|Leydig cell tumor, no International Classification of Diseases for Oncology subtype|8650/1
C0023601|T191|IS|45002009|SNOMEDCT_US|Leydig cell tumor, NOS|8650/1
C0023601|T191|PTGB|45002009|SNOMEDCT_US|Leydig cell tumour|8650/1
C0023601|T191|SYGB|45002009|SNOMEDCT_US|Leydig cell tumour, no ICD-O subtype|8650/1
C0334410|T191|PT|271489|MEDCIN|malignant Leydig cell tumor|8650/3
C0334410|T191|SY|C4213|NCI|Malignant Interstitial Cell Neoplasm|8650/3
C0334410|T191|SY|C4213|NCI|Malignant Interstitial Cell Tumor|8650/3
C0334410|T191|SY|C4213|NCI|Malignant Leydig Cell Neoplasm|8650/3
C0334410|T191|PT|C4213|NCI|Malignant Leydig Cell Tumor|8650/3
C0334410|T191|SY|C4213|NCI_CDISC|Carcinoma, Leydig Cell|8650/3
C0334410|T191|PT|C4213|NCI_CDISC|LEYDIG CELL TUMOR, MALIGNANT|8650/3
C0334410|T191|SY|C4213|NCI_CDISC|Malignant Interstitial Cell Neoplasm|8650/3
C0334410|T191|SY|C4213|NCI_CDISC|Malignant Interstitial Cell Tumor|8650/3
C0334410|T191|SY|C4213|NCI_CDISC|Malignant Leydig Cell Neoplasm|8650/3
C0334410|T191|AB|BBCC1|RCD|Malign interstitial cell tum|8650/3
C0334410|T191|SY|BBCC1|RCD|Malignant interstitial cell tumour|8650/3
C0334410|T191|PT|BBCC1|RCD|Malignant Leydig cell tumour|8650/3
C0334410|T191|SY|BBCC1|RCDAE|Malignant interstitial cell tumor|8650/3
C0334410|T191|PT|BBCC1|RCDAE|Malignant Leydig cell tumor|8650/3
C0334410|T191|SY|77870005|SNOMEDCT_US|Interstitial cell tumor, malignant|8650/3
C0334410|T191|SYGB|77870005|SNOMEDCT_US|Interstitial cell tumour, malignant|8650/3
C0334410|T191|PT|77870005|SNOMEDCT_US|Leydig cell tumor, malignant|8650/3
C0334410|T191|PTGB|77870005|SNOMEDCT_US|Leydig cell tumour, malignant|8650/3
C0334410|T191|SY|77870005|SNOMEDCT_US|Malignant interstitial cell tumor|8650/3
C0334410|T191|SYGB|77870005|SNOMEDCT_US|Malignant interstitial cell tumour|8650/3
C0334410|T191|SY|77870005|SNOMEDCT_US|Malignant Leydig cell tumor|8650/3
C0334410|T191|SYGB|77870005|SNOMEDCT_US|Malignant Leydig cell tumour|8650/3
C0346179|T191|PT|MTHU035145|ICPC2ICD10ENG|hilar cell; tumor|8660/0
C0346179|T191|PT|MTHU077073|ICPC2ICD10ENG|tumor; hilar cell|8660/0
C0346179|T191|SY|C4214|NCI|Hilar Cell Neoplasm|8660/0
C0346179|T191|SY|C4214|NCI|Hilar Cell Tumor of Ovary|8660/0
C0346179|T191|SY|C4214|NCI|Hilar Cell Tumor of the Ovary|8660/0
C0346179|T191|SY|C4214|NCI|Hilus Cell Neoplasm|8660/0
C0346179|T191|SY|C4214|NCI|Hilus Cell Tumor|8660/0
C0346179|T191|SY|C4214|NCI|Ovarian Hilar Cell Tumor|8660/0
C0346179|T191|PT|C4214|NCI|Ovarian Hilus Cell Tumor|8660/0
C0346179|T191|SY|BBCD.|RCD|Hilar cell tumour|8660/0
C0346179|T191|SY|BBCD.|RCD|Hilus cell tumour|8660/0
C0346179|T191|PT|X78X6|RCD|Hilus cell tumour of ovary|8660/0
C0346179|T191|SY|BBCD.|RCDAE|Hilar cell tumor|8660/0
C0346179|T191|SY|BBCD.|RCDAE|Hilus cell tumor|8660/0
C0346179|T191|PT|X78X6|RCDAE|Hilus cell tumor of ovary|8660/0
C0346179|T191|SY|11506001|SNOMEDCT_US|Hilar cell tumor|8660/0
C0346179|T191|SYGB|11506001|SNOMEDCT_US|Hilar cell tumour|8660/0
C0346179|T191|PT|11506001|SNOMEDCT_US|Hilus cell tumor|8660/0
C0346179|T191|PT|254868008|SNOMEDCT_US|Hilus cell tumor of ovary|8660/0
C0346179|T191|PTGB|11506001|SNOMEDCT_US|Hilus cell tumour|8660/0
C0346179|T191|PTGB|254868008|SNOMEDCT_US|Hilus cell tumour of ovary|8660/0
C0334412|T191|SY|0000029973|CHV|cell steroid tumors|8670/0
C0334412|T191|PT|0000029973|CHV|steroid cell tumor|8670/0
C0334412|T191|PT|MTHU077179|ICPC2ICD10ENG|tumor; fat cell, ovary|8670/0
C0334412|T191|PT|31613|MEDCIN|lipoid cell tumor of ovary|8670/0
C0334412|T191|SY|C4215|NCI|Lipid Cell Neoplasm of Ovary|8670/0
C0334412|T191|SY|C4215|NCI|Lipid Cell Neoplasm of the Ovary|8670/0
C0334412|T191|SY|C4215|NCI|Lipid Cell Tumor of Ovary|8670/0
C0334412|T191|SY|C4215|NCI|Lipid Cell Tumor of the Ovary|8670/0
C0334412|T191|SY|C4215|NCI|Ovarian Lipid Cell Neoplasm|8670/0
C0334412|T191|SY|C4215|NCI|Ovarian Lipid Cell Tumor|8670/0
C0334412|T191|SY|C4215|NCI|Ovarian Lipoid Cell Neoplasm|8670/0
C0334412|T191|SY|C4215|NCI|Ovarian Steroid Cell Neoplasm|8670/0
C0334412|T191|PT|C4215|NCI|Ovarian Steroid Cell Tumor|8670/0
C0334412|T191|SY|C4215|NCI|Steroid Cell Tumor of Ovary|8670/0
C0334412|T191|SY|C4215|NCI|Steroid Cell Tumor of the Ovary|8670/0
C0334412|T191|PT|BBCE.|RCD|Lipid cell tumour of ovary|8670/0
C0334412|T191|SY|BBCE.|RCD|Lipoid cell tumour of ovary|8670/0
C0334412|T191|SY|BBCE.|RCD|Masculinovoblastoma|8670/0
C0334412|T191|PT|BBCE.|RCDAE|Lipid cell tumor of ovary|8670/0
C0334412|T191|SY|BBCE.|RCDAE|Lipoid cell tumor of ovary|8670/0
C0334412|T191|PT|40761005|SNOMEDCT_US|Lipid cell tumor of ovary|8670/0
C0334412|T191|PTGB|40761005|SNOMEDCT_US|Lipid cell tumour of ovary|8670/0
C0334412|T191|SY|40761005|SNOMEDCT_US|Lipoid cell tumor of ovary|8670/0
C0334412|T191|SYGB|40761005|SNOMEDCT_US|Lipoid cell tumour of ovary|8670/0
C0334412|T191|SY|40761005|SNOMEDCT_US|Masculinovoblastoma|8670/0
C0334412|T191|SY|40761005|SNOMEDCT_US|Steroid cell tumor|8670/0
C0334412|T191|SYGB|40761005|SNOMEDCT_US|Steroid cell tumour|8670/0
C2212011|T191|PT|233162|MEDCIN|malignant steroid cell tumor of ovary|8670/3
C2212011|T191|PT|C39981|NCI|Malignant Ovarian Steroid Cell Tumor|8670/3
C1266110|T191|PT|128907008|SNOMEDCT_US|Steroid cell tumor, malignant|8670/3
C1266110|T191|PTGB|128907008|SNOMEDCT_US|Steroid cell tumour, malignant|8670/3
C0001630|T191|SY|0000000771|CHV|adrenal rest tumor|8671/0
C0001630|T191|PT|0000000771|CHV|adrenal rest tumour|8671/0
C0001630|T191|PT|31468|MEDCIN|adrenal benign rest tumor|8671/0
C0001630|T191|SY|31468|MEDCIN|adrenal rest tumor|8671/0
C0001630|T191|ET|D000314|MSH|Adrenal Cortical Rest Tumor|8671/0
C0001630|T191|MH|D000314|MSH|Adrenal Rest Tumor|8671/0
C0001630|T191|PM|D000314|MSH|Adrenal Rest Tumors|8671/0
C0001630|T191|PM|D000314|MSH|Rest Tumor, Adrenal|8671/0
C0001630|T191|PM|D000314|MSH|Rest Tumors, Adrenal|8671/0
C0001630|T191|PM|D000314|MSH|Tumor, Adrenal Rest|8671/0
C0001630|T191|PM|D000314|MSH|Tumors, Adrenal Rest|8671/0
C0001630|T191|SY|C2860|NCI|Adrenal Rest Neoplasm|8671/0
C0001630|T191|PT|C2860|NCI|Adrenal Rest Tumor|8671/0
C0001630|T191|PT|BBCF.|RCD|Adrenal rest tumour|8671/0
C0001630|T191|PT|BBCF.|RCDAE|Adrenal rest tumor|8671/0
C0001630|T191|PT|54292009|SNOMEDCT_US|Adrenal rest tumor|8671/0
C0001630|T191|PTGB|54292009|SNOMEDCT_US|Adrenal rest tumour|8671/0
C0346416|T191|AB|D3A|ICD10CM|Benign neuroendocrine tumors|8680/0
C0346416|T191|HT|D3A|ICD10CM|Benign neuroendocrine tumors|8680/0
C0346416|T191|LLT|10075443|MDR|Benign paraganglioma|8680/0
C0346416|T191|PT|333358|MEDCIN|benign neuroendocrine tumor|8680/0
C0346416|T191|PT|C48314|NCI|Benign Paraganglioma|8680/0
C0346416|T191|SY|C48314|NCI|Benign Paraganglionic Neoplasm|8680/0
C0346416|T191|SY|C48314|NCI_CDISC|Benign Neuroendocrine Cell Tumor|8680/0
C0346416|T191|SY|C48314|NCI_CDISC|Benign Paraganglionic Neoplasm|8680/0
C0346416|T191|PT|C48314|NCI_CDISC|PARAGANGLIOMA, BENIGN|8680/0
C0346416|T191|OP|X78du|RCD|Benign neuroendocrine tumour|8680/0
C0346416|T191|PT|XM1FK|RCD|Paraganglioma and glomus tumour|8680/0
C0346416|T191|AB|XM1FK|RCD|Paraganglioma+glomus tumour|8680/0
C0346416|T191|OP|X78du|RCDAE|Benign neuroendocrine tumor|8680/0
C0346416|T191|PT|XM1FK|RCDAE|Paraganglioma and glomus tumor|8680/0
C0346416|T191|AB|XM1FK|RCDAE|Paraganglioma+glomus tumor|8680/0
C0346416|T191|OA|BBD..|RCDSA|Paragangliom./glomus tumor|8680/0
C0346416|T191|OP|BBD..|RCDSA|Paragangliomas and glomus tumors|8680/0
C0346416|T191|OA|BBD..|RCDSY|Paragangliom./glomus tumour|8680/0
C0346416|T191|OP|BBD..|RCDSY|Paragangliomas and glomus tumours|8680/0
C0346416|T191|PT|255047001|SNOMEDCT_US|Benign neuroendocrine tumor|8680/0
C0346416|T191|PTGB|255047001|SNOMEDCT_US|Benign neuroendocrine tumour|8680/0
C0346416|T191|SY|107694002|SNOMEDCT_US|Paraganglioma and glomus tumor|8680/0
C0346416|T191|SYGB|107694002|SNOMEDCT_US|Paraganglioma and glomus tumour|8680/0
C0346416|T191|PT|107694002|SNOMEDCT_US|Paraganglioma, benign|8680/0
C0030421|T191|ET|0000004658|AOD|paraganglioma|8680/1
C0030421|T191|PT|0000009261|CHV|paraganglioma|8680/1
C0030421|T191|SY|0000009261|CHV|paragangliomas|8680/1
C0030421|T191|SY|HP:0002668|HPO|Carotid body tumors|8680/1
C0030421|T191|PT|HP:0002668|HPO|Paraganglioma|8680/1
C0030421|T191|SY|HP:0002668|HPO|Paragangliomas|8680/1
C0030421|T191|PT|MTHU030260|ICPC2ICD10ENG|gangliocytic; paraganglioma, unspecified site|8680/1
C0030421|T191|PT|MTHU057395|ICPC2ICD10ENG|paraganglioma; gangliocytic, unspecified site|8680/1
C0030421|T191|LLT|10073860|MDR|Paraganglioma|8680/1
C0030421|T191|LLT|10061332|MDR|Paraganglion neoplasm|8680/1
C0030421|T191|PT|10061332|MDR|Paraganglion neoplasm|8680/1
C0030421|T191|LLT|10033792|MDR|Paraganglion neoplasm NOS|8680/1
C0030421|T191|SY|31959|MEDCIN|chemodectomas|8680/1
C0030421|T191|PT|353399|MEDCIN|gangliocytic paraganglioma|8680/1
C0030421|T191|PT|97872|MEDCIN|neoplasm of paraganglia|8680/1
C0030421|T191|SY|97872|MEDCIN|paraganglia neoplasm|8680/1
C0030421|T191|SY|353399|MEDCIN|paraganglioma gangliocytic|8680/1
C0030421|T191|PT|31959|MEDCIN|paragangliomas|8680/1
C0030421|T191|PM|D010235|MSH|Gangliocytic Paraganglioma|8680/1
C0030421|T191|PM|D010235|MSH|Gangliocytic Paragangliomas|8680/1
C0030421|T191|MH|D010235|MSH|Paraganglioma|8680/1
C0030421|T191|ET|D010235|MSH|Paraganglioma, Gangliocytic|8680/1
C0030421|T191|PM|D010235|MSH|Paragangliomas|8680/1
C0030421|T191|ET|D010235|MSH|Paragangliomas 1|8680/1
C0030421|T191|ET|D010235|MSH|Paragangliomas, Familial, 1|8680/1
C0030421|T191|PM|D010235|MSH|Paragangliomas, Gangliocytic|8680/1
C0030421|T191|ET|D010235|MSH|Paragangliomata|8680/1
C0030421|T191|PN|NOCODE|MTH|Paraganglioma|8680/1
C0030421|T191|SY|C3308|NCI|Neoplasm of Paraganglion|8680/1
C0030421|T191|SY|C3308|NCI|Neoplasm of the Paraganglion|8680/1
C0030421|T191|SY|TCGA|NCI|Paraganglioma|8680/1
C0030421|T191|PT|C3308|NCI|Paraganglioma|8680/1
C0030421|T191|SY|C3308|NCI|Paraganglion Neoplasm|8680/1
C0030421|T191|SY|C3308|NCI|Paraganglion Tumor|8680/1
C0030421|T191|SY|C3308|NCI|Paraganglionic Neoplasm|8680/1
C0030421|T191|SY|C3308|NCI|Paraganglionic Tumor|8680/1
C0030421|T191|SY|C3308|NCI|Tumor of Paraganglion|8680/1
C0030421|T191|SY|C3308|NCI|Tumor of the Paraganglion|8680/1
C0030421|T191|DN|C3308|NCI_CTRP|Paraganglioma|8680/1
C0030421|T191|PT|CDR0000390305|NCI_NCI-GLOSS|paraganglioma|8680/1
C0030421|T191|SY|CDR0000639696|PDQ|Neoplasm of Paraganglion|8680/1
C0030421|T191|SY|CDR0000639696|PDQ|Neoplasm of the Paraganglion|8680/1
C0030421|T191|PT|CDR0000639696|PDQ|paraganglioma|8680/1
C0030421|T191|SY|CDR0000639696|PDQ|Paraganglion Neoplasm|8680/1
C0030421|T191|SY|CDR0000639696|PDQ|Paraganglion Tumor|8680/1
C0030421|T191|SY|CDR0000639696|PDQ|Paraganglionic Neoplasm|8680/1
C0030421|T191|SY|CDR0000639696|PDQ|Paraganglionic Tumor|8680/1
C0030421|T191|SY|CDR0000639696|PDQ|Tumor of Paraganglion|8680/1
C0030421|T191|SY|CDR0000639696|PDQ|Tumor of the Paraganglion|8680/1
C0030421|T191|PT|X77oB|RCD|Gangliocytic paraganglioma|8680/1
C0030421|T191|PT|Xa99M|RCD|Paraganglioma|8680/1
C0030421|T191|OP|BBDE.|RCDSY|Gangliocytic paraganglioma|8680/1
C0030421|T191|OP|BBD0.|RCDSY|Paraganglioma NOS|8680/1
C0030421|T191|PT|72787006|SNOMEDCT_US|Gangliocytic paraganglioma|8680/1
C0030421|T191|PT|253029009|SNOMEDCT_US|Gangliocytic paraganglioma|8680/1
C0030421|T191|PT|127027008|SNOMEDCT_US|Neoplasm of paraganglion|8680/1
C0030421|T191|PT|302833002|SNOMEDCT_US|Paraganglioma|8680/1
C0030421|T191|PT|803009|SNOMEDCT_US|Paraganglioma|8680/1
C0030421|T191|IS|803009|SNOMEDCT_US|Paraganglioma, NOS|8680/1
C1533592|T191|LLT|10075444|MDR|Malignant paraganglioma|8680/3
C1533592|T191|LLT|10026665|MDR|Malignant paraganglion neoplasm|8680/3
C1533592|T191|LLT|10033791|MDR|Paraganglion neoplasm malignant|8680/3
C1533592|T191|PT|10033791|MDR|Paraganglion neoplasm malignant|8680/3
C1533592|T191|PT|97873|MEDCIN|malignant neoplasm of paraganglia|8680/3
C1533592|T191|SY|97873|MEDCIN|malignant paraganglia neoplasm|8680/3
C1533592|T191|PT|271490|MEDCIN|malignant paraganglioma|8680/3
C1533592|T191|SY|97873|MEDCIN|malignant tumor of paraganglia|8680/3
C1533592|T191|PN|NOCODE|MTH|Malignant Paraganglionic Neoplasm|8680/3
C1533592|T191|SY|C8559|NCI|Malignant Neoplasm of Paraganglion|8680/3
C1533592|T191|SY|C8559|NCI|Malignant Neoplasm of the Paraganglion|8680/3
C1533592|T191|PT|C8559|NCI|Malignant Paraganglioma|8680/3
C1533592|T191|SY|C8559|NCI|Malignant Paraganglion Neoplasm|8680/3
C1533592|T191|SY|C8559|NCI|Malignant Paraganglion Tumor|8680/3
C1533592|T191|SY|C8559|NCI|Malignant Paraganglionic Neoplasm|8680/3
C1533592|T191|SY|C8559|NCI|Malignant Paraganglionic Tumor|8680/3
C1533592|T191|SY|C8559|NCI|Malignant Tumor of Paraganglion|8680/3
C1533592|T191|SY|C8559|NCI|Malignant Tumor of the Paraganglion|8680/3
C1533592|T191|SY|C8559|NCI|Paraganglion Neoplasm, Malignant|8680/3
C1533592|T191|SY|C8559|NCI_CDISC|Malignant Neoplasm of Paraganglion|8680/3
C1533592|T191|SY|C8559|NCI_CDISC|Malignant Paraganglion Tumor|8680/3
C1533592|T191|PT|C8559|NCI_CDISC|PARAGANGLIOMA, MALIGNANT|8680/3
C1533592|T191|PT|C8559|NCI_CPTAC|Malignant Paraganglioma|8680/3
C1533592|T191|DN|C8559|NCI_CTRP|Malignant Paraganglioma|8680/3
C1533592|T191|PT|CDR0000639698|PDQ|extra-adrenal paraganglioma|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Malignant Neoplasm of Paraganglion|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Malignant Neoplasm of the Paraganglion|8680/3
C1533592|T191|LV|CDR0000639698|PDQ|Malignant Paraganglioma|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Malignant Paraganglion Neoplasm|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Malignant Paraganglion Tumor|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Malignant Paraganglionic Neoplasm|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Malignant Paraganglionic Tumor|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Malignant Tumor of Paraganglion|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Malignant Tumor of the Paraganglion|8680/3
C1533592|T191|SY|CDR0000639698|PDQ|Paraganglion Neoplasm, Malignant|8680/3
C1533592|T191|PT|BBD1.|RCD|Malignant paraganglioma|8680/3
C1533592|T191|SY|9903002|SNOMEDCT_US|Malignant paraganglioma|8680/3
C1533592|T191|PT|9903002|SNOMEDCT_US|Paraganglioma, malignant|8680/3
C0334415|T191|PN|NOCODE|MTH|Sympathetic paraganglioma|8681/1
C0334415|T191|SY|C4216|NCI|Chromaffin Neoplasm|8681/1
C0334415|T191|SY|C4216|NCI|Chromaffin Tumor|8681/1
C0334415|T191|SY|C4216|NCI|Chromaffinoma|8681/1
C0334415|T191|PT|C4216|NCI|Sympathetic Paraganglioma|8681/1
C0334415|T191|SY|C4216|NCI|Sympathetic Paraganglionic Neoplasm|8681/1
C0334415|T191|PT|BBD2.|RCD|Sympathetic paraganglioma|8681/1
C0334415|T191|PT|31794002|SNOMEDCT_US|Sympathetic paraganglioma|8681/1
C0334416|T191|SY|C4217|NCI|Parasympathetic Extra-Adrenal Paraganglioma|8682/1
C0334416|T191|PT|C4217|NCI|Parasympathetic Paraganglioma|8682/1
C0334416|T191|SY|C4217|NCI|Parasympathetic Paraganglionic Neoplasm|8682/1
C0334416|T191|PT|BBD3.|RCD|Parasympathetic paraganglioma|8682/1
C0334416|T191|PT|52205002|SNOMEDCT_US|Parasympathetic paraganglioma|8682/1
C0030421|T191|ET|0000004658|AOD|paraganglioma|8683/0
C0030421|T191|PT|0000009261|CHV|paraganglioma|8683/0
C0030421|T191|SY|0000009261|CHV|paragangliomas|8683/0
C0030421|T191|SY|HP:0002668|HPO|Carotid body tumors|8683/0
C0030421|T191|PT|HP:0002668|HPO|Paraganglioma|8683/0
C0030421|T191|SY|HP:0002668|HPO|Paragangliomas|8683/0
C0030421|T191|PT|MTHU030260|ICPC2ICD10ENG|gangliocytic; paraganglioma, unspecified site|8683/0
C0030421|T191|PT|MTHU057395|ICPC2ICD10ENG|paraganglioma; gangliocytic, unspecified site|8683/0
C0030421|T191|LLT|10073860|MDR|Paraganglioma|8683/0
C0030421|T191|LLT|10061332|MDR|Paraganglion neoplasm|8683/0
C0030421|T191|PT|10061332|MDR|Paraganglion neoplasm|8683/0
C0030421|T191|LLT|10033792|MDR|Paraganglion neoplasm NOS|8683/0
C0030421|T191|SY|31959|MEDCIN|chemodectomas|8683/0
C0030421|T191|PT|353399|MEDCIN|gangliocytic paraganglioma|8683/0
C0030421|T191|PT|97872|MEDCIN|neoplasm of paraganglia|8683/0
C0030421|T191|SY|97872|MEDCIN|paraganglia neoplasm|8683/0
C0030421|T191|SY|353399|MEDCIN|paraganglioma gangliocytic|8683/0
C0030421|T191|PT|31959|MEDCIN|paragangliomas|8683/0
C0030421|T191|PM|D010235|MSH|Gangliocytic Paraganglioma|8683/0
C0030421|T191|PM|D010235|MSH|Gangliocytic Paragangliomas|8683/0
C0030421|T191|MH|D010235|MSH|Paraganglioma|8683/0
C0030421|T191|ET|D010235|MSH|Paraganglioma, Gangliocytic|8683/0
C0030421|T191|PM|D010235|MSH|Paragangliomas|8683/0
C0030421|T191|ET|D010235|MSH|Paragangliomas 1|8683/0
C0030421|T191|ET|D010235|MSH|Paragangliomas, Familial, 1|8683/0
C0030421|T191|PM|D010235|MSH|Paragangliomas, Gangliocytic|8683/0
C0030421|T191|ET|D010235|MSH|Paragangliomata|8683/0
C0030421|T191|PN|NOCODE|MTH|Paraganglioma|8683/0
C1334232|T191|SY|C5325|NCI|Gangliocytic Intestinal Paraganglioma|8683/0
C1334232|T191|SY|C5325|NCI|Gangliocytic Paraganglioma of Intestine|8683/0
C1334232|T191|SY|C5325|NCI|Gangliocytic Paraganglioma of the Intestine|8683/0
C1334232|T191|PT|C5325|NCI|Intestinal Gangliocytic Paraganglioma|8683/0
C0030421|T191|SY|C3308|NCI|Neoplasm of Paraganglion|8683/0
C0030421|T191|SY|C3308|NCI|Neoplasm of the Paraganglion|8683/0
C0030421|T191|PT|C3308|NCI|Paraganglioma|8683/0
C0030421|T191|SY|TCGA|NCI|Paraganglioma|8683/0
C0030421|T191|SY|C3308|NCI|Paraganglion Neoplasm|8683/0
C0030421|T191|SY|C3308|NCI|Paraganglion Tumor|8683/0
C0030421|T191|SY|C3308|NCI|Paraganglionic Neoplasm|8683/0
C0030421|T191|SY|C3308|NCI|Paraganglionic Tumor|8683/0
C0030421|T191|SY|C3308|NCI|Tumor of Paraganglion|8683/0
C0030421|T191|SY|C3308|NCI|Tumor of the Paraganglion|8683/0
C0030421|T191|DN|C3308|NCI_CTRP|Paraganglioma|8683/0
C0030421|T191|PT|CDR0000390305|NCI_NCI-GLOSS|paraganglioma|8683/0
C0030421|T191|SY|CDR0000639696|PDQ|Neoplasm of Paraganglion|8683/0
C0030421|T191|SY|CDR0000639696|PDQ|Neoplasm of the Paraganglion|8683/0
C0030421|T191|PT|CDR0000639696|PDQ|paraganglioma|8683/0
C0030421|T191|SY|CDR0000639696|PDQ|Paraganglion Neoplasm|8683/0
C0030421|T191|SY|CDR0000639696|PDQ|Paraganglion Tumor|8683/0
C0030421|T191|SY|CDR0000639696|PDQ|Paraganglionic Neoplasm|8683/0
C0030421|T191|SY|CDR0000639696|PDQ|Paraganglionic Tumor|8683/0
C0030421|T191|SY|CDR0000639696|PDQ|Tumor of Paraganglion|8683/0
C0030421|T191|SY|CDR0000639696|PDQ|Tumor of the Paraganglion|8683/0
C0030421|T191|PT|X77oB|RCD|Gangliocytic paraganglioma|8683/0
C0030421|T191|PT|Xa99M|RCD|Paraganglioma|8683/0
C0030421|T191|OP|BBDE.|RCDSY|Gangliocytic paraganglioma|8683/0
C0030421|T191|OP|BBD0.|RCDSY|Paraganglioma NOS|8683/0
C0030421|T191|PT|72787006|SNOMEDCT_US|Gangliocytic paraganglioma|8683/0
C0030421|T191|PT|253029009|SNOMEDCT_US|Gangliocytic paraganglioma|8683/0
C0030421|T191|PT|127027008|SNOMEDCT_US|Neoplasm of paraganglion|8683/0
C0030421|T191|PT|302833002|SNOMEDCT_US|Paraganglioma|8683/0
C0030421|T191|PT|803009|SNOMEDCT_US|Paraganglioma|8683/0
C0030421|T191|IS|803009|SNOMEDCT_US|Paraganglioma, NOS|8683/0
C0017671|T191|PT|0050182|CCPSS|GLOMUS JUGULARE TUMOR|8690/1
C0017671|T191|PT|0000005544|CHV|glomus jugulare tumor|8690/1
C0017671|T191|SY|0000005544|CHV|glomus jugulare tumors|8690/1
C0017671|T191|SY|0000005544|CHV|jugular paragangliomas|8690/1
C0017671|T191|DI|U000730|DXP|GLOMUS JUGULARE TUMOR|8690/1
C0017671|T191|PT|HP:0003001|HPO|Glomus jugular tumor|8690/1
C0017671|T191|SY|HP:0003001|HPO|Glomus jugulare tumor|8690/1
C0017671|T191|SY|HP:0003001|HPO|Glomus jugulare tumors|8690/1
C0017671|T191|PT|MTHU077067|ICPC2ICD10ENG|tumor; glomus jugulare|8690/1
C0017671|T191|PT|sh85055321|LCH_NW|Glomus jugulare--Tumors|8690/1
C0017671|T191|LLT|10056573|MDR|Glomus jugulare tumor|8690/1
C0017671|T191|MTH_PT|10056563|MDR|Glomus jugulare tumor|8690/1
C0017671|T191|LLT|10056563|MDR|Glomus jugulare tumour|8690/1
C0017671|T191|PT|10056563|MDR|Glomus jugulare tumour|8690/1
C0017671|T191|PT|31751|MEDCIN|neoplasm of glomus jugulare|8690/1
C0017671|T191|MH|D005925|MSH|Glomus Jugulare Tumor|8690/1
C0017671|T191|ET|D005925|MSH|Glomus Jugulare Tumors|8690/1
C0017671|T191|PM|D005925|MSH|Jugulare Tumor, Glomus|8690/1
C0017671|T191|PM|D005925|MSH|Jugulare Tumors, Glomus|8690/1
C0017671|T191|PM|D005925|MSH|Tumor, Glomus Jugulare|8690/1
C0017671|T191|PM|D005925|MSH|Tumors, Glomus Jugulare|8690/1
C0017671|T191|PN|NOCODE|MTH|Glomus Jugulare Tumor|8690/1
C0017671|T191|SY|C3061|NCI|Glomus Jugulare Neoplasm|8690/1
C0017671|T191|SY|C3061|NCI|Glomus Jugulare Tumor|8690/1
C0017671|T191|SY|C3061|NCI|Jugular Paraganglioma|8690/1
C0017671|T191|PT|C3061|NCI|Jugulotympanic Paraganglioma|8690/1
C0017671|T191|SY|C3061|NCI|Neoplasm of Glomus Jugulare|8690/1
C0017671|T191|SY|C3061|NCI|Neoplasm of the Glomus Jugulare|8690/1
C0017671|T191|SY|C3061|NCI|Tumor of Glomus Jugulare|8690/1
C0017671|T191|SY|C3061|NCI|Tumor of the Glomus Jugulare|8690/1
C0017671|T191|SY|BBD4.|RCD|Glomus jugulare tumour|8690/1
C0017671|T191|SY|BBD4.|RCD|Jugular paraganglioma|8690/1
C0017671|T191|SY|BBD4.|RCDAE|Glomus jugulare tumor|8690/1
C0017671|T191|PT|32037004|SNOMEDCT_US|Glomus jugulare tumor|8690/1
C0017671|T191|PTGB|32037004|SNOMEDCT_US|Glomus jugulare tumour|8690/1
C0017671|T191|SY|32037004|SNOMEDCT_US|Jugular paraganglioma|8690/1
C0017671|T191|SY|32037004|SNOMEDCT_US|Jugulotympanic paraganglioma|8690/1
C0017671|T191|PT|127030001|SNOMEDCT_US|Neoplasm of glomus jugulare|8690/1
C0334417|T191|PT|MTHU057396|ICPC2ICD10ENG|paraganglioma; aortic body|8691/1
C0334417|T191|PT|MTHU077065|ICPC2ICD10ENG|tumor; aortic body|8691/1
C0334417|T191|PT|97870|MEDCIN|neoplasm of aortic body|8691/1
C0334417|T191|SY|C4218|NCI|Aortic Body Neoplasm|8691/1
C0334417|T191|SY|C4218|NCI|Aortic Body Paraganglioma|8691/1
C0334417|T191|SY|C4218|NCI|Aortic Body Tumor|8691/1
C0334417|T191|PT|C4218|NCI|Aorticopulmonary Paraganglioma|8691/1
C0334417|T191|SY|C4218|NCI|Neoplasm of Aortic Body|8691/1
C0334417|T191|SY|C4218|NCI|Neoplasm of the Aortic Body|8691/1
C0334417|T191|SY|C4218|NCI|Paraganglioma of Aortic Body|8691/1
C0334417|T191|SY|C4218|NCI|Paraganglioma of the Aortic Body|8691/1
C0334417|T191|SY|C4218|NCI|Tumor of Aortic Body|8691/1
C0334417|T191|SY|C4218|NCI|Tumor of the Aortic Body|8691/1
C0334417|T191|SY|BBD5.|RCD|Aortic body paraganglioma|8691/1
C0334417|T191|SY|BBD5.|RCD|Aortic body tumour|8691/1
C0334417|T191|SY|BBD5.|RCDAE|Aortic body tumor|8691/1
C0334417|T191|SY|53320004|SNOMEDCT_US|Aortic body paraganglioma|8691/1
C0334417|T191|PT|53320004|SNOMEDCT_US|Aortic body tumor|8691/1
C0334417|T191|PTGB|53320004|SNOMEDCT_US|Aortic body tumour|8691/1
C0334417|T191|SY|53320004|SNOMEDCT_US|Aorticopulmonary paraganglioma|8691/1
C0334417|T191|PT|127029006|SNOMEDCT_US|Neoplasm of aortic body|8691/1
C0007279|T191|SY|0000002480|CHV|body carotid tumours|8692/1
C0007279|T191|PT|0000002480|CHV|carotid body tumor|8692/1
C0007279|T191|SY|0000002480|CHV|carotid body tumors|8692/1
C0007279|T191|SY|0000002480|CHV|carotid body tumour|8692/1
C0007279|T191|SY|0000002480|CHV|paraganglioma carotid body|8692/1
C0007279|T191|DI|U000300|DXP|CAROTID BODY, TUMOR|8692/1
C0007279|T191|PT|HP:0030074|HPO|Chemodectoma|8692/1
C0007279|T191|SY|HP:0030074|HPO|Chemodectomas|8692/1
C0007279|T191|PT|MTHU057398|ICPC2ICD10ENG|paraganglioma; carotid body|8692/1
C0007279|T191|PT|MTHU077066|ICPC2ICD10ENG|tumor; carotid body|8692/1
C0007279|T191|PT|sh85020417|LCH_NW|Carotid body--Tumors|8692/1
C0007279|T191|LLT|10007689|MDR|Carotid body tumor|8692/1
C0007279|T191|MTH_PT|10007690|MDR|Carotid body tumor|8692/1
C0007279|T191|LLT|10007690|MDR|Carotid body tumour|8692/1
C0007279|T191|PT|10007690|MDR|Carotid body tumour|8692/1
C0007279|T191|LLT|10075392|MDR|Glomus caroticum tumor|8692/1
C0007279|T191|LLT|10075388|MDR|Glomus caroticum tumour|8692/1
C0007279|T191|PT|31752|MEDCIN|carotid body tumor|8692/1
C0007279|T191|PM|D002345|MSH|Carotid Body Paraganglioma|8692/1
C0007279|T191|PM|D002345|MSH|Carotid Body Paragangliomas|8692/1
C0007279|T191|MH|D002345|MSH|Carotid Body Tumor|8692/1
C0007279|T191|ET|D002345|MSH|Carotid Body Tumors|8692/1
C0007279|T191|ET|D002345|MSH|Paraganglioma, Carotid Body|8692/1
C0007279|T191|PM|D002345|MSH|Paragangliomas, Carotid Body|8692/1
C0007279|T191|PM|D002345|MSH|Tumor, Carotid Body|8692/1
C0007279|T191|PM|D002345|MSH|Tumors, Carotid Body|8692/1
C0007279|T191|PN|NOCODE|MTH|Carotid Body Paraganglioma|8692/1
C0007279|T191|SY|C2932|NCI|Carotid Body Chemodectoma|8692/1
C0007279|T191|PT|C2932|NCI|Carotid Body Paraganglioma|8692/1
C0007279|T191|SY|C2932|NCI|Carotid Body Tumor|8692/1
C0007279|T191|SY|C2932|NCI|Chemodectoma|8692/1
C0007279|T191|SY|C2932|NCI|Paraganglioma of Carotid Body|8692/1
C0007279|T191|SY|C2932|NCI|Paraganglioma of the Carotid Body|8692/1
C0007279|T191|SY|C2932|NCI|Tumor of Carotid Body|8692/1
C0007279|T191|SY|C2932|NCI|Tumor of the Carotid Body|8692/1
C0007279|T191|SY|BBD6.|RCD|Carotid body paraganglioma|8692/1
C0007279|T191|SY|BBD6.|RCD|Carotid body tumour|8692/1
C0007279|T191|SY|BBD6.|RCDAE|Carotid body tumor|8692/1
C0007279|T191|SY|30699005|SNOMEDCT_US|Carotid body paraganglioma|8692/1
C0007279|T191|PT|30699005|SNOMEDCT_US|Carotid body tumor|8692/1
C0007279|T191|PTGB|30699005|SNOMEDCT_US|Carotid body tumour|8692/1
C0007279|T191|PT|127028003|SNOMEDCT_US|Neoplasm of carotid body|8692/1
C0030422|T191|PT|0000009262|CHV|chemodectoma|8693/1
C0030422|T191|SY|NOCODE|DXP|CHEMODECTOMA|8693/1
C0030422|T191|SY|NOCODE|DXP|PARAGANGLIOMA, NONCHROMAFFIN|8693/1
C0030422|T191|PT|sh85092239|LCH_NW|Nonchromaffin paraganglioma|8693/1
C0030422|T191|LLT|10051227|MDR|Chemodectoma|8693/1
C0030422|T191|PT|10051227|MDR|Chemodectoma|8693/1
C0030422|T191|PT|351586|MEDCIN|extra-adrenal paraganglioma|8693/1
C0030422|T191|SY|351586|MEDCIN|neoplasm of paraganglioma extra-adrenal|8693/1
C0030422|T191|ET|D010236|MSH|Chemodectoma|8693/1
C0030422|T191|ET|D010236|MSH|Chemodectomas|8693/1
C0030422|T191|PM|D010236|MSH|Extra-Adrenal Paraganglioma|8693/1
C0030422|T191|PM|D010236|MSH|Extra-Adrenal Paragangliomas|8693/1
C0030422|T191|PM|D010236|MSH|Non-Chromaffin Paraganglioma|8693/1
C0030422|T191|PM|D010236|MSH|Non-Chromaffin Paragangliomas|8693/1
C0030422|T191|PM|D010236|MSH|Nonchromaffin Paraganglioma|8693/1
C0030422|T191|PM|D010236|MSH|Nonchromaffin Paragangliomas|8693/1
C0030422|T191|PM|D010236|MSH|Paraganglioma, Extra Adrenal|8693/1
C0030422|T191|MH|D010236|MSH|Paraganglioma, Extra-Adrenal|8693/1
C0030422|T191|PM|D010236|MSH|Paraganglioma, Non Chromaffin|8693/1
C0030422|T191|ET|D010236|MSH|Paraganglioma, Non-Chromaffin|8693/1
C0030422|T191|ET|D010236|MSH|Paraganglioma, Nonchromaffin|8693/1
C0030422|T191|PM|D010236|MSH|Paragangliomas, Extra-Adrenal|8693/1
C0030422|T191|ET|D010236|MSH|Paragangliomas, Familial Nonchromaffin, 1|8693/1
C0030422|T191|PM|D010236|MSH|Paragangliomas, Non-Chromaffin|8693/1
C0030422|T191|PM|D010236|MSH|Paragangliomas, Nonchromaffin|8693/1
C0030422|T191|PN|NOCODE|MTH|Extra-Adrenal Paraganglioma|8693/1
C0030422|T191|PT|C3309|NCI|Extra-Adrenal Paraganglioma|8693/1
C0030422|T191|SY|C3309|NCI|Extra-Adrenal Paraganglionic Neoplasm|8693/1
C0030422|T191|SY|C3309|NCI|Extraadrenal Paraganglioma|8693/1
C0030422|T191|DN|C3309|NCI_CTRP|Extra-Adrenal Paraganglioma|8693/1
C0030422|T191|SY|Xa99O|RCD|Chemodectoma|8693/1
C0030422|T191|PT|Xa99O|RCD|Extra-adrenal paraganglioma|8693/1
C0030422|T191|SY|Xa99O|RCD|Non-chromaffin paraganglioma|8693/1
C0030422|T191|SY|Xa99O|RCD|Nonchromaffin paraganglioma|8693/1
C0030422|T191|AB|XE1wW|RCDSY|Extra-adrenal paragangl.NOS|8693/1
C0030422|T191|PT|XE1wW|RCDSY|Extra-adrenal paraganglioma, NOS|8693/1
C0030422|T191|SY|51747000|SNOMEDCT_US|Chemodectoma|8693/1
C0030422|T191|SY|302834008|SNOMEDCT_US|Chemodectoma|8693/1
C0030422|T191|PT|51747000|SNOMEDCT_US|Extra-adrenal paraganglioma|8693/1
C0030422|T191|PT|302834008|SNOMEDCT_US|Extra-adrenal paraganglioma|8693/1
C0030422|T191|IS|51747000|SNOMEDCT_US|Extra-adrenal paraganglioma, NOS|8693/1
C0030422|T191|SY|302834008|SNOMEDCT_US|Non-chromaffin paraganglioma|8693/1
C0030422|T191|SY|51747000|SNOMEDCT_US|Nonchromaffin paraganglioma|8693/1
C0030422|T191|IS|51747000|SNOMEDCT_US|Nonchromaffin paraganglioma, NOS|8693/1
C0334418|T191|PT|271491|MEDCIN|malignant extra-adrenal paraganglioma|8693/3
C4763506|T191|PT|C157246|NCI|Composite Paraganglioma|8693/3
C0334418|T191|PT|C4219|NCI|Malignant Extra-Adrenal Paraganglioma|8693/3
C0334418|T191|AB|BBD8.|RCD|Mal non-chromaf paraganglioma|8693/3
C0334418|T191|AB|BBD8.|RCD|Malig extra-adr paraganglioma|8693/3
C0334418|T191|AB|BBD8.|RCD|Malig nonchromaf paraganglioma|8693/3
C0334418|T191|PT|BBD8.|RCD|Malignant extra-adrenal paraganglioma|8693/3
C0334418|T191|SY|BBD8.|RCD|Malignant non-chromaffin paraganglioma|8693/3
C0334418|T191|SY|BBD8.|RCD|Malignant nonchromaffin paraganglioma|8693/3
C4763506|T191|PT|817953005|SNOMEDCT_US|Composite paraganglioma|8693/3
C0334418|T191|PT|32512003|SNOMEDCT_US|Extra-adrenal paraganglioma, malignant|8693/3
C0334418|T191|SY|32512003|SNOMEDCT_US|Malignant extra-adrenal paraganglioma|8693/3
C0334418|T191|SY|32512003|SNOMEDCT_US|Malignant non-chromaffin paraganglioma|8693/3
C0334418|T191|SY|32512003|SNOMEDCT_US|Nonchromaffin paraganglioma, malignant|8693/3
C4551683|T191|ET|0000004641|AOD|pheochromocytoma|8700/0
C4551683|T191|SY|0000009623|CHV|chromaffin tumor|8700/0
C4551683|T191|SY|0000009623|CHV|phaeochromocytoma|8700/0
C4551683|T191|PT|0000009623|CHV|pheochromocytoma|8700/0
C4551683|T191|SY|0000009623|CHV|pheochromocytoma syndrome|8700/0
C4551683|T191|SY|0000009623|CHV|pheochromocytomas|8700/0
C4551683|T191|ET|2012-7663|CSP|chromaffinoma|8700/0
C4551683|T191|PT|2012-7663|CSP|pheochromocytoma|8700/0
C4551683|T191|SY|NOCODE|DXP|CHROMAFFINOMA, MEDULLARY|8700/0
C4551683|T191|SY|NOCODE|DXP|PARAGANGLIOMA, MEDULLARY|8700/0
C4551683|T191|PT|HP:0006748|HPO|Adrenal pheochromocytoma|8700/0
C4551683|T191|SY|HP:0006748|HPO|Pheochromocytoma, adrenal|8700/0
C4551683|T191|SY|HP:0006748|HPO|Pheochromocytomas, adrenal|8700/0
C4551683|T191|LLT|10034800|MDR|Phaeochromocytoma|8700/0
C4551683|T191|PT|10034800|MDR|Phaeochromocytoma|8700/0
C4551683|T191|LLT|10034876|MDR|Pheochromocytoma|8700/0
C4551683|T191|MTH_PT|10034800|MDR|Pheochromocytoma|8700/0
C4551683|T191|SY|351578|MEDCIN|adrenal neoplasm of uncertain behavior pheochromocytoma|8700/0
C4551683|T191|PT|351578|MEDCIN|pheochromocytoma|8700/0
C4551683|T191|PN|NOCODE|MTH|Adrenal Gland Pheochromocytoma|8700/0
C4551683|T191|SY|C3326|NCI|Adrenal Gland Chromaffin Paraganglioma|8700/0
C4551683|T191|SY|C3326|NCI|Adrenal Gland Chromaffinoma|8700/0
C4551683|T191|SY|C3326|NCI|Adrenal Gland Paraganglioma|8700/0
C4551683|T191|PT|C3326|NCI|Adrenal Gland Pheochromocytoma|8700/0
C4551683|T191|SY|TCGA|NCI|Adrenal Gland Pheochromocytoma|8700/0
C4551683|T191|SY|C3326|NCI|Adrenal Medullary Paraganglioma|8700/0
C4551683|T191|SY|C3326|NCI|Adrenal Medullary Pheochromocytoma|8700/0
C4551683|T191|SY|C3326|NCI|Adrenal Pheochromocytoma|8700/0
C4551683|T191|SY|C3326|NCI|Chromaffin Paraganglioma of the Adrenal Gland|8700/0
C4551683|T191|SY|C3326|NCI|Intraadrenal Paraganglioma|8700/0
C4551683|T191|AB|C3326|NCI|PCC|8700/0
C4551683|T191|SY|C3326|NCI|Pheochromocytoma|8700/0
C4551683|T191|DN|C3326|NCI_CTRP|Pheochromocytoma|8700/0
C4551683|T191|PT|CDR0000322877|NCI_NCI-GLOSS|pheochromocytoma|8700/0
C0474822|T191|PT|X77oF|RCD|Benign phaeochromocytoma|8700/0
C0474822|T191|AB|XaBA3|RCD|Benign phaeochromocytoma morph|8700/0
C0474822|T191|PT|XaBA3|RCD|Benign phaeochromocytoma morphology|8700/0
C4551683|T191|SY|Xa99P|RCD|Chromaffin paraganglioma|8700/0
C4551683|T191|SY|Xa99P|RCD|Chromaffin tumour|8700/0
C4551683|T191|SY|Xa99P|RCD|Chromaffinoma|8700/0
C4551683|T191|PT|Xa99P|RCD|Phaeochromocytoma|8700/0
C0474822|T191|PT|X77oF|RCDAE|Benign pheochromocytoma|8700/0
C0474822|T191|AB|XaBA3|RCDAE|Benign pheochromocytoma morph|8700/0
C0474822|T191|PT|XaBA3|RCDAE|Benign pheochromocytoma morphology|8700/0
C4551683|T191|SY|Xa99P|RCDAE|Chromaffin tumor|8700/0
C4551683|T191|PT|Xa99P|RCDAE|Pheochromocytoma|8700/0
C4551683|T191|PT|BBD9.|RCDSA|Pheochromocytoma NOS|8700/0
C4551683|T191|PT|BBD9.|RCDSY|Phaeochromocytoma NOS|8700/0
C4551683|T191|SY|302835009|SNOMEDCT_US|Adrenal medullary paraganglioma|8700/0
C4551683|T191|SY|85583005|SNOMEDCT_US|Adrenal medullary paraganglioma|8700/0
C0474822|T191|OAP|189177006|SNOMEDCT_US|Benign phaeochromocytoma|8700/0
C0474822|T191|OF|189177006|SNOMEDCT_US|Benign phaeochromocytoma|8700/0
C0474822|T191|PTGB|307575002|SNOMEDCT_US|Benign phaeochromocytoma|8700/0
C0474822|T191|PTGB|253032007|SNOMEDCT_US|Benign phaeochromocytoma|8700/0
C0474822|T191|SYGB|307575002|SNOMEDCT_US|Benign phaeochromocytoma morphology|8700/0
C0474822|T191|OAP|189177006|SNOMEDCT_US|Benign pheochromocytoma|8700/0
C0474822|T191|PT|307575002|SNOMEDCT_US|Benign pheochromocytoma|8700/0
C0474822|T191|PT|253032007|SNOMEDCT_US|Benign pheochromocytoma|8700/0
C0474822|T191|SY|307575002|SNOMEDCT_US|Benign pheochromocytoma morphology|8700/0
C4551683|T191|OAP|399258001|SNOMEDCT_US|Chromaffin cell neoplasm|8700/0
C4551683|T191|SY|85583005|SNOMEDCT_US|Chromaffin cell neoplasm|8700/0
C4551683|T191|SY|85583005|SNOMEDCT_US|Chromaffin paraganglioma|8700/0
C4551683|T191|SY|302835009|SNOMEDCT_US|Chromaffin paraganglioma|8700/0
C4551683|T191|SY|85583005|SNOMEDCT_US|Chromaffin tumor|8700/0
C4551683|T191|SY|302835009|SNOMEDCT_US|Chromaffin tumor|8700/0
C4551683|T191|SYGB|85583005|SNOMEDCT_US|Chromaffin tumour|8700/0
C4551683|T191|SYGB|302835009|SNOMEDCT_US|Chromaffin tumour|8700/0
C4551683|T191|SY|85583005|SNOMEDCT_US|Chromaffinoma|8700/0
C4551683|T191|SY|302835009|SNOMEDCT_US|Chromaffinoma|8700/0
C4551683|T191|PTGB|85583005|SNOMEDCT_US|Phaeochromocytoma|8700/0
C4551683|T191|PTGB|302835009|SNOMEDCT_US|Phaeochromocytoma|8700/0
C4551683|T191|IS|85583005|SNOMEDCT_US|Phaeochromocytoma, NOS|8700/0
C4551683|T191|PT|302835009|SNOMEDCT_US|Pheochromocytoma|8700/0
C4551683|T191|PT|85583005|SNOMEDCT_US|Pheochromocytoma|8700/0
C4551683|T191|IS|85583005|SNOMEDCT_US|Pheochromocytoma, NOS|8700/0
C0334419|T191|PT|MTHU047281|ICPC2ICD10ENG|malignant; pheochromocytoma, unspecified site|8700/3
C0334419|T191|PT|MTHU028073|ICPC2ICD10ENG|pheochromocytoma; malignant, unspecified site|8700/3
C0334419|T191|PT|10051710|MDR|Phaeochromocytoma malignant|8700/3
C0334419|T191|LLT|10051710|MDR|Phaeochromocytoma malignant|8700/3
C0334419|T191|MTH_LLT|10051710|MDR|Pheochromocytoma malignant|8700/3
C0334419|T191|MTH_PT|10051710|MDR|Pheochromocytoma malignant|8700/3
C0334419|T191|PT|236340|MEDCIN|malignant paraganglioma of adrenal gland|8700/3
C0334419|T191|PT|34858|MEDCIN|malignant pheochromocytoma|8700/3
C0334419|T191|PT|236342|MEDCIN|malignant pheochromocytoma of adrenal gland|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Adrenal Gland Chromaffin Neoplasm|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Adrenal Gland Chromaffin Paraganglioma|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Adrenal Gland Chromaffin Tumor|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Adrenal Gland Chromaffinoma|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Adrenal Gland Paraganglioma|8700/3
C0334419|T191|PT|C4220|NCI|Malignant Adrenal Gland Pheochromocytoma|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Adrenal Medullary Paraganglioma|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Adrenal Medullary Pheochromocytoma|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Adrenal Pheochromocytoma|8700/3
C0334419|T191|SY|C4220|NCI|Malignant Pheochromocytoma|8700/3
C0334419|T191|SY|C4220|NCI|Pheochromoblastoma|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Adrenal Gland Chromaffin Neoplasm|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Adrenal Gland Chromaffin Paraganglioma|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Adrenal Gland Chromaffin Tumor|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Adrenal Gland Chromaffinoma|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Adrenal Gland Paraganglioma|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Adrenal Medullary Paraganglioma|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Adrenal Medullary Pheochromocytoma|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Adrenal Pheochromocytoma|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Malignant Pheochromocytoma|8700/3
C0334419|T191|SY|C4220|NCI_CDISC|Pheochromoblastoma|8700/3
C0334419|T191|PT|C4220|NCI_CDISC|PHEOCHROMOCYTOMA, MALIGNANT|8700/3
C0334419|T191|PT|BBDA.|RCD|Malignant phaeochromocytoma|8700/3
C0334419|T191|SY|BBDA.|RCD|Phaeochromoblastoma|8700/3
C0334419|T191|PT|BBDA.|RCDAE|Malignant pheochromocytoma|8700/3
C0334419|T191|SY|BBDA.|RCDAE|Pheochromoblastoma|8700/3
C0334419|T191|SY|29370006|SNOMEDCT_US|Adrenal medullary paraganglioma, malignant|8700/3
C5231203|T191|PTGB|817952000|SNOMEDCT_US|Composite phaeochromocytoma|8700/3
C5231203|T191|PT|817952000|SNOMEDCT_US|Composite pheochromocytoma|8700/3
C0334419|T191|PTGB|21851000119103|SNOMEDCT_US|Malignant phaeochromocytoma|8700/3
C0334419|T191|PTGB|29370006|SNOMEDCT_US|Malignant phaeochromocytoma|8700/3
C0334419|T191|PT|29370006|SNOMEDCT_US|Malignant pheochromocytoma|8700/3
C0334419|T191|PT|21851000119103|SNOMEDCT_US|Malignant pheochromocytoma|8700/3
C0334419|T191|SYGB|29370006|SNOMEDCT_US|Phaeochromoblastoma|8700/3
C0334419|T191|SYGB|29370006|SNOMEDCT_US|Phaeochromocytoma, malignant|8700/3
C0334419|T191|SY|29370006|SNOMEDCT_US|Pheochromoblastoma|8700/3
C0334419|T191|SY|29370006|SNOMEDCT_US|Pheochromocytoma, malignant|8700/3
C1266111|T191|PT|MTHU032305|ICPC2ICD10ENG|glomoid; sarcoma|8710/3
C1266111|T191|PT|MTHU065899|ICPC2ICD10ENG|sarcoma; glomoid|8710/3
C1266111|T191|PT|271524|MEDCIN|glomangiosarcoma|8710/3
C1266111|T191|SY|C4221|NCI|Glomangiosarcoma|8710/3
C1266111|T191|SY|C4221|NCI|Malignant Glomus Neoplasm|8710/3
C1266111|T191|PT|C4221|NCI|Malignant Glomus Tumor|8710/3
C1266111|T191|PT|BBDB.|RCD|Glomangiosarcoma|8710/3
C1266111|T191|SY|BBDB.|RCD|Glomoid sarcoma|8710/3
C1266111|T191|PT|13875003|SNOMEDCT_US|Glomangiosarcoma|8710/3
C1266111|T191|SY|13875003|SNOMEDCT_US|Glomoid sarcoma|8710/3
C1266111|T191|PT|128908003|SNOMEDCT_US|Glomus tumor, malignant|8710/3
C1266111|T191|PTGB|128908003|SNOMEDCT_US|Glomus tumour, malignant|8710/3
C0017653|T191|PT|0000005534|CHV|glomus tumor|8711/0
C0017653|T191|SY|0000005534|CHV|glomus tumors|8711/0
C0017653|T191|SY|0000005534|CHV|glomus tumour|8711/0
C0017653|T191|SY|0000005534|CHV|tumor glomus|8711/0
C0017653|T191|PT|NOCODE|COSTAR|Glomus Tumor|8711/0
C0017653|T191|LLT|10018380|MDR|Glomus tumor|8711/0
C0017653|T191|MTH_PT|10018381|MDR|Glomus tumor|8711/0
C0017653|T191|LLT|10018381|MDR|Glomus tumour|8711/0
C0017653|T191|PT|10018381|MDR|Glomus tumour|8711/0
C0017653|T191|MH|D005918|MSH|Glomus Tumor|8711/0
C0017653|T191|PM|D005918|MSH|Glomus Tumors|8711/0
C0017653|T191|PM|D005918|MSH|Tumor, Glomus|8711/0
C0017653|T191|PM|D005918|MSH|Tumors, Glomus|8711/0
C0017653|T191|PN|NOCODE|MTH|Glomus Tumor|8711/0
C0017653|T191|SY|C3060|NCI|Glomus Neoplasm|8711/0
C0017653|T191|PT|C3060|NCI|Glomus Tumor|8711/0
C0017653|T191|PT|BBDC.|RCD|Glomus tumour|8711/0
C0017653|T191|PT|BBDC.|RCDAE|Glomus tumor|8711/0
C0017653|T191|PT|403969002|SNOMEDCT_US|Glomus tumor|8711/0
C0017653|T191|PT|10438002|SNOMEDCT_US|Glomus tumor|8711/0
C0017653|T191|OAS|189193002|SNOMEDCT_US|Glomus tumor|8711/0
C0017653|T191|PTGB|403969002|SNOMEDCT_US|Glomus tumour|8711/0
C0017653|T191|PTGB|10438002|SNOMEDCT_US|Glomus tumour|8711/0
C0017653|T191|OAP|393567008|SNOMEDCT_US|Glomus tumour|8711/0
C0017653|T191|OAS|189193002|SNOMEDCT_US|Glomus tumour|8711/0
C0017653|T191|OF|393567008|SNOMEDCT_US|Glomus tumour|8711/0
C1333824|T191|PT|C27496|NCI|Glomangiomatosis|8711/1
C1333824|T191|PT|703603008|SNOMEDCT_US|Glomangiomatosis|8711/1
C1266111|T191|PT|MTHU032305|ICPC2ICD10ENG|glomoid; sarcoma|8711/3
C1266111|T191|PT|MTHU065899|ICPC2ICD10ENG|sarcoma; glomoid|8711/3
C1266111|T191|PT|271524|MEDCIN|glomangiosarcoma|8711/3
C1266111|T191|SY|C4221|NCI|Glomangiosarcoma|8711/3
C1266111|T191|SY|C4221|NCI|Malignant Glomus Neoplasm|8711/3
C1266111|T191|PT|C4221|NCI|Malignant Glomus Tumor|8711/3
C1266111|T191|PT|BBDB.|RCD|Glomangiosarcoma|8711/3
C1266111|T191|SY|BBDB.|RCD|Glomoid sarcoma|8711/3
C1266111|T191|PT|13875003|SNOMEDCT_US|Glomangiosarcoma|8711/3
C1266111|T191|SY|13875003|SNOMEDCT_US|Glomoid sarcoma|8711/3
C1266111|T191|PT|128908003|SNOMEDCT_US|Glomus tumor, malignant|8711/3
C1266111|T191|PTGB|128908003|SNOMEDCT_US|Glomus tumour, malignant|8711/3
C0334421|T191|PT|0000029974|CHV|glomangioma|8712/0
C0334421|T191|SY|0000029974|CHV|glomangiomas|8712/0
C0334421|T191|ET|2007-0683|CSP|glomangioma|8712/0
C0334421|T191|PT|MTHU032181|ICPC2ICD10ENG|glomangioma|8712/0
C0334421|T191|PEP|D005918|MSH|Glomangioma|8712/0
C0334421|T191|PM|D005918|MSH|Glomangiomas|8712/0
C0334421|T191|PN|NOCODE|MTH|Glomangioma|8712/0
C0334421|T191|PT|C4222|NCI|Glomangioma|8712/0
C0334421|T191|PT|BBDD.|RCD|Glomangioma|8712/0
C0334421|T191|PT|7429002|SNOMEDCT_US|Glomangioma|8712/0
C0334422|T191|PT|MTHU032180|ICPC2ICD10ENG|glomangiomyoma|8713/0
C0334422|T191|PT|C4223|NCI|Glomangiomyoma|8713/0
C0334422|T191|PT|X77oG|RCD|Glomangiomyoma|8713/0
C0334422|T191|OAP|189745002|SNOMEDCT_US|Glomangiomyoma|8713/0
C0334422|T191|OF|189745002|SNOMEDCT_US|Glomangiomyoma|8713/0
C0334422|T191|PT|34550005|SNOMEDCT_US|Glomangiomyoma|8713/0
C1302808|T191|MH|D000077777|MSH|Myopericytoma|8713/1
C1302808|T191|PM|D000077777|MSH|Myopericytomas|8713/1
C1302808|T191|PN|NOCODE|MTH|Myopericytoma|8713/1
C1302808|T191|OP|C50401|NCI|Hemangiopericytoma|8713/1
C1302808|T191|PT|C50401|NCI|Myopericytoma|8713/1
C1302808|T191|OP|C50401|NCI|Solitary Myofibroma|8713/1
C1302808|T191|PT|400065005|SNOMEDCT_US|Myopericytoma|8713/1
C3839685|T191|PT|C121791|NCI|Benign PEComa|8714/0
C3839685|T191|SY|C121791|NCI|Benign PEComa, NOS|8714/0
C3839685|T191|SY|C121791|NCI|Benign PEComa, Not Otherwise Specified|8714/0
C3839685|T191|SY|C121791|NCI|Typical PEComa|8714/0
C3839685|T191|SY|703604002|SNOMEDCT_US|PEComa, benign|8714/0
C3839685|T191|PT|703604002|SNOMEDCT_US|Perivascular epithelioid tumor, benign|8714/0
C3839685|T191|PTGB|703604002|SNOMEDCT_US|Perivascular epithelioid tumour, benign|8714/0
C3839062|T191|PT|C121792|NCI|Malignant PEComa|8714/3
C3839062|T191|SY|C121792|NCI|Malignant PEComa, NOS|8714/3
C3839062|T191|SY|C121792|NCI|Malignant PEComa, Not Otherwise Specified|8714/3
C3839062|T191|SY|703605001|SNOMEDCT_US|PEComa, malignant|8714/3
C3839062|T191|PT|703605001|SNOMEDCT_US|Perivascular epithelioid tumor, malignant|8714/3
C3839062|T191|PTGB|703605001|SNOMEDCT_US|Perivascular epithelioid tumour, malignant|8714/3
C0027962|T191|PT|0029638|CCPSS|NEVUS MELANOCYTIC|8720/0
C0027962|T191|PT|0044443|CCPSS|NEVUS PIGMENTED|8720/0
C0027962|T191|SY|0000008684|CHV|melanocytic naevi|8720/0
C0027962|T191|SY|0000008684|CHV|melanocytic naevus|8720/0
C0027962|T191|SY|0000008684|CHV|melanocytic nevi|8720/0
C0027962|T191|SY|0000008684|CHV|melanocytic nevus|8720/0
C0027962|T191|PT|0000008684|CHV|mole|8720/0
C0027962|T191|SY|0000008684|CHV|moles|8720/0
C0027962|T191|SY|0000008684|CHV|pigmented mole|8720/0
C0027962|T191|SY|0000008684|CHV|pigmented nevi|8720/0
C0027962|T191|SY|0000008684|CHV|pigmented nevus|8720/0
C0027962|T191|PT|U000489|COSTAR|PIGMENTED MOLE|8720/0
C0027962|T191|PT|NOCODE|COSTAR|Pigmented Nevus|8720/0
C3665593|T191|ET|0727-0083|CSP|mole|8720/0
C3665593|T191|PT|0727-0083|CSP|pigmented nevus|8720/0
C0027962|T191|GT|MELANOSIS|CST|NERVUS PIGMENTED|8720/0
C0027962|T191|GT|MELANOSIS|CST|NEVUS MELANOTIC|8720/0
C0027962|T191|FI|U002796|DXP|NEVUS PIGMENTATION|8720/0
C0027962|T191|SY|HP:0000995|HPO|Beauty mark|8720/0
C0027962|T191|SY|HP:0000995|HPO|Melanocytic naevus|8720/0
C0027962|T191|SY|HP:0000995|HPO|Melanocytic nevi|8720/0
C0027962|T191|PT|HP:0000995|HPO|Melanocytic nevus|8720/0
C0027962|T191|ET|HP:0003764|HPO|Naevi|8720/0
C0027962|T191|SY|HP:0000995|HPO|Nevocellular nevi|8720/0
C0027962|T191|SY|HP:0000995|HPO|Pigmented naevi|8720/0
C0027962|T191|SY|HP:0000995|HPO|Pigmented nevi|8720/0
C0027962|T191|HT|D22|ICD10|Melanocytic naevi|8720/0
C0027962|T191|PT|D22.9|ICD10|Melanocytic naevi, unspecified|8720/0
C0027962|T191|HT|D22|ICD10AE|Melanocytic nevi|8720/0
C0027962|T191|PT|D22.9|ICD10AE|Melanocytic nevi, unspecified|8720/0
C0027962|T191|AB|D22|ICD10CM|Melanocytic nevi|8720/0
C0027962|T191|HT|D22|ICD10CM|Melanocytic nevi|8720/0
C0027962|T191|PT|D22.9|ICD10CM|Melanocytic nevi, unspecified|8720/0
C0027962|T191|AB|D22.9|ICD10CM|Melanocytic nevi, unspecified|8720/0
C0027962|T191|ET|D22|ICD10CM|nevus NOS|8720/0
C0027962|T191|PT|S82007|ICPC2P|Naevus;pigmented|8720/0
C0027962|T191|MTH_PT|S82007|ICPC2P|Nevus;pigmented|8720/0
C0027962|T191|PTN|S82007|ICPC2P|pigmented naevus|8720/0
C0027962|T191|MTH_PTN|S82007|ICPC2P|pigmented nevus|8720/0
C0027962|T191|LLT|10027145|MDR|Melanocytic naevus|8720/0
C0027962|T191|PT|10027145|MDR|Melanocytic naevus|8720/0
C0027962|T191|LLT|10062797|MDR|Melanocytic nevus|8720/0
C0027962|T191|MTH_PT|10027145|MDR|Melanocytic nevus|8720/0
C0027962|T191|LLT|10028677|MDR|Naevi melanocytic|8720/0
C0027962|T191|LLT|10028678|MDR|Naevi pigmented|8720/0
C0027962|T191|LLT|10073897|MDR|Naevus melanotic|8720/0
C0027962|T191|OL|10029218|MDR|Nervus pigmented|8720/0
C0027962|T191|MTH_LLT|10028677|MDR|Nevi melanocytic|8720/0
C0027962|T191|MTH_LLT|10028678|MDR|Nevi pigmented|8720/0
C0027962|T191|LLT|10029385|MDR|Nevus melanotic|8720/0
C0027962|T191|LLT|10035031|MDR|Pigmented naevus|8720/0
C0027962|T191|LLT|10062799|MDR|Pigmented nevus|8720/0
C3665593|T191|SY|277704|MEDCIN|benign pigmented nevus|8720/0
C3665593|T191|PT|277704|MEDCIN|benign pigmented nevus of skin|8720/0
C0027962|T191|PM|D009508|MSH|Melanocytic Nevi|8720/0
C0027962|T191|PM|D009508|MSH|Melanocytic Nevus|8720/0
C0027962|T191|ET|D009508|MSH|Nevi, Melanocytic|8720/0
C0027962|T191|ET|D009508|MSH|Nevi, Pigmented|8720/0
C0027962|T191|ET|D009508|MSH|Nevus, Melanocytic|8720/0
C0027962|T191|MH|D009508|MSH|Nevus, Pigmented|8720/0
C0027962|T191|ET|D009508|MSH|Pigmented Moles|8720/0
C0027962|T191|PM|D009508|MSH|Pigmented Nevi|8720/0
C0027962|T191|PM|D009508|MSH|Pigmented Nevus|8720/0
C0027962|T191|PN|NOCODE|MTH|Melanocytic nevus|8720/0
C3665593|T191|PN|NOCODE|MTH|Melanocytic nevus of skin|8720/0
C0027962|T191|SY|NOCODE|MTH|NEVI MELANOCYTIC|8720/0
C0027962|T191|SY|NOCODE|MTH|NEVI PIGMENTED|8720/0
C0027962|T191|PT|C7570|NCI|Melanocytic Nevus|8720/0
C0027962|T191|SY|C7570|NCI|Melanotic Nevus|8720/0
C0027962|T191|SY|C7570|NCI|Mole|8720/0
C0027962|T191|SY|C7570|NCI|Mole of Skin|8720/0
C0027962|T191|SY|C7570|NCI|Nevus|8720/0
C3665593|T191|PT|C27816|NCI|Pigmented Nevus|8720/0
C0027962|T191|PT|CDR0000046286|NCI_NCI-GLOSS|mole|8720/0
C0027962|T191|PT|CDR0000046271|NCI_NCI-GLOSS|nevus|8720/0
C3665593|T191|SY|Xa99Q|RCD|Melanocytic naevus|8720/0
C3665593|T191|SY|X78Uv|RCD|Melanocytic naevus of skin|8720/0
C3665593|T191|SY|X78Uv|RCD|Mole|8720/0
C3665593|T191|SY|X78Uv|RCD|Mole of skin|8720/0
C3665593|T191|PT|Xa99Q|RCD|Pigmented naevus|8720/0
C3665593|T191|SY|X78Uv|RCD|Pigmented naevus of skin|8720/0
C3665593|T191|SY|Xa99Q|RCDAE|Melanocytic nevus|8720/0
C3665593|T191|SY|X78Uv|RCDAE|Melanocytic nevus of skin|8720/0
C3665593|T191|PT|Xa99Q|RCDAE|Pigmented nevus|8720/0
C3665593|T191|SY|X78Uv|RCDAE|Pigmented nevus of skin|8720/0
C0027962|T191|OA|ByuGN|RCDSA|Melanocytic nevi, unspecif|8720/0
C0027962|T191|OP|ByuGN|RCDSA|Melanocytic nevi, unspecified|8720/0
C0027962|T191|IS|Xa07S|RCDSA|Pigmented nevus NOS|8720/0
C0027962|T191|OA|ByuGN|RCDSY|Melanocytic naevi, unspecif|8720/0
C0027962|T191|OP|ByuGN|RCDSY|Melanocytic naevi, unspecified|8720/0
C0027962|T191|IS|Xa07S|RCDSY|Pigmented naevus NOS|8720/0
C1302707|T191|OAP|400094003|SNOMEDCT_US|Acquired melanocytic naevus|8720/0
C1302707|T191|PTGB|399899001|SNOMEDCT_US|Acquired melanocytic naevus|8720/0
C1302707|T191|OAP|400094003|SNOMEDCT_US|Acquired melanocytic nevus|8720/0
C1302707|T191|PT|399899001|SNOMEDCT_US|Acquired melanocytic nevus|8720/0
C3266058|T191|PTGB|449767002|SNOMEDCT_US|Intramucosal naevus|8720/0
C3266058|T191|PT|449767002|SNOMEDCT_US|Intramucosal nevus|8720/0
C4518825|T191|PTGB|733523000|SNOMEDCT_US|Lentiginous melanocytic naevus|8720/0
C4518825|T191|PT|733523000|SNOMEDCT_US|Lentiginous melanocytic nevus|8720/0
C0027962|T191|PTGB|400096001|SNOMEDCT_US|Melanocytic naevus|8720/0
C0027962|T191|SYGB|21119008|SNOMEDCT_US|Melanocytic naevus|8720/0
C3665593|T191|OAS|109265005|SNOMEDCT_US|Melanocytic naevus of skin|8720/0
C3665593|T191|PTGB|400010006|SNOMEDCT_US|Melanocytic naevus of skin|8720/0
C0027962|T191|PT|400096001|SNOMEDCT_US|Melanocytic nevus|8720/0
C0027962|T191|SY|21119008|SNOMEDCT_US|Melanocytic nevus|8720/0
C3665593|T191|PT|400010006|SNOMEDCT_US|Melanocytic nevus of skin|8720/0
C3665593|T191|OAS|109265005|SNOMEDCT_US|Melanocytic nevus of skin|8720/0
C0027962|T191|SY|400096001|SNOMEDCT_US|Mole|8720/0
C3665593|T191|SY|400010006|SNOMEDCT_US|Mole of skin|8720/0
C0027962|T191|SYGB|21119008|SNOMEDCT_US|Naevus|8720/0
C0027962|T191|SY|21119008|SNOMEDCT_US|Nevus|8720/0
C0027962|T191|OAS|189051001|SNOMEDCT_US|Pigmented naevus|8720/0
C0027962|T191|PTGB|21119008|SNOMEDCT_US|Pigmented naevus|8720/0
C3665593|T191|OAS|109265005|SNOMEDCT_US|Pigmented naevus of skin|8720/0
C3665593|T191|SYGB|400010006|SNOMEDCT_US|Pigmented naevus of skin|8720/0
C0027962|T191|PT|21119008|SNOMEDCT_US|Pigmented nevus|8720/0
C0027962|T191|OAS|189051001|SNOMEDCT_US|Pigmented nevus|8720/0
C3665593|T191|SY|400010006|SNOMEDCT_US|Pigmented nevus of skin|8720/0
C3665593|T191|OAS|109265005|SNOMEDCT_US|Pigmented nevus of skin|8720/0
C0027962|T191|SY|21119008|SNOMEDCT_US|Pigmented nevus, no ICD-O subtype|8720/0
C0027962|T191|SY|21119008|SNOMEDCT_US|Pigmented nevus, no International Classification of Diseases for Oncology subtype|8720/0
C0027962|T191|IS|21119008|SNOMEDCT_US|Pigmented nevus, NOS|8720/0
C0027962|T191|IT|0019|WHO|NAEVI MELANOCYTIC|8720/0
C0027962|T191|IT|0019|WHO|NAEVI PIGMENTED|8720/0
C0346040|T191|SY|0000029975|CHV|in situ melanoma|8720/2
C0346040|T191|PT|0000029975|CHV|melanoma in situ|8720/2
C0346040|T191|HT|D03|ICD10|Melanoma in situ|8720/2
C0346040|T191|PT|D03.9|ICD10|Melanoma in situ, unspecified|8720/2
C0346040|T191|AB|D03|ICD10CM|Melanoma in situ|8720/2
C0346040|T191|HT|D03|ICD10CM|Melanoma in situ|8720/2
C0346040|T191|AB|D03.9|ICD10CM|Melanoma in situ, unspecified|8720/2
C0346040|T191|PT|D03.9|ICD10CM|Melanoma in situ, unspecified|8720/2
C0346040|T191|PT|MTHU048094|ICPC2ICD10ENG|melanoma in situ|8720/2
C0346040|T191|PT|MTHU048120|ICPC2ICD10ENG|melanoma in situ; skin|8720/2
C0346040|T191|PT|MTHU035641|ICPC2ICD10ENG|skin; melanoma in situ|8720/2
C0346040|T191|LLT|10027148|MDR|Melanoma in situ|8720/2
C0346040|T191|PT|274864|MEDCIN|malignant melanoma of skin stage 0|8720/2
C0346040|T191|PT|333245|MEDCIN|Melanoma in situ|8720/2
C0346040|T191|PT|231605|MEDCIN|melanoma in situ of skin|8720/2
C4520764|T191|PN|NOCODE|MTH|Stage 0 Cutaneous Melanoma AJCC v6 and v7|8720/2
C0346040|T191|PN|NOCODE|MTH|Stage 0 Skin Melanoma|8720/2
C4520764|T191|SY|C8423|NCI|Cutaneous Melanoma in situ|8720/2
C4520764|T191|SY|C8423|NCI|Malignant Cutaneous Melanoma in situ|8720/2
C4520764|T191|SY|C8423|NCI|Malignant Skin Melanoma in situ|8720/2
C4520764|T191|SY|TCGA|NCI|Melanoma in situ|8720/2
C4520764|T191|SY|C8423|NCI|Melanoma In Situ|8720/2
C4520764|T191|SY|C8423|NCI|Melanoma in situ of Skin|8720/2
C4520764|T191|SY|C8423|NCI|Melanoma in situ of the Skin|8720/2
C4520764|T191|SY|C8423|NCI|Skin Melanoma in situ|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Cutaneous Melanoma|8720/2
C4520764|T191|PT|C8423|NCI|Stage 0 Cutaneous Melanoma AJCC v6 and v7|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Malignant Cutaneous Melanoma|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Malignant Melanoma|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Malignant Skin Melanoma|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Melanoma|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Melanoma of Skin|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Melanoma of the Skin|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Skin Melanoma AJCC v6|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Skin Melanoma AJCC v6 and v7|8720/2
C4520764|T191|SY|C8423|NCI|Stage 0 Skin Melanoma AJCC v7|8720/2
C4520764|T191|PT|C8423|NCI_CPTAC|Stage 0 Cutaneous Melanoma AJCC v6 and v7|8720/2
C4520764|T191|PT|CDR0000522541|NCI_NCI-GLOSS|melanoma in situ|8720/2
C4520764|T191|PT|CDR0000352156|NCI_NCI-GLOSS|stage 0 melanoma|8720/2
C0346040|T191|SY|CDR0000042623|PDQ|melanoma, stage 0|8720/2
C0346040|T191|PSC|CDR0000042623|PDQ|stage 0 melanoma|8720/2
C0346040|T191|AB|X78TH|RCD|In situ malign melanoma skin|8720/2
C0346040|T191|SY|X78TH|RCD|In situ malignant melanoma of skin|8720/2
C0346040|T191|SY|X78TH|RCD|In situ melanoma of skin|8720/2
C0346040|T191|SY|X78TH|RCD|ISM - In situ melanoma of skin|8720/2
C0346040|T191|SY|X78TH|RCD|ISMM - In situ malignant melanoma of skin|8720/2
C0346040|T191|AB|X78TH|RCD|ISMM - In situ MM of skin|8720/2
C0346040|T191|PT|X77oN|RCD|Melanoma in situ|8720/2
C0346040|T191|PT|X78TH|RCD|Melanoma in situ of skin|8720/2
C0346040|T191|OA|ByuFF|RCDSY|Melanoma in situ, unspecif|8720/2
C0346040|T191|OP|ByuFF|RCDSY|Melanoma in situ, unspecified|8720/2
C0346040|T191|SY|109266006|SNOMEDCT_US|In situ malignant melanoma of skin|8720/2
C0346040|T191|SY|109266006|SNOMEDCT_US|In situ melanoma of skin|8720/2
C0346040|T191|SY|109266006|SNOMEDCT_US|ISM - In situ melanoma of skin|8720/2
C0346040|T191|SY|109266006|SNOMEDCT_US|ISMM - In situ malignant melanoma of skin|8720/2
C0346040|T191|OAP|189758001|SNOMEDCT_US|Melanoma in situ|8720/2
C0346040|T191|OF|189758001|SNOMEDCT_US|Melanoma in situ|8720/2
C0346040|T191|PT|77986002|SNOMEDCT_US|Melanoma in situ|8720/2
C0346040|T191|OAP|189320002|SNOMEDCT_US|Melanoma in situ of skin|8720/2
C0346040|T191|OF|189320002|SNOMEDCT_US|Melanoma in situ of skin|8720/2
C0346040|T191|SY|109266006|SNOMEDCT_US|Melanoma in situ of skin|8720/2
C0025202|T191|ET|0000004558|AOD|melanoma|8720/3
C0025202|T191|SY|BI00601|BI|malignant melanoma|8720/3
C0025202|T191|PT|BI00601|BI|melanoma|8720/3
C0025202|T191|SY|0000007894|CHV|cutaneous melanoma|8720/3
C0025202|T191|SY|0000007894|CHV|malignant melanoma|8720/3
C0025202|T191|SY|0000007894|CHV|malignant melanomas|8720/3
C0025202|T191|SY|0000007894|CHV|melanocarcinoma|8720/3
C0025202|T191|PT|0000007894|CHV|melanoma|8720/3
C0025202|T191|SY|0000007894|CHV|melanoma malignant|8720/3
C0025202|T191|SY|0000007894|CHV|melanoma syndrome|8720/3
C0025202|T191|SY|0000007894|CHV|melanomas|8720/3
C0025202|T191|SY|0000007894|CHV|melanosarcoma|8720/3
C0025202|T191|SY|0000007894|CHV|nevocarcinoma|8720/3
C0025202|T191|PT|467|COSTAR|MALIGNANT MELANOMA|8720/3
C0025202|T191|PT|475|COSTAR|MELANOMA|8720/3
C0025202|T191|PT|2020-2434|CSP|melanoma|8720/3
C0025202|T191|GT|MELANOMA SKIN|CST|MALIGNANT MELANOMA|8720/3
C0025202|T191|GT|MELANOMA SKIN|CST|MELANOMA MALIGNANT|8720/3
C0025202|T191|DI|U001151|DXP|MELANOMA, MALIGNANT|8720/3
C0025202|T191|ET|HP:0002861|HPO|Cancer of skin pigment cells|8720/3
C0025202|T191|SY|HP:0002861|HPO|Malignant melanoma|8720/3
C0025202|T191|PT|HP:0002861|HPO|Melanoma|8720/3
C0025202|T191|PT|MTHU048175|ICPC2ICD10ENG|melanoma|8720/3
C0025202|T191|PT|S77003|ICPC2P|Melanoma|8720/3
C0025202|T191|PTN|S77003|ICPC2P|melanoma|8720/3
C0025202|T191|PT|U002889|LCH|Melanoma|8720/3
C0025202|T191|PT|sh85083381|LCH_NW|Melanoma|8720/3
C0025202|T191|LA|LA14279-6|LNC|Melanoma|8720/3
C0025202|T191|LLT|10025650|MDR|Malignant melanoma|8720/3
C0025202|T191|PT|10025650|MDR|Malignant melanoma|8720/3
C0025202|T191|LLT|10053571|MDR|Melanoma|8720/3
C0025202|T191|LLT|10027150|MDR|Melanoma malignant|8720/3
C0025202|T191|PT|352914|MEDCIN|malignant melanoma|8720/3
C0025202|T191|SY|352914|MEDCIN|malignant neoplasm melanoma|8720/3
C0025202|T191|PT|321|MEDLINEPLUS|Melanoma|8720/3
C0025202|T191|ET|D008545|MSH|Malignant Melanoma|8720/3
C0025202|T191|PM|D008545|MSH|Malignant Melanomas|8720/3
C0025202|T191|MH|D008545|MSH|Melanoma|8720/3
C0025202|T191|PM|D008545|MSH|Melanoma, Malignant|8720/3
C0025202|T191|PM|D008545|MSH|Melanomas|8720/3
C0025202|T191|PM|D008545|MSH|Melanomas, Malignant|8720/3
C0025202|T191|PT|475|MTH|MALIGNANT MELANOMA|8720/3
C0025202|T191|PN|NOCODE|MTH|melanoma|8720/3
C0545071|T191|PN|NOCODE|MTH|Minimal Deviation Melanoma|8720/3
C1334386|T191|SY|C5317|NCI|Leptomeningeal Melanoma|8720/3
C0025202|T191|SY|C3224|NCI|Malignant Melanoma|8720/3
C0025202|T191|PT|C3224|NCI|Melanoma|8720/3
C0025202|T191|SY|TCGA|NCI|Melanoma|8720/3
C1334386|T191|SY|C5317|NCI|Melanoma of Leptomeninges|8720/3
C1334386|T191|SY|C5317|NCI|Melanoma of the Leptomeninges|8720/3
C1334386|T191|PT|C5317|NCI|Meningeal Melanoma|8720/3
C0545071|T191|PT|C48612|NCI|Minimal Deviation Melanoma|8720/3
C0545071|T191|SY|TCGA|NCI|Minimal Deviation Melanoma|8720/3
C0025202|T191|SY|C3224|NCI_CDISC|Malignant Melanoma|8720/3
C0025202|T191|PT|C3224|NCI_CDISC|MELANOMA, MALIGNANT|8720/3
C0025202|T191|PT|C3224|NCI_CPTAC|Melanoma|8720/3
C0025202|T191|PT|10053571|NCI_CTEP-SDC|Melanoma|8720/3
C0025202|T191|PT|C3224|NCI_CTRP|Melanoma|8720/3
C0025202|T191|DN|C3224|NCI_CTRP|Melanoma|8720/3
C0025202|T191|PT|CDR0000045135|NCI_NCI-GLOSS|melanoma|8720/3
C0025202|T191|PT|C3224|NCI_NICHD|Melanoma|8720/3
C0025202|T191|PSC|CDR0000038833|PDQ|melanoma|8720/3
C0025202|T191|PT|Xa99S|RCD|Malignant melanoma|8720/3
C0025202|T191|SY|Xa99S|RCD|MM - Malignant melanoma|8720/3
C0025202|T191|OP|XE1wX|RCDSY|Malignant melanoma NOS|8720/3
C1302571|T191|PT|399634005|SNOMEDCT_US|Choroidal melanoma, diffuse|8720/3
C0025202|T191|PT|2092003|SNOMEDCT_US|Malignant melanoma|8720/3
C0025202|T191|OAS|154501005|SNOMEDCT_US|Malignant melanoma|8720/3
C0025202|T191|OAS|269577007|SNOMEDCT_US|Malignant melanoma|8720/3
C0025202|T191|PT|372244006|SNOMEDCT_US|Malignant melanoma|8720/3
C0025202|T191|SY|2092003|SNOMEDCT_US|Malignant melanoma, no ICD-O subtype|8720/3
C0025202|T191|SY|2092003|SNOMEDCT_US|Malignant melanoma, no International Classification of Diseases for Oncology subtype|8720/3
C0025202|T191|IS|2092003|SNOMEDCT_US|Malignant melanoma, NOS|8720/3
C0545071|T191|SY|399475009|SNOMEDCT_US|MDM - Minimal deviation melanoma|8720/3
C0025202|T191|SY|2092003|SNOMEDCT_US|Melanoma|8720/3
C0025202|T191|OAS|269577007|SNOMEDCT_US|Melanoma - malignant|8720/3
C0025202|T191|OAS|154501005|SNOMEDCT_US|Melanoma - malignant|8720/3
C0025202|T191|IS|2092003|SNOMEDCT_US|Melanoma, NOS|8720/3
C0025202|T191|SY|372244006|SNOMEDCT_US|Melanosarcoma|8720/3
C1334386|T191|PT|726420002|SNOMEDCT_US|Meningeal melanoma|8720/3
C0545071|T191|PT|399475009|SNOMEDCT_US|Minimal deviation melanoma|8720/3
C0025202|T191|SY|2092003|SNOMEDCT_US|MM - Malignant melanoma|8720/3
C1302476|T191|PT|399521000|SNOMEDCT_US|Necrotic melanoma|8720/3
C0025202|T191|PT|1084|WHO|MELANOMA MALIGNANT|8720/3
C0860594|T191|SY|0000050761|CHV|malignant melanoma metastatic|8720/6
C0860594|T191|PT|0000050761|CHV|metastatic malignant melanoma|8720/6
C0860594|T191|LLT|10027480|MDR|Metastatic malignant melanoma|8720/6
C0860594|T191|PT|10027480|MDR|Metastatic malignant melanoma|8720/6
C0860594|T191|PT|31663|MEDCIN|metastatic malignant melanoma|8720/6
C0860594|T191|PT|372158004|SNOMEDCT_US|Malignant melanoma, metastatic|8720/6
C0860594|T191|PT|443493003|SNOMEDCT_US|Metastatic malignant melanoma|8720/6
C0334424|T191|SY|0000029976|CHV|melanoma nodular|8721/3
C0334424|T191|SY|0000029976|CHV|melanomas nodular|8721/3
C0334424|T191|PT|0000029976|CHV|nodular melanoma|8721/3
C0334424|T191|PT|HP:0012058|HPO|Nodular melanoma|8721/3
C0334424|T191|LA|LA27884-8|LNC|Nodular melanoma|8721/3
C0334424|T191|LLT|10029488|MDR|Nodular melanoma|8721/3
C0334424|T191|PT|10029488|MDR|Nodular melanoma|8721/3
C0334424|T191|PT|31664|MEDCIN|nodular melanoma of skin|8721/3
C0334424|T191|SY|C4225|NCI|Nodular Malignant Melanoma|8721/3
C0334424|T191|SY|C4225|NCI|Nodular Malignant Melanoma of Skin|8721/3
C0334424|T191|SY|C4225|NCI|Nodular Malignant Melanoma of the Skin|8721/3
C0334424|T191|SY|C4225|NCI|Nodular Malignant Skin Melanoma|8721/3
C0334424|T191|PT|C4225|NCI|Nodular Melanoma|8721/3
C0334424|T191|SY|TCGA|NCI|Nodular Melanoma|8721/3
C0334424|T191|SY|CDR0000039906|PDQ|malignant melanoma, nodular|8721/3
C0334424|T191|SY|CDR0000039906|PDQ|melanoma, nodular malignant|8721/3
C0334424|T191|PT|CDR0000039906|PDQ|nodular malignant melanoma|8721/3
C0334424|T191|SY|CDR0000039906|PDQ|Nodular Malignant Melanoma of Skin|8721/3
C0334424|T191|SY|CDR0000039906|PDQ|Nodular Malignant Melanoma of the Skin|8721/3
C0334424|T191|SY|CDR0000039906|PDQ|Nodular Malignant Skin Melanoma|8721/3
C0334424|T191|SY|CDR0000039906|PDQ|Nodular Melanoma|8721/3
C0334424|T191|SY|BBE2.|RCD|NM - Nodular melanoma|8721/3
C0334424|T191|SY|X78TD|RCD|NM - Nodular melanoma of skin|8721/3
C0334424|T191|AB|X78TD|RCD|Nodular malig melanoma of skin|8721/3
C0334424|T191|PT|X78TD|RCD|Nodular malignant melanoma of skin|8721/3
C0334424|T191|PT|BBE2.|RCD|Nodular melanoma|8721/3
C0334424|T191|SY|X78TD|RCD|Nodular melanoma of skin|8721/3
C0334424|T191|SY|2142002|SNOMEDCT_US|NM - Nodular melanoma|8721/3
C0334424|T191|SY|254731001|SNOMEDCT_US|NM - Nodular melanoma of skin|8721/3
C0334424|T191|PT|254731001|SNOMEDCT_US|Nodular malignant melanoma of skin|8721/3
C0334424|T191|PT|2142002|SNOMEDCT_US|Nodular melanoma|8721/3
C0334424|T191|SY|254731001|SNOMEDCT_US|Nodular melanoma of skin|8721/3
C0334425|T191|PT|C4226|NCI|Balloon Cell Nevus|8722/0
C0334425|T191|PT|BBE3.|RCD|Balloon cell naevus|8722/0
C0334425|T191|PT|BBE3.|RCDAE|Balloon cell nevus|8722/0
C0334425|T191|PTGB|8276007|SNOMEDCT_US|Balloon cell naevus|8722/0
C0334425|T191|PT|8276007|SNOMEDCT_US|Balloon cell nevus|8722/0
C0334426|T191|PT|352915|MEDCIN|Balloon cell malignant melanoma|8722/3
C0334426|T191|SY|352915|MEDCIN|malignant neoplasm melanoma balloon cell|8722/3
C0334426|T191|PN|NOCODE|MTH|Balloon cell malignant melanoma|8722/3
C0334426|T191|SY|C4227|NCI|Balloon Cell Malignant Melanoma|8722/3
C0334426|T191|SY|C4227|NCI|Balloon Cell Malignant Melanoma of Skin|8722/3
C0334426|T191|SY|C4227|NCI|Balloon Cell Malignant Melanoma of the Skin|8722/3
C0334426|T191|SY|C4227|NCI|Balloon Cell Malignant Skin Melanoma|8722/3
C0334426|T191|PT|C4227|NCI|Balloon Cell Melanoma|8722/3
C0334426|T191|SY|C4227|NCI|Balloon Cell Skin Melanoma|8722/3
C0334426|T191|PT|BBE4.|RCD|Balloon cell melanoma|8722/3
C0334426|T191|PT|403922007|SNOMEDCT_US|Balloon cell malignant melanoma|8722/3
C0334426|T191|PT|39274007|SNOMEDCT_US|Balloon cell melanoma|8722/3
C0474824|T191|SY|0000037070|CHV|halo naevus|8723/0
C0474824|T191|SY|0000037070|CHV|halo nevi|8723/0
C0474824|T191|PT|0000037070|CHV|halo nevus|8723/0
C0474824|T191|SY|0000037070|CHV|halos nevi|8723/0
C0474824|T191|SY|0000037070|CHV|naevus halo|8723/0
C0474824|T191|SY|0000037070|CHV|nevus halo|8723/0
C0474824|T191|PTN|S82014|ICPC2P|halo naevus|8723/0
C0474824|T191|MTH_PTN|S82014|ICPC2P|halo nevus|8723/0
C0474824|T191|PT|S82014|ICPC2P|Naevus;halo|8723/0
C0474824|T191|MTH_PT|S82014|ICPC2P|Nevus;halo|8723/0
C0474824|T191|LLT|10019097|MDR|Halo naevus|8723/0
C0474824|T191|LLT|10062794|MDR|Halo nevus|8723/0
C0474824|T191|ET|D055882|MSH|Halo Nevi|8723/0
C0474824|T191|PM|D055882|MSH|Halo Nevus|8723/0
C0474824|T191|ET|D055882|MSH|Leukoderma Acquisitum Centrifugum of Sutton|8723/0
C0474824|T191|ET|D055882|MSH|Nevi, Halo|8723/0
C0474824|T191|MH|D055882|MSH|Nevus, Halo|8723/0
C0474824|T191|PN|NOCODE|MTH|Halo nevus|8723/0
C0474824|T191|PT|C7602|NCI|Halo Nevus|8723/0
C0474824|T191|PT|XaBAv|RCD|Halo naevus|8723/0
C0474824|T191|SY|XaBAv|RCD|Sutton's naevus|8723/0
C0474824|T191|PT|XaBAv|RCDAE|Halo nevus|8723/0
C0474824|T191|SY|XaBAv|RCDAE|Sutton's nevus|8723/0
C0474824|T191|PT|BBE5.|RCDSA|Halo nevus|8723/0
C0474824|T191|PT|BBE5.|RCDSY|Halo naevus|8723/0
C0474824|T191|OAP|307602007|SNOMEDCT_US|Halo naevus|8723/0
C0474824|T191|PTGB|78325005|SNOMEDCT_US|Halo naevus|8723/0
C0474824|T191|PTGB|398028009|SNOMEDCT_US|Halo naevus|8723/0
C0474824|T191|PT|398028009|SNOMEDCT_US|Halo nevus|8723/0
C0474824|T191|PT|78325005|SNOMEDCT_US|Halo nevus|8723/0
C0474824|T191|OAP|307602007|SNOMEDCT_US|Halo nevus|8723/0
C0474824|T191|OAS|307602007|SNOMEDCT_US|Sutton's naevus|8723/0
C0474824|T191|SYGB|398028009|SNOMEDCT_US|Sutton's naevus|8723/0
C0474824|T191|OAS|307602007|SNOMEDCT_US|Sutton's nevus|8723/0
C0474824|T191|SY|398028009|SNOMEDCT_US|Sutton's nevus|8723/0
C0334427|T191|SY|C4228|NCI|Regressing Malignant Melanoma|8723/3
C0334427|T191|PT|C4228|NCI|Regressing Melanoma|8723/3
C0334427|T191|PT|C4228|NCI_CPTAC|Regressing Melanoma|8723/3
C0334427|T191|PT|X77oJ|RCD|Regressing malignant melanoma|8723/3
C0334427|T191|AB|X77oJ|RCDSY|Malign melanoma, regressing|8723/3
C0334427|T191|SY|X77oJ|RCDSY|Malignant melanoma, regressing|8723/3
C0334427|T191|PT|39896009|SNOMEDCT_US|Malignant melanoma, regressing|8723/3
C0334427|T191|OAP|189750008|SNOMEDCT_US|Regressing malignant melanoma|8723/3
C0334427|T191|OF|189750008|SNOMEDCT_US|Regressing malignant melanoma|8723/3
C0334430|T191|SY|C4229|NCI|Neural Nevus|8725/0
C0334430|T191|PT|C4229|NCI|Neuronevus|8725/0
C0334430|T191|PT|BBE7.|RCD|Neuronaevus|8725/0
C0334430|T191|PT|BBE7.|RCDAE|Neuronevus|8725/0
C0334430|T191|PTGB|17930004|SNOMEDCT_US|Neuronaevus|8725/0
C0334430|T191|PT|17930004|SNOMEDCT_US|Neuronevus|8725/0
C2004458|T191|PT|MTHU047127|ICPC2ICD10ENG|magnocellular; nevus, unspecified site|8726/0
C2004458|T191|PT|MTHU048090|ICPC2ICD10ENG|melanocytoma; eyeball|8726/0
C2004458|T191|PT|MTHU051600|ICPC2ICD10ENG|nevus; magnocellular, unspecified site|8726/0
C2004458|T191|LLT|10057531|MDR|Ocular melanocytoma|8726/0
C2004458|T191|PT|38592|MEDCIN|ocular melanocytoma|8726/0
C2004458|T191|SY|C4230|NCI|Magnocellular Nevus|8726/0
C2004458|T191|SY|C4230|NCI|Melanocytoma of Eyeball|8726/0
C2004458|T191|PT|C4230|NCI|Melanocytoma of the Eyeball|8726/0
C2004458|T191|PT|BBE8.|RCD|Magnocellular naevus|8726/0
C2004458|T191|SY|BBE8.|RCD|Melanocytoma of the eyeball|8726/0
C2004458|T191|PT|BBE8.|RCDAE|Magnocellular nevus|8726/0
C2004458|T191|PTGB|26325004|SNOMEDCT_US|Magnocellular naevus|8726/0
C2004458|T191|PT|26325004|SNOMEDCT_US|Magnocellular nevus|8726/0
C2004458|T191|SY|26325004|SNOMEDCT_US|Melanocytoma of the eyeball|8726/0
C0205748|T191|PT|BI00571|BI|atypical nevi|8727/0
C0205748|T191|PT|BI00584|BI|dysplastic nevi|8727/0
C0205748|T191|SY|0000020703|CHV|atypical naevus|8727/0
C0205748|T191|SY|0000020703|CHV|atypical nevi|8727/0
C0205748|T191|SY|0000020703|CHV|atypical nevis|8727/0
C0205748|T191|SY|0000020703|CHV|atypical nevus|8727/0
C0205748|T191|SY|0000020703|CHV|dysplastic naevus|8727/0
C0205748|T191|PT|0000020703|CHV|dysplastic nevi|8727/0
C0205748|T191|SY|0000020703|CHV|dysplastic nevis|8727/0
C0205748|T191|SY|0000020703|CHV|dysplastic nevus|8727/0
C0205748|T191|SY|0000020703|CHV|naevus dysplastic|8727/0
C0205748|T191|SY|HP:0001062|HPO|Atypical mole|8727/0
C0205748|T191|PT|HP:0001062|HPO|Atypical nevus|8727/0
C0205748|T191|ET|HP:0001062|HPO|Dysplastic Nevus|8727/0
C0205748|T191|ET|D22|ICD10CM|atypical nevus|8727/0
C0205748|T191|PT|10062805|MDR|Dysplastic naevus|8727/0
C0205748|T191|LLT|10062805|MDR|Dysplastic naevus|8727/0
C0205748|T191|LLT|10013961|MDR|Dysplastic nevus|8727/0
C0205748|T191|MTH_PT|10062805|MDR|Dysplastic nevus|8727/0
C0205748|T191|PT|214042|MEDCIN|dysplastic nevus|8727/0
C0205748|T191|PEP|D004416|MSH|Dysplastic Nevi|8727/0
C0205748|T191|PM|D004416|MSH|Dysplastic Nevus|8727/0
C0205748|T191|PM|D004416|MSH|Nevi, Dysplastic|8727/0
C0205748|T191|ET|D004416|MSH|Nevus, Dysplastic|8727/0
C0205748|T191|PN|NOCODE|MTH|Dysplastic Nevus|8727/0
C0205748|T191|SY|C3694|NCI|Atypical Nevus|8727/0
C0205748|T191|SY|C3694|NCI|Clark Nevus|8727/0
C0205748|T191|SY|C3694|NCI|Clark's Nevus|8727/0
C0205748|T191|PT|C3694|NCI|Dysplastic Nevus|8727/0
C0205748|T191|SY|C3694|NCI|Lentiginous Nevus|8727/0
C0205748|T191|AB|C3694|NCI|NAD|8727/0
C0205748|T191|SY|C3694|NCI|Nevus with Architectural Disorder|8727/0
C0205748|T191|SY|C3694|NCI|Nevus with Architectural Disorder and Cytologic Atypia of Melanocytes|8727/0
C0205748|T191|PT|CDR0000046161|NCI_NCI-GLOSS|dysplastic nevi|8727/0
C0205748|T191|PT|CDR0000044279|NCI_NCI-GLOSS|dysplastic nevus|8727/0
C0205748|T191|SY|X77oS|RCD|Atypical naevus|8727/0
C0205748|T191|SY|X78VI|RCD|Atypical naevus of skin|8727/0
C0205748|T191|SY|X77oS|RCD|DN - Dysplastic naevus|8727/0
C0205748|T191|PT|X77oS|RCD|Dysplastic naevus|8727/0
C0205748|T191|PT|X78VI|RCD|Dysplastic naevus of skin|8727/0
C0205748|T191|SY|X77oS|RCDAE|Atypical nevus|8727/0
C0205748|T191|SY|X78VI|RCDAE|Atypical nevus of skin|8727/0
C0205748|T191|SY|X77oS|RCDAE|DN - Dysplastic nevus|8727/0
C0205748|T191|PT|X77oS|RCDAE|Dysplastic nevus|8727/0
C0205748|T191|PT|X78VI|RCDAE|Dysplastic nevus of skin|8727/0
C0205748|T191|SYGB|61814002|SNOMEDCT_US|Atypical naevus|8727/0
C0205748|T191|SYGB|254818000|SNOMEDCT_US|Atypical naevus of skin|8727/0
C0205748|T191|SY|61814002|SNOMEDCT_US|Atypical nevus|8727/0
C0205748|T191|SY|254818000|SNOMEDCT_US|Atypical nevus of skin|8727/0
C0205748|T191|SYGB|61814002|SNOMEDCT_US|DN - Dysplastic naevus|8727/0
C0205748|T191|SY|61814002|SNOMEDCT_US|DN - Dysplastic nevus|8727/0
C0205748|T191|OF|189759009|SNOMEDCT_US|Dysplastic naevus|8727/0
C0205748|T191|PTGB|61814002|SNOMEDCT_US|Dysplastic naevus|8727/0
C0205748|T191|OAP|189759009|SNOMEDCT_US|Dysplastic naevus|8727/0
C0205748|T191|PTGB|254818000|SNOMEDCT_US|Dysplastic naevus of skin|8727/0
C0205748|T191|OAP|189759009|SNOMEDCT_US|Dysplastic nevus|8727/0
C0205748|T191|PT|61814002|SNOMEDCT_US|Dysplastic nevus|8727/0
C0205748|T191|PT|254818000|SNOMEDCT_US|Dysplastic nevus of skin|8727/0
C1266112|T191|SY|C6890|NCI|Diffuse Melanocytosis|8728/0
C1266112|T191|SY|C6890|NCI|Diffuse Melanosis|8728/0
C1266112|T191|SY|C6890|NCI|Diffuse Meningeal Melanocytosis|8728/0
C1266112|T191|PT|C6890|NCI|Meningeal Melanocytosis|8728/0
C1266112|T191|PT|128729004|SNOMEDCT_US|Diffuse melanocytosis|8728/0
C1266113|T191|PT|356639|MEDCIN|Melanocytoma of meninges|8728/1
C1266113|T191|SY|356639|MEDCIN|meningeal neoplasm primary melanocytoma|8728/1
C1266113|T191|PN|NOCODE|MTH|Meningeal melanocytoma|8728/1
C1266113|T191|SY|C4662|NCI|Leptomeningeal Melanocytoma|8728/1
C1266113|T191|SY|C4662|NCI|Melanocytoma of Meninges|8728/1
C1266113|T191|SY|C4662|NCI|Melanocytoma of the Meninges|8728/1
C1266113|T191|PT|C4662|NCI|Meningeal Melanocytoma|8728/1
C1266113|T191|SY|C4662|NCI|Meninges Melanocytoma|8728/1
C1266113|T191|PT|Xa0RR|RCD|Melanocytoma of meninges|8728/1
C1266113|T191|PT|277527003|SNOMEDCT_US|Melanocytoma of meninges|8728/1
C1266113|T191|PT|128730009|SNOMEDCT_US|Meningeal melanocytoma|8728/1
C1266114|T191|PT|235569|MEDCIN|malignant melanomatosis of meninges|8728/3
C1266114|T191|SY|235569|MEDCIN|meningeal melanomatosis|8728/3
C1266114|T191|PN|NOCODE|MTH|Meningeal melanomatosis|8728/3
C1266114|T191|SY|C6891|NCI|Leptomeningeal Melanomatosis|8728/3
C1266114|T191|PT|C6891|NCI|Meningeal Melanomatosis|8728/3
C1266114|T191|PT|128731008|SNOMEDCT_US|Meningeal melanomatosis|8728/3
C0334432|T191|SY|0000029978|CHV|achromic naevus|8730/0
C0334432|T191|SY|0000029978|CHV|achromic nevus|8730/0
C0334432|T191|SY|0000029978|CHV|naevus depigmentosus|8730/0
C0334432|T191|SY|0000029978|CHV|nevus achromic|8730/0
C0334432|T191|PT|0000029978|CHV|nevus depigmentosus|8730/0
C0334432|T191|SY|0000029978|CHV|non-pigmented nevus|8730/0
C0334432|T191|PT|C27095|NCI|Nonpigmented Nevus|8730/0
C0334432|T191|SY|BBE9.|RCD|Achromic naevus|8730/0
C0334432|T191|SY|BBE9.|RCD|Hypochromic naevus|8730/0
C0334432|T191|SY|BBE9.|RCD|Naevus depigmentosus|8730/0
C0334432|T191|PT|BBE9.|RCD|Non-pigmented naevus|8730/0
C0334432|T191|SY|BBE9.|RCDAE|Achromic nevus|8730/0
C0334432|T191|SY|BBE9.|RCDAE|Hypochromic nevus|8730/0
C0334432|T191|SY|BBE9.|RCDAE|Nevus depigmentosus|8730/0
C0334432|T191|PT|BBE9.|RCDAE|Non-pigmented nevus|8730/0
C0334432|T191|PTGB|403541001|SNOMEDCT_US|Achromic naevus|8730/0
C0334432|T191|SYGB|112680001|SNOMEDCT_US|Achromic naevus|8730/0
C0334432|T191|SY|112680001|SNOMEDCT_US|Achromic nevus|8730/0
C0334432|T191|PT|403541001|SNOMEDCT_US|Achromic nevus|8730/0
C0334432|T191|SYGB|403541001|SNOMEDCT_US|Hypochromic naevus|8730/0
C0334432|T191|SYGB|112680001|SNOMEDCT_US|Hypochromic naevus|8730/0
C0334432|T191|SY|112680001|SNOMEDCT_US|Hypochromic nevus|8730/0
C0334432|T191|SY|403541001|SNOMEDCT_US|Hypochromic nevus|8730/0
C0334432|T191|SYGB|403541001|SNOMEDCT_US|Naevus depigmentosus|8730/0
C0334432|T191|SYGB|112680001|SNOMEDCT_US|Naevus depigmentosus|8730/0
C0334432|T191|SY|403541001|SNOMEDCT_US|Nevus depigmentosus|8730/0
C0334432|T191|SY|112680001|SNOMEDCT_US|Nevus depigmentosus|8730/0
C0334432|T191|SYGB|112680001|SNOMEDCT_US|Non-pigmented naevus|8730/0
C0334432|T191|SY|112680001|SNOMEDCT_US|Non-pigmented nevus|8730/0
C0334432|T191|PTGB|112680001|SNOMEDCT_US|Nonpigmented naevus|8730/0
C0334432|T191|PT|112680001|SNOMEDCT_US|Nonpigmented nevus|8730/0
C0206735|T191|LLT|10072454|MDR|Amelanotic melanoma|8730/3
C0206735|T191|PM|D018328|MSH|Amelanotic Melanoma|8730/3
C0206735|T191|PM|D018328|MSH|Amelanotic Melanomas|8730/3
C0206735|T191|MH|D018328|MSH|Melanoma, Amelanotic|8730/3
C0206735|T191|PM|D018328|MSH|Melanomas, Amelanotic|8730/3
C0206735|T191|PN|NOCODE|MTH|Melanoma, Amelanotic|8730/3
C0206735|T191|PT|C3802|NCI|Amelanotic Melanoma|8730/3
C0206735|T191|PT|C3802|NCI_CDISC|MELANOMA, AMELANOTIC, MALIGNANT|8730/3
C0206735|T191|PT|C3802|NCI_CPTAC|Amelanotic Melanoma|8730/3
C0206735|T191|PT|CDR0000044526|NCI_NCI-GLOSS|amelanotic melanoma|8730/3
C0206735|T191|PT|BBEA.|RCD|Amelanotic melanoma|8730/3
C0206735|T191|PT|70594002|SNOMEDCT_US|Amelanotic melanoma|8730/3
C0334433|T191|SY|0000029979|CHV|junction nevus|8740/0
C0334433|T191|SY|0000029979|CHV|junctional melanocytic nevus|8740/0
C0334433|T191|SY|0000029979|CHV|junctional naevus|8740/0
C0334433|T191|PT|0000029979|CHV|junctional nevus|8740/0
C0334433|T191|PTN|S82015|ICPC2P|junctional naevus|8740/0
C0334433|T191|MTH_PTN|S82015|ICPC2P|junctional nevus|8740/0
C0334433|T191|PT|S82015|ICPC2P|Naevus;junctional|8740/0
C0334433|T191|MTH_PT|S82015|ICPC2P|Nevus;junctional|8740/0
C0334433|T191|LLT|10023245|MDR|Junctional naevus|8740/0
C0334433|T191|LLT|10062796|MDR|Junctional nevus|8740/0
C0334433|T191|SY|C4231|NCI|Intraepidermal Nevus|8740/0
C0334433|T191|SY|C4231|NCI|Intraepidermal Nevus of Skin|8740/0
C0334433|T191|SY|C4231|NCI|Intraepidermal Nevus of the Skin|8740/0
C0334433|T191|SY|C4231|NCI|Junction Nevus|8740/0
C0334433|T191|SY|C4231|NCI|Junctional Melanocytic Nevus|8740/0
C0334433|T191|SY|C4231|NCI|Junctional Melanocytoma|8740/0
C0334433|T191|PT|C4231|NCI|Junctional Nevus|8740/0
C0334433|T191|SY|C4231|NCI|Junctional Nevus of Skin|8740/0
C0334433|T191|SY|C4231|NCI|Junctional Nevus of the Skin|8740/0
C0334433|T191|SY|C4231|NCI|Junctional Skin Nevus|8740/0
C0334433|T191|PT|CDR0000044285|NCI_NCI-GLOSS|junctional nevus|8740/0
C0334433|T191|SY|X78Ux|RCD|Intra-epidermal naevus of skin|8740/0
C0334433|T191|SY|BBEB.|RCD|Intraepidermal naevus|8740/0
C0334433|T191|AB|X78Ux|RCD|Junction melanocyt naevus skin|8740/0
C0334433|T191|SY|BBEB.|RCD|Junction naevus|8740/0
C0334433|T191|SY|BBEB.|RCD|Junctional melanocytic naevus|8740/0
C0334433|T191|PT|X78Ux|RCD|Junctional melanocytic naevus of skin|8740/0
C0334433|T191|PT|BBEB.|RCD|Junctional naevus|8740/0
C0334433|T191|SY|X78Ux|RCDAE|Intra-epidermal nevus of skin|8740/0
C0334433|T191|SY|BBEB.|RCDAE|Intraepidermal nevus|8740/0
C0334433|T191|AB|X78Ux|RCDAE|Junction melanocyt nevus skin|8740/0
C0334433|T191|SY|BBEB.|RCDAE|Junction nevus|8740/0
C0334433|T191|SY|BBEB.|RCDAE|Junctional melanocytic nevus|8740/0
C0334433|T191|PT|X78Ux|RCDAE|Junctional melanocytic nevus of skin|8740/0
C0334433|T191|PT|BBEB.|RCDAE|Junctional nevus|8740/0
C0334433|T191|SYGB|254802006|SNOMEDCT_US|Intra-epidermal naevus of skin|8740/0
C0334433|T191|SY|254802006|SNOMEDCT_US|Intra-epidermal nevus of skin|8740/0
C0334433|T191|SYGB|30494009|SNOMEDCT_US|Intraepidermal naevus|8740/0
C0334433|T191|SY|30494009|SNOMEDCT_US|Intraepidermal nevus|8740/0
C0334433|T191|SYGB|30494009|SNOMEDCT_US|Junction naevus|8740/0
C0334433|T191|SY|30494009|SNOMEDCT_US|Junction nevus|8740/0
C0334433|T191|SYGB|30494009|SNOMEDCT_US|Junctional melanocytic naevus|8740/0
C0334433|T191|PTGB|254802006|SNOMEDCT_US|Junctional melanocytic naevus of skin|8740/0
C0334433|T191|SY|30494009|SNOMEDCT_US|Junctional melanocytic nevus|8740/0
C0334433|T191|PT|254802006|SNOMEDCT_US|Junctional melanocytic nevus of skin|8740/0
C0334433|T191|SY|30494009|SNOMEDCT_US|Junctional melanocytoma|8740/0
C0334433|T191|PTGB|30494009|SNOMEDCT_US|Junctional naevus|8740/0
C0334433|T191|PT|30494009|SNOMEDCT_US|Junctional nevus|8740/0
C0334433|T191|IS|30494009|SNOMEDCT_US|Junctional nevus, NOS|8740/0
C0334434|T191|PT|231652|MEDCIN|malignant melanoma of skin in junctional nevus|8740/3
C0334434|T191|SY|C4232|NCI|Malignant Melanoma in Junctional Nevus|8740/3
C0334434|T191|SY|C4232|NCI|Malignant Melanoma of Skin in Junctional Nevus|8740/3
C0334434|T191|SY|C4232|NCI|Malignant Melanoma of the Skin in Junctional Nevus|8740/3
C0334434|T191|SY|C4232|NCI|Malignant Skin Melanoma in Junctional Nevus|8740/3
C0334434|T191|PT|C4232|NCI|Melanoma in Junctional Nevus|8740/3
C0334434|T191|AB|BBEC.|RCD|Malig melanoma in junct naevus|8740/3
C0334434|T191|PT|BBEC.|RCD|Malignant melanoma in junctional naevus|8740/3
C0334434|T191|AB|BBEC.|RCDAE|Malig melanoma in junct nevus|8740/3
C0334434|T191|PT|BBEC.|RCDAE|Malignant melanoma in junctional nevus|8740/3
C0334434|T191|PTGB|915007|SNOMEDCT_US|Malignant melanoma in junctional naevus|8740/3
C0334434|T191|PT|915007|SNOMEDCT_US|Malignant melanoma in junctional nevus|8740/3
C0334435|T191|PT|231606|MEDCIN|precancerous melanosis of skin|8741/2
C0334435|T191|PN|NOCODE|MTH|Precancerous melanosis|8741/2
C0334435|T191|PT|C4233|NCI|Precancerous Melanosis|8741/2
C0334435|T191|AB|X508j|RCD|Melanosis circumscr precancer|8741/2
C0334435|T191|SY|X508j|RCD|Melanosis circumscripta precancerosa of Dubreuilh|8741/2
C0334435|T191|PT|X508j|RCD|Precancerous melanosis|8741/2
C0334435|T191|OP|BBED.|RCDSY|Precancerous melanosis NOS|8741/2
C0334435|T191|SY|238701007|SNOMEDCT_US|Melanosis circumscripta precancerosa of Dubreuilh|8741/2
C0334435|T191|OAP|253036005|SNOMEDCT_US|Precancerous melanosis|8741/2
C0334435|T191|PT|238701007|SNOMEDCT_US|Precancerous melanosis|8741/2
C0334435|T191|PT|38969003|SNOMEDCT_US|Precancerous melanosis|8741/2
C0334435|T191|IS|38969003|SNOMEDCT_US|Precancerous melanosis, NOS|8741/2
C0431098|T191|PT|C66753|NCI|Malignant Melanoma in Precancerous Melanosis|8741/3
C0431098|T191|AB|BBEE.|RCD|Malig melanoma in preca melais|8741/3
C0431098|T191|PT|BBEE.|RCD|Malignant melanoma in precancerous melais|8741/3
C0431098|T191|SY|18450009|SNOMEDCT_US|Malignant melanoma in melanosis|8741/3
C0431098|T191|IS|18450009|SNOMEDCT_US|Malignant melanoma in precancerous melais|8741/3
C0431098|T191|PT|18450009|SNOMEDCT_US|Malignant melanoma in precancerous melanosis|8741/3
C0149722|T191|SY|0000016666|CHV|hutchinson's melanotic freckle|8742/2
C0149722|T191|PT|0000016666|CHV|lentigo maligna|8742/2
C0149722|T191|SY|0000016666|CHV|lentigo malignant|8742/2
C0149722|T191|SY|0000016666|CHV|melanotic freckle|8742/2
C0149722|T191|PT|U000411|COSTAR|LENTIGO MALIGNA|8742/2
C0149722|T191|OP|S80004|ICPC2P|Hutchinsons melanotic freckle|8742/2
C0149722|T191|PT|S79009|ICPC2P|Hutchinsons melanotic freckle|8742/2
C0149722|T191|PTN|S79009|ICPC2P|Hutchinsons melanotic freckle|8742/2
C0149722|T191|LLT|10020473|MDR|Hutchinson's melanotic freckle|8742/2
C0149722|T191|OL|10020476|MDR|Hutchison's melanotic freckle|8742/2
C0149722|T191|LLT|10024218|MDR|Lentigo maligna|8742/2
C0149722|T191|PT|10024218|MDR|Lentigo maligna|8742/2
C0149722|T191|LLT|10027160|MDR|Melanotic freckle of Hutchinson|8742/2
C0149722|T191|PT|314842|MEDCIN|lentigo maligna|8742/2
C0149722|T191|PM|D018327|MSH|Freckle, Hutchinson's Melanotic|8742/2
C0149722|T191|ET|D018327|MSH|Freckle, Melanotic|8742/2
C0149722|T191|PM|D018327|MSH|Freckles, Melanotic|8742/2
C0149722|T191|PM|D018327|MSH|Hutchinson Melanotic Freckle|8742/2
C0149722|T191|MH|D018327|MSH|Hutchinson's Melanotic Freckle|8742/2
C0149722|T191|PM|D018327|MSH|Hutchinsons Melanotic Freckle|8742/2
C0149722|T191|ET|D018327|MSH|Lentigo Maligna|8742/2
C0149722|T191|ET|D018327|MSH|Lentigo, Malignant|8742/2
C0149722|T191|PM|D018327|MSH|Lentigos, Malignant|8742/2
C0149722|T191|PM|D018327|MSH|Malignant Lentigo|8742/2
C0149722|T191|PM|D018327|MSH|Malignant Lentigos|8742/2
C0149722|T191|ET|D018327|MSH|Melanotic Freckle|8742/2
C0149722|T191|PM|D018327|MSH|Melanotic Freckle, Hutchinson's|8742/2
C0149722|T191|PM|D018327|MSH|Melanotic Freckles|8742/2
C0149722|T191|SY|C43372|NCI|Hutchinson's Melanotic Freckle|8742/2
C0149722|T191|PT|C43372|NCI|Lentigo Maligna|8742/2
C0149722|T191|PT|Xa99X|RCD|Lentigo maligna|8742/2
C0149722|T191|SY|Xa99X|RCD|LM - Lentigo maligna|8742/2
C0149722|T191|OA|BBEF.|RCDSY|Hutchinson melanot freckle|8742/2
C0149722|T191|OP|BBEF.|RCDSY|Hutchinson's melanotic freckle|8742/2
C0149722|T191|SY|61217001|SNOMEDCT_US|Hutchinson melanotic freckle|8742/2
C0149722|T191|PT|61217001|SNOMEDCT_US|Hutchinson's melanotic freckle|8742/2
C0149722|T191|IS|61217001|SNOMEDCT_US|Hutchinson's melanotic freckle, NOS|8742/2
C0149722|T191|SY|61217001|SNOMEDCT_US|Lentigo maligna|8742/2
C0149722|T191|PT|302836005|SNOMEDCT_US|Lentigo maligna|8742/2
C0149722|T191|SY|302836005|SNOMEDCT_US|LM - Lentigo maligna|8742/2
C0149722|T191|IT|0019|WHO|LENTIGO MALIGNA|8742/2
C2739810|T191|PT|HP:0012059|HPO|Lentigo maligna melanoma|8742/3
C2739810|T191|LA|LA27885-5|LNC|Lentigo maligna melanoma|8742/3
C2739810|T191|LLT|10024219|MDR|Lentigo maligna melanoma|8742/3
C2739810|T191|PT|31662|MEDCIN|lentigo maligna melanoma of skin|8742/3
C2739810|T191|PT|C9151|NCI|Lentigo Maligna Melanoma|8742/3
C2739810|T191|SY|TCGA|NCI|Lentigo Maligna Melanoma|8742/3
C2739810|T191|SY|C9151|NCI|Malignant Lentigo Melanoma|8742/3
C2739810|T191|DN|C9151|NCI_CTRP|Lentigo Maligna Melanoma|8742/3
C2739810|T191|PT|CDR0000039902|PDQ|lentigo maligna malignant melanoma|8742/3
C2739810|T191|SY|CDR0000039902|PDQ|Lentigo Maligna Melanoma|8742/3
C2739810|T191|SY|CDR0000039902|PDQ|Malignant Lentigo Melanoma|8742/3
C2739810|T191|SY|CDR0000039902|PDQ|malignant melanoma, lentigo maligna malignant|8742/3
C2739810|T191|SY|CDR0000039902|PDQ|melanoma, lentigo maligna malignant|8742/3
C2739810|T191|PT|Xa99Y|RCD|Lentigo maligna melanoma|8742/3
C2739810|T191|SY|Xa99Y|RCD|LMM - Lentigo maligna melanoma|8742/3
C2739810|T191|OP|BBEG.|RCDSY|Malignant melanoma in Hutchinson's melanotic freckle|8742/3
C2739810|T191|OA|BBEG.|RCDSY|MM Hutchin melanot freckle|8742/3
C2739810|T191|SY|44474009|SNOMEDCT_US|Lentigo maligna melanoma|8742/3
C2739810|T191|PT|302837001|SNOMEDCT_US|Lentigo maligna melanoma|8742/3
C2739810|T191|SY|302837001|SNOMEDCT_US|LMM - Lentigo maligna melanoma|8742/3
C2739810|T191|SY|44474009|SNOMEDCT_US|Malignant melanoma in Hutchinson melanotic freckle|8742/3
C2739810|T191|PT|44474009|SNOMEDCT_US|Malignant melanoma in Hutchinson's melanotic freckle|8742/3
C0334438|T191|SY|0000029980|CHV|melanoma superficial spreading|8743/3
C0334438|T191|PT|0000029980|CHV|superficial spreading melanoma|8743/3
C0334438|T191|PT|HP:0012057|HPO|Superficial spreading melanoma|8743/3
C0334438|T191|LA|LA27883-0|LNC|Superficial spreading melanoma|8743/3
C0334438|T191|LLT|10042547|MDR|Superficial spreading melanoma|8743/3
C0334438|T191|LLT|10042553|MDR|Superficial spreading melanoma stage unspecified|8743/3
C0334438|T191|PT|10042553|MDR|Superficial spreading melanoma stage unspecified|8743/3
C0334438|T191|SY|31665|MEDCIN|superficial spreading malignant melanoma|8743/3
C0334438|T191|PT|31665|MEDCIN|superficial spreading malignant melanoma of skin|8743/3
C0334438|T191|PN|NOCODE|MTH|Superficial spreading malignant melanoma of skin|8743/3
C0334438|T191|SY|C9152|NCI|Cutaneous Superficial Spreading Melanoma|8743/3
C0334438|T191|SY|C9152|NCI|Pagetoid Melanoma|8743/3
C0334438|T191|AB|C9152|NCI|SSM|8743/3
C0334438|T191|SY|C9152|NCI|Superficial Spreading Malignant Melanoma of Skin|8743/3
C0334438|T191|SY|C9152|NCI|Superficial Spreading Malignant Melanoma of the Skin|8743/3
C0334438|T191|SY|C9152|NCI|Superficial Spreading Malignant Skin Melanoma|8743/3
C0334438|T191|PT|C9152|NCI|Superficial Spreading Melanoma|8743/3
C0334438|T191|SY|TCGA|NCI|Superficial Spreading Melanoma|8743/3
C0334438|T191|SY|C9152|NCI|Superficial Spreading Melanoma of Skin|8743/3
C0334438|T191|SY|C9152|NCI|Superficial Spreading Melanoma of the Skin|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|Cutaneous Superficial Spreading Melanoma|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|malignant melanoma, superficial spreading|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|melanoma, superficial spreading malignant|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|Pagetoid Melanoma|8743/3
C0334438|T191|AB|CDR0000039903|PDQ|SSM|8743/3
C0334438|T191|PT|CDR0000039903|PDQ|superficial spreading malignant melanoma|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|Superficial Spreading Malignant Melanoma of Skin|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|Superficial Spreading Malignant Melanoma of the Skin|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|Superficial Spreading Malignant Skin Melanoma|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|Superficial Spreading Melanoma|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|Superficial Spreading Melanoma of Skin|8743/3
C0334438|T191|SY|CDR0000039903|PDQ|Superficial Spreading Melanoma of the Skin|8743/3
C0334438|T191|AB|X78TC|RCD|SMM - Superfic spread melanoma|8743/3
C0334438|T191|SY|X78TC|RCD|SMM - Superficial spreading melanoma of skin|8743/3
C0334438|T191|AB|BBEH.|RCD|SSM - Superfic spread melanoma|8743/3
C0334438|T191|SY|BBEH.|RCD|SSM - Superficial spreading melanoma|8743/3
C0334438|T191|AB|BBEH.|RCD|SSMM - Superfic spread melanom|8743/3
C0334438|T191|SY|X78TC|RCD|SSMM - Superficial spreading malignant melanoma of skin|8743/3
C0334438|T191|SY|BBEH.|RCD|SSMM - Superficial spreading melanoma|8743/3
C0334438|T191|AB|X78TC|RCD|SSMM-Superfic spread MM skin|8743/3
C0334438|T191|AB|X78TC|RCD|Superfic spread melanoma skin|8743/3
C0334438|T191|PT|X78TC|RCD|Superficial spreading malignant melanoma of skin|8743/3
C0334438|T191|PT|BBEH.|RCD|Superficial spreading melanoma|8743/3
C0334438|T191|SY|X78TC|RCD|Superficial spreading melanoma of skin|8743/3
C0334438|T191|AB|X78TC|RCD|Superficial spreading MM skin|8743/3
C0334438|T191|SY|254730000|SNOMEDCT_US|SMM - Superficial spreading melanoma of skin|8743/3
C0334438|T191|SY|55320002|SNOMEDCT_US|SSM - Superficial spreading melanoma|8743/3
C0334438|T191|SY|254730000|SNOMEDCT_US|SSMM - Superficial spreading malignant melanoma of skin|8743/3
C0334438|T191|SY|55320002|SNOMEDCT_US|SSMM - Superficial spreading melanoma|8743/3
C0334438|T191|PT|254730000|SNOMEDCT_US|Superficial spreading malignant melanoma of skin|8743/3
C0334438|T191|PT|55320002|SNOMEDCT_US|Superficial spreading melanoma|8743/3
C0334438|T191|SY|254730000|SNOMEDCT_US|Superficial spreading melanoma of skin|8743/3
C0346037|T191|PT|0000048913|CHV|acral lentiginous melanoma|8744/3
C0346037|T191|PT|HP:0012060|HPO|Acral lentiginous melanoma|8744/3
C0346037|T191|LA|LA27886-3|LNC|Acral lentiginous melanoma|8744/3
C0346037|T191|LLT|10000583|MDR|Acral lentiginous melanoma|8744/3
C0346037|T191|PT|10000583|MDR|Acral lentiginous melanoma|8744/3
C0346037|T191|PT|231654|MEDCIN|acral lentiginous melanoma of skin|8744/3
C0346037|T191|SY|231654|MEDCIN|malignant acral lentiginous melanoma|8744/3
C0346037|T191|PN|NOCODE|MTH|Acral Lentiginous Malignant Melanoma|8744/3
C0346037|T191|SY|C4022|NCI|Acral Lentiginous Malignant Melanoma|8744/3
C0346037|T191|PT|C4022|NCI|Acral Lentiginous Melanoma|8744/3
C0346037|T191|SY|TCGA|NCI|Acral Lentiginous Melanoma|8744/3
C0346037|T191|DN|C4022|NCI_CTRP|Acral Lentiginous Melanoma|8744/3
C0346037|T191|PT|CDR0000039905|PDQ|acral lentiginous malignant melanoma|8744/3
C0346037|T191|SY|CDR0000039905|PDQ|Acral Lentiginous Melanoma|8744/3
C0346037|T191|SY|CDR0000039905|PDQ|malignant melanoma, acral lentiginous|8744/3
C0346037|T191|SY|CDR0000039905|PDQ|melanoma, acral lentiginous malignant|8744/3
C0346037|T191|AB|X78TE|RCD|Acral lentigin melanoma skin|8744/3
C0346037|T191|PT|X78TE|RCD|Acral lentiginous malignant melanoma of skin|8744/3
C0346037|T191|SY|X78TE|RCD|Acral lentiginous melanoma of skin|8744/3
C0346037|T191|AB|X78TE|RCD|Acral lentiginous MM of skin|8744/3
C0346037|T191|SY|X78TE|RCD|ALM - Acral lentiginous melanoma of skin|8744/3
C0346037|T191|AB|X78TE|RCD|ALM-Acral lentig melanoma skin|8744/3
C0346037|T191|SY|X78TE|RCD|ALMM - Acral lentiginous malignant melanoma of skin|8744/3
C0346037|T191|AB|X78TE|RCD|ALMM-Acral lentiginous MM skin|8744/3
C0346037|T191|AB|X77oK|RCD|Malig acral lentigin melanoma|8744/3
C0346037|T191|PT|X77oK|RCD|Malignant acral lentiginous melanoma|8744/3
C0346037|T191|AB|X77oK|RCDSY|Acral lentig melanoma,malig|8744/3
C0346037|T191|SY|X77oK|RCDSY|Acral lentiginous melanoma, malignant|8744/3
C0346037|T191|PT|254732008|SNOMEDCT_US|Acral lentiginous malignant melanoma of skin|8744/3
C0346037|T191|SY|254732008|SNOMEDCT_US|Acral lentiginous melanoma of skin|8744/3
C0346037|T191|PT|16974005|SNOMEDCT_US|Acral lentiginous melanoma, malignant|8744/3
C0346037|T191|SY|254732008|SNOMEDCT_US|ALM - Acral lentiginous melanoma of skin|8744/3
C0346037|T191|SY|254732008|SNOMEDCT_US|ALMM - Acral lentiginous malignant melanoma of skin|8744/3
C0346037|T191|OAP|189755003|SNOMEDCT_US|Malignant acral lentiginous melanoma|8744/3
C0346037|T191|OF|189755003|SNOMEDCT_US|Malignant acral lentiginous melanoma|8744/3
C1333280|T191|LPN|LP344944-6|LNC|Desmoplastic melanoma|8745/3
C1333280|T191|CN|MTHU062818|LNC|Desmoplastic melanoma|8745/3
C1333280|T191|PT|10072449|MDR|Desmoplastic melanoma|8745/3
C1333280|T191|LLT|10072449|MDR|Desmoplastic melanoma|8745/3
C0334439|T191|PT|352917|MEDCIN|Desmoplastic malignant melanoma|8745/3
C0334439|T191|SY|352917|MEDCIN|malignant neoplasm melanoma desmoplastic|8745/3
C1275203|T191|SY|352920|MEDCIN|malignant neoplasm melanoma neurotrophic|8745/3
C1275203|T191|PT|352920|MEDCIN|neurotrophic malignant melanoma|8745/3
C0334439|T191|PN|NOCODE|MTH|Malignant desmoplastic melanoma|8745/3
C1275203|T191|PN|NOCODE|MTH|Neurotropic malignant melanoma|8745/3
C1333280|T191|PT|C37257|NCI|Desmoplastic Melanoma|8745/3
C1333280|T191|SY|TCGA|NCI|Desmoplastic Melanoma|8745/3
C1333280|T191|PT|CDR0000321367|NCI_NCI-GLOSS|desmoplastic melanoma|8745/3
C0334439|T191|AB|X77oL|RCD|Malign desmoplastic melanoma|8745/3
C0334439|T191|PT|X77oL|RCD|Malignant desmoplastic melanoma|8745/3
C1275203|T191|SY|X77oL|RCD|Malignant neurotropic melanoma|8745/3
C0334439|T191|AB|X77oL|RCDSY|Desmoplas melanom,malignant|8745/3
C0334439|T191|SY|X77oL|RCDSY|Desmoplastic melanoma, malignant|8745/3
C0334439|T191|PT|403924008|SNOMEDCT_US|Desmoplastic malignant melanoma|8745/3
C0334439|T191|SY|51757004|SNOMEDCT_US|Desmoplastic melanoma, amelanotic|8745/3
C0334439|T191|PT|51757004|SNOMEDCT_US|Desmoplastic melanoma, malignant|8745/3
C0334439|T191|OAP|189751007|SNOMEDCT_US|Malignant desmoplastic melanoma|8745/3
C0334439|T191|OF|189751007|SNOMEDCT_US|Malignant desmoplastic melanoma|8745/3
C1275203|T191|SY|399644007|SNOMEDCT_US|Malignant neurotropic melanoma|8745/3
C1275203|T191|SY|51757004|SNOMEDCT_US|Malignant neurotropic melanoma|8745/3
C1275203|T191|PT|403925009|SNOMEDCT_US|Neurotropic malignant melanoma|8745/3
C1275203|T191|PT|399644007|SNOMEDCT_US|Neurotropic melanoma, malignant|8745/3
C1275203|T191|SY|51757004|SNOMEDCT_US|Neurotropic melanoma, malignant|8745/3
C1266115|T191|LA|LA27887-1|LNC|Mucosal-lentiginous melanoma|8746/3
C1266115|T191|PT|231656|MEDCIN|mucosal lentiginous melanoma|8746/3
C1266115|T191|SY|C48622|NCI|Mucosal Lentiginous Malignant Melanoma|8746/3
C1266115|T191|SY|TCGA|NCI|Mucosal Lentiginous Melanoma|8746/3
C1266115|T191|PT|C48622|NCI|Mucosal Lentiginous Melanoma|8746/3
C1266115|T191|PT|128732001|SNOMEDCT_US|Mucosal lentiginous melanoma|8746/3
C0206737|T191|SY|0000021060|CHV|dermal nevus|8750/0
C0206737|T191|SY|0000021060|CHV|intradermal melanocytic nevus|8750/0
C0206737|T191|SY|0000021060|CHV|intradermal naevus|8750/0
C0206737|T191|SY|0000021060|CHV|intradermal nevi|8750/0
C0206737|T191|PT|0000021060|CHV|intradermal nevus|8750/0
C0206737|T191|PT|NOCODE|COSTAR|Dermal Nevus|8750/0
C0206737|T191|PTN|S82016|ICPC2P|intradermal naevus|8750/0
C0206737|T191|MTH_PTN|S82016|ICPC2P|intradermal nevus|8750/0
C0206737|T191|PT|S82016|ICPC2P|Naevus;intradermal|8750/0
C0206737|T191|MTH_PT|S82016|ICPC2P|Nevus;intradermal|8750/0
C0206737|T191|LLT|10049663|MDR|Intradermal naevus|8750/0
C0206737|T191|LLT|10058537|MDR|Intradermal nevus|8750/0
C0206737|T191|PM|D018330|MSH|Intradermal Nevi|8750/0
C0206737|T191|PM|D018330|MSH|Intradermal Nevus|8750/0
C0206737|T191|ET|D018330|MSH|Nevi, Intradermal|8750/0
C0206737|T191|MH|D018330|MSH|Nevus, Intradermal|8750/0
C0206737|T191|SY|C3804|NCI|Dermal Nevus|8750/0
C0206737|T191|PT|C3804|NCI|Intradermal Nevus|8750/0
C0206737|T191|SY|Xa99Z|RCD|Cellular naevus|8750/0
C0206737|T191|PT|Xa99Z|RCD|Dermal cellular naevus|8750/0
C0206737|T191|SY|Xa99Z|RCD|Dermal naevus|8750/0
C0206737|T191|SY|Xa99Z|RCD|IDN - Intradermal naevus|8750/0
C0206737|T191|SY|Xa99Z|RCD|Intradermal melanocytic naevus|8750/0
C0206737|T191|OP|BBEJ.|RCD|Intradermal naevus|8750/0
C0206737|T191|SY|Xa99Z|RCDAE|Cellular nevus|8750/0
C0206737|T191|PT|Xa99Z|RCDAE|Dermal cellular nevus|8750/0
C0206737|T191|SY|Xa99Z|RCDAE|Dermal nevus|8750/0
C0206737|T191|SY|Xa99Z|RCDAE|IDN - Intradermal nevus|8750/0
C0206737|T191|SY|Xa99Z|RCDAE|Intradermal melanocytic nevus|8750/0
C0206737|T191|OP|BBEJ.|RCDAE|Intradermal nevus|8750/0
C0206737|T191|SYGB|302838006|SNOMEDCT_US|Cellular naevus|8750/0
C0206737|T191|SY|302838006|SNOMEDCT_US|Cellular nevus|8750/0
C0206737|T191|PTGB|302838006|SNOMEDCT_US|Dermal cellular naevus|8750/0
C0206737|T191|PT|302838006|SNOMEDCT_US|Dermal cellular nevus|8750/0
C0206737|T191|SYGB|302838006|SNOMEDCT_US|Dermal naevus|8750/0
C0206737|T191|SYGB|112681002|SNOMEDCT_US|Dermal naevus|8750/0
C0206737|T191|SY|302838006|SNOMEDCT_US|Dermal nevus|8750/0
C0206737|T191|SY|112681002|SNOMEDCT_US|Dermal nevus|8750/0
C0206737|T191|SYGB|302838006|SNOMEDCT_US|IDN - Intradermal naevus|8750/0
C0206737|T191|SY|302838006|SNOMEDCT_US|IDN - Intradermal nevus|8750/0
C0206737|T191|SYGB|302838006|SNOMEDCT_US|Intradermal melanocytic naevus|8750/0
C0206737|T191|SY|302838006|SNOMEDCT_US|Intradermal melanocytic nevus|8750/0
C0206737|T191|PTGB|112681002|SNOMEDCT_US|Intradermal naevus|8750/0
C0206737|T191|PT|112681002|SNOMEDCT_US|Intradermal nevus|8750/0
C0259781|T191|SY|0000025232|CHV|compound naevus|8760/0
C0259781|T191|PT|0000025232|CHV|compound nevus|8760/0
C0259781|T191|SY|0000025232|CHV|nevus compound|8760/0
C0259781|T191|PT|U000194|COSTAR|COMPOUND NEVUS|8760/0
C0259781|T191|PTN|S82013|ICPC2P|compound naevus|8760/0
C0259781|T191|MTH_PTN|S82013|ICPC2P|compound nevus|8760/0
C0259781|T191|PT|S82013|ICPC2P|Naevus;compound|8760/0
C0259781|T191|MTH_PT|S82013|ICPC2P|Nevus;compound|8760/0
C0259781|T191|LLT|10058171|MDR|Compound naevus|8760/0
C0259781|T191|LLT|10058131|MDR|Compound nevus|8760/0
C0259781|T191|PT|214041|MEDCIN|compound nevus|8760/0
C0259781|T191|PT|C3901|NCI|Compound Nevus|8760/0
C0259781|T191|SY|C3901|NCI|Compound Nevus of Skin|8760/0
C0259781|T191|SY|C3901|NCI|Compound Nevus of the Skin|8760/0
C0259781|T191|PT|CDR0000044274|NCI_NCI-GLOSS|compound nevus|8760/0
C0259781|T191|PT|BBEK.|RCD|Compound naevus|8760/0
C0259781|T191|PT|X78V0|RCD|Compound naevus of skin|8760/0
C0259781|T191|SY|BBEK.|RCD|Dermal and epidermal naevus|8760/0
C0259781|T191|PT|BBEK.|RCDAE|Compound nevus|8760/0
C0259781|T191|PT|X78V0|RCDAE|Compound nevus of skin|8760/0
C0259781|T191|SY|BBEK.|RCDAE|Dermal and epidermal nevus|8760/0
C1302809|T047|PTGB|787085004|SNOMEDCT_US|Acantholytic epidermal naevus|8760/0
C1302809|T047|PTGB|400067002|SNOMEDCT_US|Acantholytic epidermal naevus|8760/0
C1302809|T047|PT|787085004|SNOMEDCT_US|Acantholytic epidermal nevus|8760/0
C1302809|T047|PT|400067002|SNOMEDCT_US|Acantholytic epidermal nevus|8760/0
C0259781|T191|PTGB|49409001|SNOMEDCT_US|Compound naevus|8760/0
C0259781|T191|PTGB|254805008|SNOMEDCT_US|Compound naevus of skin|8760/0
C0259781|T191|PT|49409001|SNOMEDCT_US|Compound nevus|8760/0
C0259781|T191|PT|254805008|SNOMEDCT_US|Compound nevus of skin|8760/0
C0259781|T191|SYGB|49409001|SNOMEDCT_US|Dermal and epidermal naevus|8760/0
C0259781|T191|SY|49409001|SNOMEDCT_US|Dermal and epidermal nevus|8760/0
C1302848|T191|PTGB|787086003|SNOMEDCT_US|Epidermolytic epidermal naevus|8760/0
C1302848|T191|PTGB|400142003|SNOMEDCT_US|Epidermolytic epidermal naevus|8760/0
C1302848|T191|PT|787086003|SNOMEDCT_US|Epidermolytic epidermal nevus|8760/0
C1302848|T191|PT|400142003|SNOMEDCT_US|Epidermolytic epidermal nevus|8760/0
C1302879|T191|PTGB|787087007|SNOMEDCT_US|Inflammatory epidermal naevus|8760/0
C1302879|T191|PTGB|400197008|SNOMEDCT_US|Inflammatory epidermal naevus|8760/0
C1302879|T191|PT|787087007|SNOMEDCT_US|Inflammatory epidermal nevus|8760/0
C1302879|T191|PT|400197008|SNOMEDCT_US|Inflammatory epidermal nevus|8760/0
C1883045|T191|PT|C66754|NCI|Small Congenital Melanocytic Nevus|8761/0
C1266116|T191|OAP|128881008|SNOMEDCT_US|Small congenital naevus|8761/0
C1266116|T191|OAP|128881008|SNOMEDCT_US|Small congenital nevus|8761/0
C1842036|T191|PT|0000029981|CHV|bathing trunk nevus|8761/1
C1842036|T191|SY|0000029981|CHV|congenital giant naevus pigmented|8761/1
C1842036|T191|SY|0000029981|CHV|congenital giant pigmented nevus|8761/1
C1842036|T191|SY|0000029981|CHV|nevus pigmented congenital giant|8761/1
C1842036|T191|PT|HP:0005600|HPO|Congenital giant melanocytic nevus|8761/1
C1842036|T191|SY|HP:0005600|HPO|Giant pigmented hairy nevus|8761/1
C1842036|T191|SY|HP:0005600|HPO|Giant pigmented mole|8761/1
C1842036|T191|SY|HP:0005600|HPO|Giant pigmented nevus|8761/1
C1842036|T191|PT|MTHU084210|ICPC2ICD10ENG|bathing trunk; nevus|8761/1
C1842036|T191|PT|MTHU051611|ICPC2ICD10ENG|nevus; bathing trunk|8761/1
C1842036|T191|CE|C536819|MSH|Giant congenital pigmented nevus|8761/1
C1842036|T191|CE|C536819|MSH|Giant pigmented hairy nevus|8761/1
C1842036|T191|NM|C536819|MSH|Melanocytic nevus syndrome, congenital|8761/1
C1842036|T191|PN|NOCODE|MTH|GIANT PIGMENTED HAIRY NEVUS|8761/1
C1842036|T191|SY|C4234|NCI|Bathing Trunk Nevus|8761/1
C1842036|T191|PT|C4234|NCI|Giant Congenital Nevus|8761/1
C1842036|T191|SY|C4234|NCI|Giant Pigmented Nevus of Skin|8761/1
C1842036|T191|SY|C4234|NCI|Giant Pigmented Nevus of the Skin|8761/1
C1842036|T191|SY|BBEL.|RCD|Bathing trunk naevus|8761/1
C1842036|T191|SY|X78VD|RCD|Bathing trunk naevus|8761/1
C1842036|T191|AB|BBEL.|RCD|Cong giant pigmented naevus|8761/1
C1842036|T191|AB|X78VD|RCD|Congen giant pigme naevus skin|8761/1
C1842036|T191|SY|BBEL.|RCD|Congenital giant pigmented naevus|8761/1
C1842036|T191|PT|X78VD|RCD|Congenital giant pigmented naevus of skin|8761/1
C1842036|T191|PT|BBEL.|RCD|Giant pigmented naevus|8761/1
C1842036|T191|SY|X78VD|RCD|Giant pigmented naevus of skin|8761/1
C1842036|T191|SY|X78VD|RCDAE|Bathing trunk nevus|8761/1
C1842036|T191|SY|BBEL.|RCDAE|Bathing trunk nevus|8761/1
C1842036|T191|AB|BBEL.|RCDAE|Cong giant pigmented nevus|8761/1
C1842036|T191|AB|X78VD|RCDAE|Congen giant pigme nevus skin|8761/1
C1842036|T191|SY|BBEL.|RCDAE|Congenital giant pigmented nevus|8761/1
C1842036|T191|PT|X78VD|RCDAE|Congenital giant pigmented nevus of skin|8761/1
C1842036|T191|PT|BBEL.|RCDAE|Giant pigmented nevus|8761/1
C1842036|T191|SY|X78VD|RCDAE|Giant pigmented nevus of skin|8761/1
C1842036|T191|SYGB|254815002|SNOMEDCT_US|Bathing trunk naevus|8761/1
C1842036|T191|SY|254815002|SNOMEDCT_US|Bathing trunk nevus|8761/1
C1842036|T191|SYGB|10291008|SNOMEDCT_US|Congenital giant pigmented naevus|8761/1
C1842036|T191|PTGB|254815002|SNOMEDCT_US|Congenital giant pigmented naevus of skin|8761/1
C1842036|T191|SY|10291008|SNOMEDCT_US|Congenital giant pigmented nevus|8761/1
C1842036|T191|PT|254815002|SNOMEDCT_US|Congenital giant pigmented nevus of skin|8761/1
C1842036|T191|PTGB|10291008|SNOMEDCT_US|Giant pigmented naevus|8761/1
C1842036|T191|SYGB|254815002|SNOMEDCT_US|Giant pigmented naevus of skin|8761/1
C1842036|T191|PT|10291008|SNOMEDCT_US|Giant pigmented nevus|8761/1
C1842036|T191|SY|254815002|SNOMEDCT_US|Giant pigmented nevus of skin|8761/1
C1842036|T191|IS|10291008|SNOMEDCT_US|Giant pigmented nevus, NOS|8761/1
C1842036|T191|SYGB|10291008|SNOMEDCT_US|Intermediate and giant congenital naevus|8761/1
C1842036|T191|SY|10291008|SNOMEDCT_US|Intermediate and giant congenital nevus|8761/1
C1883039|T191|PT|C4235|NCI|Melanoma Arising in Giant Congenital Nevus|8761/3
C0334441|T191|PT|BBEM.|RCD|Malignant melanoma in giant pigmented naevus|8761/3
C0334441|T191|AB|BBEM.|RCD|MM in giant pigmented naevus|8761/3
C0334441|T191|PT|BBEM.|RCDAE|Malignant melanoma in giant pigmented nevus|8761/3
C0334441|T191|AB|BBEM.|RCDAE|MM in giant pigmented nevus|8761/3
C0334441|T191|SYGB|75931002|SNOMEDCT_US|Malignant melanoma in congenital melanocytic naevus|8761/3
C0334441|T191|SY|75931002|SNOMEDCT_US|Malignant melanoma in congenital melanocytic nevus|8761/3
C0334441|T191|PTGB|75931002|SNOMEDCT_US|Malignant melanoma in giant pigmented naevus|8761/3
C0334441|T191|PT|75931002|SNOMEDCT_US|Malignant melanoma in giant pigmented nevus|8761/3
C1266117|T191|PT|C66755|NCI|Proliferative Dermal Lesion in Congenital Nevus|8762/1
C1266117|T191|PTGB|128733006|SNOMEDCT_US|Proliferative dermal lesion in congenital naevus|8762/1
C1266117|T191|PT|128733006|SNOMEDCT_US|Proliferative dermal lesion in congenital nevus|8762/1
C0206739|T191|SY|0000021062|CHV|benign juvenile melanoma|8770/0
C0206739|T191|SY|0000021062|CHV|juvenile melanoma|8770/0
C0206739|T191|SY|0000021062|CHV|naevus spitz|8770/0
C0206739|T191|SY|0000021062|CHV|nevus spitz|8770/0
C0206739|T191|SY|0000021062|CHV|spitz naevus|8770/0
C0206739|T191|PT|0000021062|CHV|spitz nevus|8770/0
C0206739|T191|LLT|10023255|MDR|Juvenile melanoma|8770/0
C0206739|T191|LLT|10023256|MDR|Juvenile melanoma benign|8770/0
C0206739|T191|PT|10023256|MDR|Juvenile melanoma benign|8770/0
C0206739|T191|LLT|10041632|MDR|Spitz naevus|8770/0
C0206739|T191|LLT|10062802|MDR|Spitz nevus|8770/0
C0206739|T191|MH|D018332|MSH|Nevus, Epithelioid and Spindle Cell|8770/0
C0206739|T191|ET|D018332|MSH|Nevus, Spindle Cell and Epithelioid|8770/0
C0206739|T191|PM|D018332|MSH|Nevus, Spitz|8770/0
C0206739|T191|ET|D018332|MSH|Spitz Nevus|8770/0
C0206739|T191|PN|NOCODE|MTH|Epithelioid and spindle cell nevus|8770/0
C0206739|T191|SY|C27007|NCI|Benign Juvenile Melanoma|8770/0
C0206739|T191|SY|C27007|NCI|Juvenile Nevus|8770/0
C0206739|T191|SY|C27007|NCI|Spindle and/ or Epithelioid Cell Nevus|8770/0
C0206739|T191|PT|C27007|NCI|Spitz Nevus|8770/0
C0206739|T191|OP|X78V7|RCD|Epithelioid and spindle cell naevus|8770/0
C0206739|T191|OA|X78V7|RCD|Epithelioid+spindle cell naev|8770/0
C0206739|T191|IS|X78V7|RCD|Juvenile melanoma|8770/0
C0206739|T191|IS|X78V7|RCD|Juvenile naevus|8770/0
C0206739|T191|IS|X78V7|RCD|Spindle and epithelioid naevus|8770/0
C0206739|T191|IS|X78V7|RCD|Spitz naevus|8770/0
C0206739|T191|OP|X78V7|RCDAE|Epithelioid and spindle cell nevus|8770/0
C0206739|T191|IS|X78V7|RCDAE|Juvenile nevus|8770/0
C0206739|T191|IS|X78V7|RCDAE|Spindle and epithelioid nevus|8770/0
C0206739|T191|IS|X78V7|RCDAE|Spitz nevus|8770/0
C0206739|T191|PT|BBEN.|RCDSA|Epithelioid and spindle cell nevus|8770/0
C0206739|T191|SY|BBEN.|RCDSA|Juvenila nevus|8770/0
C0206739|T191|SY|BBEN.|RCDSA|Spitz nevus|8770/0
C0206739|T191|AB|BBEN.|RCDSY|Epithel.+spindle cell naev.|8770/0
C0206739|T191|PT|BBEN.|RCDSY|Epithelioid and spindle cell naevus|8770/0
C0206739|T191|SY|BBEN.|RCDSY|Juvenila melanoma|8770/0
C0206739|T191|SY|BBEN.|RCDSY|Juvenila naevus|8770/0
C0206739|T191|SY|BBEN.|RCDSY|Spitz naevus|8770/0
C0206739|T191|PTGB|88082008|SNOMEDCT_US|Epithelioid and spindle cell naevus|8770/0
C0206739|T191|PTGB|254811006|SNOMEDCT_US|Epithelioid and spindle cell naevus|8770/0
C0206739|T191|PT|88082008|SNOMEDCT_US|Epithelioid and spindle cell nevus|8770/0
C0206739|T191|PT|254811006|SNOMEDCT_US|Epithelioid and spindle cell nevus|8770/0
C0206739|T191|SY|88082008|SNOMEDCT_US|Juvenila melanoma|8770/0
C0206739|T191|SY|88082008|SNOMEDCT_US|Juvenila nevus|8770/0
C0206739|T191|SY|88082008|SNOMEDCT_US|Juvenile melanoma|8770/0
C0206739|T191|SY|254811006|SNOMEDCT_US|Juvenile melanoma|8770/0
C0206739|T191|SYGB|88082008|SNOMEDCT_US|Juvenile naevus|8770/0
C0206739|T191|SYGB|254811006|SNOMEDCT_US|Juvenile naevus|8770/0
C0206739|T191|SY|88082008|SNOMEDCT_US|Juvenile nevus|8770/0
C0206739|T191|SY|254811006|SNOMEDCT_US|Juvenile nevus|8770/0
C0206739|T191|SYGB|88082008|SNOMEDCT_US|Pigmented spindle cell naevus of Reed|8770/0
C0206739|T191|SY|88082008|SNOMEDCT_US|Pigmented spindle cell nevus of Reed|8770/0
C0206739|T191|SYGB|254811006|SNOMEDCT_US|Spindle and epithelioid naevus|8770/0
C0206739|T191|SY|254811006|SNOMEDCT_US|Spindle and epithelioid nevus|8770/0
C0206739|T191|SYGB|254811006|SNOMEDCT_US|Spitz naevus|8770/0
C0206739|T191|SYGB|88082008|SNOMEDCT_US|Spitz naevus|8770/0
C0206739|T191|SY|254811006|SNOMEDCT_US|Spitz nevus|8770/0
C0206739|T191|SY|88082008|SNOMEDCT_US|Spitz nevus|8770/0
C0334442|T191|PT|C66756|NCI|Mixed Epithelioid and Spindle Cell Melanoma|8770/3
C0334442|T191|PT|C66756|NCI_CPTAC|Mixed Epithelioid and Spindle Cell Melanoma|8770/3
C0334442|T191|AB|BBET.|RCD|Mix epith+spindl cell melanoma|8770/3
C0334442|T191|PT|BBET.|RCD|Mixed epithelioid and spindle cell melanoma|8770/3
C0334442|T191|PT|50813003|SNOMEDCT_US|Mixed epithelioid and spindle cell melanoma|8770/3
C0259820|T191|PT|C66757|NCI|Epithelioid Cell Nevus|8771/0
C0259820|T191|PT|X77oQ|RCD|Epithelioid cell naevus|8771/0
C0259820|T191|PT|X77oQ|RCDAE|Epithelioid cell nevus|8771/0
C0259820|T191|OF|189760004|SNOMEDCT_US|Epithelioid cell naevus|8771/0
C0259820|T191|PTGB|11099005|SNOMEDCT_US|Epithelioid cell naevus|8771/0
C0259820|T191|OAP|189760004|SNOMEDCT_US|Epithelioid cell naevus|8771/0
C0259820|T191|OAP|189760004|SNOMEDCT_US|Epithelioid cell nevus|8771/0
C0259820|T191|PT|11099005|SNOMEDCT_US|Epithelioid cell nevus|8771/0
C0334443|T191|PN|NOCODE|MTH|Epithelioid Cell Melanoma|8771/3
C0334443|T191|SY|C4236|NCI|Epithelioid Cell Malignant Melanoma|8771/3
C0334443|T191|PT|C4236|NCI|Epithelioid Cell Melanoma|8771/3
C0334443|T191|SY|C4236|NCI|Epithelioid Melanoma|8771/3
C0334443|T191|PT|C4236|NCI_CPTAC|Epithelioid Cell Melanoma|8771/3
C0334443|T191|PT|BBEP.|RCD|Epithelioid cell melanoma|8771/3
C0334443|T191|PT|37138001|SNOMEDCT_US|Epithelioid cell melanoma|8771/3
C0206738|T191|PT|0000021061|CHV|spindle cell nevus|8772/0
C0206738|T191|ET|D018331|MSH|Nevi, Spindle Cell|8772/0
C0206738|T191|MH|D018331|MSH|Nevus, Spindle Cell|8772/0
C0206738|T191|PM|D018331|MSH|Spindle Cell Nevi|8772/0
C0206738|T191|PM|D018331|MSH|Spindle Cell Nevus|8772/0
C0206738|T191|PN|NOCODE|MTH|Nevus, Spindle Cell|8772/0
C0206738|T191|PT|C66758|NCI|Spindle Cell Nevus|8772/0
C0206738|T191|PT|X77oR|RCD|Spindle cell naevus|8772/0
C0206738|T191|PT|X77oR|RCDAE|Spindle cell nevus|8772/0
C0206738|T191|OP|BBEa.|RCDSA|Spindle cell nevus|8772/0
C0206738|T191|OP|BBEa.|RCDSY|Spindle cell naevus|8772/0
C0206738|T191|PTGB|810003|SNOMEDCT_US|Spindle cell naevus|8772/0
C0206738|T191|PTGB|253038006|SNOMEDCT_US|Spindle cell naevus|8772/0
C0206738|T191|PT|810003|SNOMEDCT_US|Spindle cell nevus|8772/0
C0206738|T191|PT|253038006|SNOMEDCT_US|Spindle cell nevus|8772/0
C0334444|T191|SY|352916|MEDCIN|malignant neoplasm melanoma spindle cell|8772/3
C0334444|T191|PT|352916|MEDCIN|Spindle cell malignant melanoma|8772/3
C0334444|T191|PN|NOCODE|MTH|Spindle Cell Melanoma|8772/3
C0334444|T191|SY|C4237|NCI|Malignant Spindle Cell Melanoma|8772/3
C0334444|T191|SY|C4237|NCI|Spindle Cell Malignant Melanoma|8772/3
C0334444|T191|PT|C4237|NCI|Spindle Cell Melanoma|8772/3
C0334444|T191|PT|C4237|NCI_CPTAC|Spindle Cell Melanoma|8772/3
C0334444|T191|PT|Xa99a|RCD|Spindle cell melanoma|8772/3
C0334444|T191|OP|BBEQ.|RCDSY|Spindle cell melanoma NOS|8772/3
C0334444|T191|PT|403923002|SNOMEDCT_US|Spindle cell malignant melanoma|8772/3
C0334444|T191|PT|68827007|SNOMEDCT_US|Spindle cell melanoma|8772/3
C0334444|T191|IS|68827007|SNOMEDCT_US|Spindle cell melanoma, NOS|8772/3
C0334444|T191|SY|68827007|SNOMEDCT_US|Spitzoid malignant melanoma|8772/3
C0334444|T191|SY|403923002|SNOMEDCT_US|Spitzoid malignant melanoma|8772/3
C0334445|T191|PT|MTHU048251|ICPC2ICD10ENG|melanoma; spindle cell type A|8773/3
C0334445|T191|PT|MTHU069004|ICPC2ICD10ENG|spindle cell; melanoma, type A|8773/3
C0334445|T191|SY|C4238|NCI|Malignant Spindle Cell Type A Melanoma|8773/3
C0334445|T191|SY|C4238|NCI|Spindle Cell Type A Malignant Melanoma|8773/3
C0334445|T191|PT|C4238|NCI|Type A Spindle Cell Melanoma|8773/3
C0334445|T191|PT|BBER.|RCD|Spindle cell melanoma - type A|8773/3
C0334445|T191|SY|24653009|SNOMEDCT_US|Spindle cell melanoma - type A|8773/3
C0334445|T191|PT|24653009|SNOMEDCT_US|Spindle cell melanoma, type A|8773/3
C0334446|T191|PT|MTHU048252|ICPC2ICD10ENG|melanoma; spindle cell type B|8774/3
C0334446|T191|PT|MTHU069005|ICPC2ICD10ENG|spindle cell; melanoma, type B|8774/3
C0334446|T191|SY|C4239|NCI|Malignant Spindle Cell Type B Melanoma|8774/3
C0334446|T191|SY|C4239|NCI|Spindle Cell Type B Malignant Melanoma|8774/3
C0334446|T191|PT|C4239|NCI|Type B Spindle Cell Melanoma|8774/3
C0334446|T191|PT|BBES.|RCD|Spindle cell melanoma - type B|8774/3
C0334446|T191|SY|40244008|SNOMEDCT_US|Spindle cell melanoma - type B|8774/3
C0334446|T191|PT|40244008|SNOMEDCT_US|Spindle cell melanoma, type B|8774/3
C0206736|T191|PT|0000021059|CHV|blue nevus|8780/0
C0206736|T191|SY|0000021059|CHV|nevus blue|8780/0
C0206736|T191|PT|U000011|COSTAR|BLUE NEVUS|8780/0
C0206736|T191|PT|MTHU012041|ICPC2ICD10ENG|blue nevus; Jadassohn|8780/0
C0206736|T191|PT|MTHU040526|ICPC2ICD10ENG|Jadassohn; blue nevus|8780/0
C0206736|T191|PTN|S82005|ICPC2P|blue naevus|8780/0
C0206736|T191|MTH_PTN|S82005|ICPC2P|blue nevus|8780/0
C0206736|T191|PT|S82005|ICPC2P|Naevus;blue|8780/0
C0206736|T191|MTH_PT|S82005|ICPC2P|Nevus;blue|8780/0
C0206736|T191|LLT|10005882|MDR|Blue naevus|8780/0
C0206736|T191|LLT|10062788|MDR|Blue nevus|8780/0
C0206736|T191|SY|277702|MEDCIN|benign blue nevus neoplasm|8780/0
C0206736|T191|PT|277702|MEDCIN|benign blue nevus of skin|8780/0
C0206736|T191|ET|D018329|MSH|Blue Nevi|8780/0
C0206736|T191|ET|D018329|MSH|Blue Nevus|8780/0
C0206736|T191|PM|D018329|MSH|Nevi, Blue|8780/0
C0206736|T191|MH|D018329|MSH|Nevus, Blue|8780/0
C0206736|T191|PN|NOCODE|MTH|Nevus, Blue|8780/0
C0206736|T191|PT|C3803|NCI|Blue Nevus|8780/0
C0206736|T191|SY|C3803|NCI|Blue Nevus of Skin|8780/0
C0206736|T191|SY|C3803|NCI|Blue Nevus of the Skin|8780/0
C0206736|T191|SY|C3803|NCI|Blue Skin Nevus|8780/0
C0206736|T191|PT|Xa99b|RCD|Blue naevus|8780/0
C0206736|T191|PT|X78V2|RCD|Blue naevus of skin|8780/0
C0206736|T191|SY|Xa99b|RCD|Jadassohn's blue naevus|8780/0
C0206736|T191|PT|Xa99b|RCDAE|Blue nevus|8780/0
C0206736|T191|PT|X78V2|RCDAE|Blue nevus of skin|8780/0
C0206736|T191|SY|Xa99b|RCDAE|Jadassohn's blue nevus|8780/0
C0206736|T191|OP|BBEU.|RCDSA|Blue nevus NOS|8780/0
C0206736|T191|OP|BBEU.|RCDSY|Blue naevus NOS|8780/0
C0206736|T191|OAS|189051001|SNOMEDCT_US|Blue naevus|8780/0
C0206736|T191|PTGB|63166000|SNOMEDCT_US|Blue naevus|8780/0
C0206736|T191|PTGB|254806009|SNOMEDCT_US|Blue naevus of skin|8780/0
C0206736|T191|OAS|189051001|SNOMEDCT_US|Blue nevus|8780/0
C0206736|T191|PT|63166000|SNOMEDCT_US|Blue nevus|8780/0
C0206736|T191|PT|254806009|SNOMEDCT_US|Blue nevus of skin|8780/0
C0206736|T191|IS|63166000|SNOMEDCT_US|Blue nevus, NOS|8780/0
C0206736|T191|SY|63166000|SNOMEDCT_US|Dermal melanocytoma|8780/0
C0206736|T191|SYGB|63166000|SNOMEDCT_US|Jadassohn's blue naevus|8780/0
C0206736|T191|SY|63166000|SNOMEDCT_US|Jadassohn's blue nevus|8780/0
C0334447|T191|LA|LA27889-7|LNC|Melanoma arising from blue nevus|8780/3
C0334447|T191|LLT|10072447|MDR|Blue naevus-like melanoma|8780/3
C0334447|T191|LLT|10072453|MDR|Blue nevus-like melanoma|8780/3
C0334447|T191|LLT|10072448|MDR|Malignant blue naevus|8780/3
C0334447|T191|PT|10072448|MDR|Malignant blue naevus|8780/3
C0334447|T191|LLT|10072455|MDR|Malignant blue nevus|8780/3
C0334447|T191|MTH_PT|10072448|MDR|Malignant blue nevus|8780/3
C0334447|T191|PT|231661|MEDCIN|malignant blue nevus of skin|8780/3
C0334447|T191|SY|C4240|NCI|Blue Nevus-Like Melanoma|8780/3
C0334447|T191|SY|C4240|NCI|Malignant Blue Nevus|8780/3
C0334447|T191|SY|C4240|NCI|Malignant Blue Nevus of Skin|8780/3
C0334447|T191|SY|C4240|NCI|Malignant Blue Nevus of the Skin|8780/3
C0334447|T191|SY|C4240|NCI|Malignant Cutaneous Blue Nevus|8780/3
C0334447|T191|SY|C4240|NCI|Malignant Skin Blue Nevus|8780/3
C0334447|T191|PT|C4240|NCI|Melanoma Arising from Blue Nevus|8780/3
C0334447|T191|SY|TCGA|NCI|Melanoma Arising from Blue Nevus|8780/3
C0334447|T191|SY|BBEV.|RCD|Malignant blue naevus|8780/3
C0334447|T191|PT|XaBAw|RCD|Malignant blue naevus of skin|8780/3
C0334447|T191|SY|BBEV.|RCDAE|Malignant blue nevus|8780/3
C0334447|T191|PT|XaBAw|RCDAE|Malignant blue nevus of skin|8780/3
C0334447|T191|PT|BBEV.|RCDSA|Blue nevus, malignant|8780/3
C0334447|T191|PT|BBEV.|RCDSY|Blue naevus, malignant|8780/3
C0334447|T191|PTGB|67159000|SNOMEDCT_US|Blue naevus, malignant|8780/3
C0334447|T191|PT|67159000|SNOMEDCT_US|Blue nevus, malignant|8780/3
C0334447|T191|SYGB|67159000|SNOMEDCT_US|Malignant blue naevus|8780/3
C0334447|T191|PTGB|307603002|SNOMEDCT_US|Malignant blue naevus of skin|8780/3
C0334447|T191|SY|67159000|SNOMEDCT_US|Malignant blue nevus|8780/3
C0334447|T191|PT|307603002|SNOMEDCT_US|Malignant blue nevus of skin|8780/3
C0334447|T191|SYGB|307603002|SNOMEDCT_US|Malignant melanoma in blue naevus|8780/3
C0334447|T191|SY|307603002|SNOMEDCT_US|Malignant melanoma in blue nevus|8780/3
C0334448|T191|PT|0000029982|CHV|cellular blue nevus|8790/0
C0334448|T191|PM|D018329|MSH|Blue Nevi, Cellular|8790/0
C0334448|T191|ET|D018329|MSH|Blue Nevus, Cellular|8790/0
C0334448|T191|ET|D018329|MSH|Cellular Blue Nevi|8790/0
C0334448|T191|PEP|D018329|MSH|Cellular Blue Nevus|8790/0
C0334448|T191|PM|D018329|MSH|Nevi, Cellular Blue|8790/0
C0334448|T191|PM|D018329|MSH|Nevus, Cellular Blue|8790/0
C0334448|T191|PT|C4241|NCI|Cellular Blue Nevus|8790/0
C0334448|T191|SY|C4241|NCI|Cellular Blue Nevus of Skin|8790/0
C0334448|T191|SY|C4241|NCI|Cellular Blue Nevus of the Skin|8790/0
C0334448|T191|PT|BBEW.|RCD|Cellular blue naevus|8790/0
C0334448|T191|PT|X78V4|RCD|Cellular blue naevus of skin|8790/0
C0334448|T191|PT|BBEW.|RCDAE|Cellular blue nevus|8790/0
C0334448|T191|PT|X78V4|RCDAE|Cellular blue nevus of skin|8790/0
C0334448|T191|PTGB|88006009|SNOMEDCT_US|Cellular blue naevus|8790/0
C0334448|T191|PTGB|254808005|SNOMEDCT_US|Cellular blue naevus of skin|8790/0
C0334448|T191|PT|88006009|SNOMEDCT_US|Cellular blue nevus|8790/0
C0334448|T191|PT|254808005|SNOMEDCT_US|Cellular blue nevus of skin|8790/0
C0334450|T191|PT|0037083|CCPSS|SOFT TISSUE TUMOR BENIGN|8800/0
C0334450|T191|PT|0000029983|CHV|benign neoplasm of soft tissue|8800/0
C0334450|T191|SY|0000029983|CHV|soft tissue benign tumor|8800/0
C0334450|T191|SY|0000029983|CHV|soft tissue tumor benign|8800/0
C0334450|T191|PTN|L97009|ICPC2P|benign neoplasm of the soft tissue|8800/0
C0334450|T191|OP|L71006|ICPC2P|Neoplasm benign;soft tissue|8800/0
C0334450|T191|PT|L97009|ICPC2P|Neoplasm benign;soft tissue|8800/0
C0334450|T191|LLT|10061004|MDR|Benign soft tissue neoplasm|8800/0
C0334450|T191|PT|10061004|MDR|Benign soft tissue neoplasm|8800/0
C0334450|T191|LLT|10004459|MDR|Benign soft tissue neoplasm NOS|8800/0
C0334450|T191|HG|10041294|MDR|Soft tissue neoplasms benign|8800/0
C0334450|T191|PT|333298|MEDCIN|benign soft tissue neoplasm|8800/0
C0334450|T191|SY|333298|MEDCIN|neoplasm - soft tissue benign|8800/0
C0334450|T191|SY|C4242|NCI|Benign Neoplasm of Soft Tissue|8800/0
C0334450|T191|SY|C4242|NCI|Benign Neoplasm of the Soft Tissue|8800/0
C0334450|T191|PT|C4242|NCI|Benign Soft Tissue Neoplasm|8800/0
C0334450|T191|SY|C4242|NCI|Benign Soft Tissue Tumor|8800/0
C0334450|T191|SY|C4242|NCI|Benign Tumor of Soft Tissue|8800/0
C0334450|T191|SY|C4242|NCI|Benign Tumor of the Soft Tissue|8800/0
C0334450|T191|PT|XM1FL|RCD|Benign soft tissue tumour|8800/0
C0334450|T191|PT|X78qp|RCD|Benign tumour of soft tissue|8800/0
C0334450|T191|OP|B75..|RCD|Other benign neoplasms of connective and soft tissue|8800/0
C0334450|T191|OA|B75..|RCD|Other soft tissue benign neop|8800/0
C0334450|T191|PT|XM1FL|RCDAE|Benign soft tissue tumor|8800/0
C0334450|T191|PT|X78qp|RCDAE|Benign tumor of soft tissue|8800/0
C0334450|T191|OP|BBF0.|RCDSA|Soft tissue tumor, benign|8800/0
C0334450|T191|OP|BBF0.|RCDSY|Soft tissue tumour, benign|8800/0
C0334450|T191|SY|92069005|SNOMEDCT_US|Benign neoplasm of connective and other soft tissues|8800/0
C0334450|T191|IS|92069005|SNOMEDCT_US|Benign neoplasm of connective and other soft tissues, NOS|8800/0
C0334450|T191|PT|92069005|SNOMEDCT_US|Benign neoplasm of soft tissue|8800/0
C0334450|T191|SY|92069005|SNOMEDCT_US|Benign neoplasm of soft tissues|8800/0
C0334450|T191|SY|47623001|SNOMEDCT_US|Benign soft tissue tumor|8800/0
C0334450|T191|SYGB|47623001|SNOMEDCT_US|Benign soft tissue tumour|8800/0
C0334450|T191|SY|92069005|SNOMEDCT_US|Benign tumor of soft tissue|8800/0
C0334450|T191|SYGB|92069005|SNOMEDCT_US|Benign tumour of soft tissue|8800/0
C0334450|T191|OAP|189019002|SNOMEDCT_US|Other benign neoplasms of connective and soft tissue|8800/0
C0334450|T191|PT|47623001|SNOMEDCT_US|Soft tissue tumor, benign|8800/0
C0334450|T191|PTGB|47623001|SNOMEDCT_US|Soft tissue tumour, benign|8800/0
C1261473|T191|DE|0000004530|AOD|sarcoma|8800/3
C1261473|T191|PT|0020102|CCPSS|SARCOMA|8800/3
C1261473|T191|SD|NEO024|CCSR_10|Sarcoma|8800/3
C1261473|T191|PT|U000602|COSTAR|SARCOMA|8800/3
C1261473|T191|PT|2000-8986|CSP|sarcoma|8800/3
C1261473|T191|PT|SARCOMA|CST|SARCOMA|8800/3
C1261473|T191|SY|HP:0100242|HPO|Cancer of connective tissue|8800/3
C1261473|T191|SY|HP:0100242|HPO|Malignant connective tissue tumor|8800/3
C1261473|T191|PT|HP:0100242|HPO|Sarcoma|8800/3
C1261473|T191|PT|A79013|ICPC2P|Sarcoma|8800/3
C1261473|T191|PTN|A79013|ICPC2P|sarcoma|8800/3
C1261473|T191|PT|U004213|LCH|Sarcoma|8800/3
C1261473|T191|PT|sh85117504|LCH_NW|Sarcoma|8800/3
C1261473|T191|LLT|10039491|MDR|Sarcoma|8800/3
C1261473|T191|PT|10039491|MDR|Sarcoma|8800/3
C1261473|T191|LLT|10039494|MDR|Sarcoma NOS|8800/3
C1261473|T191|PT|271492|MEDCIN|sarcoma|8800/3
C1261473|T191|MH|D012509|MSH|Sarcoma|8800/3
C1261473|T191|ET|D012509|MSH|Sarcoma, Soft Tissue|8800/3
C1261473|T191|PM|D012509|MSH|Sarcomas|8800/3
C1261473|T191|PM|D012509|MSH|Sarcomas, Soft Tissue|8800/3
C1261473|T191|PM|D012509|MSH|Soft Tissue Sarcoma|8800/3
C1261473|T191|PM|D012509|MSH|Soft Tissue Sarcomas|8800/3
C1261473|T191|PN|NOCODE|MTH|Sarcoma|8800/3
C1261473|T191|PT|C9118|NCI|Sarcoma|8800/3
C1261473|T191|SY|TCGA|NCI|Sarcoma|8800/3
C1261473|T191|SY|C9118|NCI|Sarcoma of Soft Tissue and Bone|8800/3
C1261473|T191|SY|C9118|NCI|Sarcoma of the Soft Tissue and Bone|8800/3
C1261473|T191|SY|C9118|NCI_CDISC|Mesenchymal Tumor, Malignant|8800/3
C1261473|T191|SY|C9118|NCI_CDISC|Sarcoma|8800/3
C1261473|T191|SY|C9118|NCI_CDISC|Sarcoma of Soft Tissue and Bone|8800/3
C1261473|T191|SY|C9118|NCI_CDISC|Sarcoma of the Soft Tissue and Bone|8800/3
C1261473|T191|PT|C9118|NCI_CDISC|SARCOMA, MALIGNANT|8800/3
C1261473|T191|PT|C9118|NCI_CPTAC|Sarcoma|8800/3
C1261473|T191|PT|C9118|NCI_CTRP|Sarcoma|8800/3
C1261473|T191|DN|C9118|NCI_CTRP|Sarcoma|8800/3
C1261473|T191|PT|CDR0000045562|NCI_NCI-GLOSS|sarcoma|8800/3
C1261473|T191|PT|C9118|NCI_NICHD|Sarcoma|8800/3
C1261473|T191|SY|CDR0000039253|PDQ|sarcoma|8800/3
C1261473|T191|SY|CDR0000039253|PDQ|Sarcoma of Soft Tissue and Bone|8800/3
C1261473|T191|SY|CDR0000039253|PDQ|Sarcoma of the Soft Tissue and Bone|8800/3
C1261473|T191|ET|45270|PSY|Sarcomas|8800/3
C1261473|T191|SY|Xa99e|RCD|Malignant mesenchymal tumour|8800/3
C1261473|T191|PT|Xa99e|RCD|Sarcoma|8800/3
C1261473|T191|SY|Xa99e|RCD|Soft tissue sarcoma|8800/3
C1261473|T191|SY|Xa99e|RCDAE|Malignant mesenchymal tumor|8800/3
C1261473|T191|OP|BBF1.|RCDSY|Sarcoma NOS|8800/3
C1261473|T191|SY|2424003|SNOMEDCT_US|Malignant mesenchymal tumor|8800/3
C1261473|T191|SYGB|2424003|SNOMEDCT_US|Malignant mesenchymal tumour|8800/3
C1261473|T191|SY|2424003|SNOMEDCT_US|Mesenchymal tumor, malignant|8800/3
C1261473|T191|SYGB|2424003|SNOMEDCT_US|Mesenchymal tumour, malignant|8800/3
C4041089|T191|PT|708979005|SNOMEDCT_US|Poorly differentiated sarcoma|8800/3
C4304633|T191|PT|719952009|SNOMEDCT_US|Primary sarcoma|8800/3
C1261473|T191|PT|424413001|SNOMEDCT_US|Sarcoma|8800/3
C1261473|T191|PT|2424003|SNOMEDCT_US|Sarcoma|8800/3
C1261473|T191|OAS|269634000|SNOMEDCT_US|Sarcoma NOS|8800/3
C1261473|T191|SY|2424003|SNOMEDCT_US|Sarcoma, no ICD-O subtype|8800/3
C1261473|T191|SY|2424003|SNOMEDCT_US|Sarcoma, no International Classification of Diseases for Oncology subtype|8800/3
C1261473|T191|IS|2424003|SNOMEDCT_US|Sarcoma, NOS|8800/3
C1261473|T191|PT|1047|WHO|SARCOMA|8800/3
C0748505|T191|PT|0025086|CCPSS|SARCOMA METASTATIC|8800/6
C0748505|T191|PT|10068595|MDR|Sarcoma metastatic|8800/6
C0748505|T191|LLT|10068595|MDR|Sarcoma metastatic|8800/6
C0748505|T191|PT|352268|MEDCIN|Metastatic sarcoma|8800/6
C0748505|T191|SY|352268|MEDCIN|sarcoma metastatic|8800/6
C0748505|T191|PT|C152076|NCI|Metastatic Sarcoma|8800/6
C0748505|T191|PT|C152076|NCI_CPTAC|Metastatic Sarcoma|8800/6
C0748505|T191|PT|443144000|SNOMEDCT_US|Metastatic sarcoma|8800/6
C0748505|T191|PT|372152003|SNOMEDCT_US|Sarcoma, metastatic|8800/6
C0334451|T191|LLT|10039500|MDR|Sarcomatosis|8800/9
C0334451|T191|PT|10039500|MDR|Sarcomatosis|8800/9
C0334451|T191|PT|C4243|NCI|Sarcomatosis|8800/9
C0334451|T191|PT|Xa99g|RCD|Sarcomatosis|8800/9
C0334451|T191|OP|BBF2.|RCDSY|Sarcomatosis NOS|8800/9
C0334451|T191|PT|9395006|SNOMEDCT_US|Sarcomatosis|8800/9
C0334451|T191|IS|9395006|SNOMEDCT_US|Sarcomatosis, NOS|8800/9
C0205945|T191|SY|0000020754|CHV|sarcoma spindle cell|8801/3
C0205945|T191|PT|0000020754|CHV|spindle cell sarcoma|8801/3
C0205945|T191|PT|MTHU065933|ICPC2ICD10ENG|sarcoma; spindle cell|8801/3
C0205945|T191|PT|MTHU069007|ICPC2ICD10ENG|spindle cell; sarcoma|8801/3
C0205945|T191|PT|10049067|MDR|Spindle cell sarcoma|8801/3
C0205945|T191|LLT|10049067|MDR|Spindle cell sarcoma|8801/3
C0205945|T191|PT|271493|MEDCIN|spindle cell sarcoma|8801/3
C0205945|T191|PEP|D012509|MSH|Sarcoma, Spindle Cell|8801/3
C0205945|T191|PM|D012509|MSH|Sarcomas, Spindle Cell|8801/3
C0205945|T191|PM|D012509|MSH|Spindle Cell Sarcoma|8801/3
C0205945|T191|PM|D012509|MSH|Spindle Cell Sarcomas|8801/3
C0205945|T191|PT|C27005|NCI|Spindle Cell Sarcoma|8801/3
C0205945|T191|PT|C27005|NCI_CPTAC|Spindle Cell Sarcoma|8801/3
C0205945|T191|PT|CDR0000044298|NCI_NCI-GLOSS|spindle cell sarcoma|8801/3
C0205945|T191|PT|BBF3.|RCD|Spindle cell sarcoma|8801/3
C0205945|T191|PT|9801004|SNOMEDCT_US|Spindle cell sarcoma|8801/3
C3839767|T191|PTGB|703606000|SNOMEDCT_US|Pleomorphic hyalinising angiectatic tumour|8802/1
C3839767|T191|PT|703606000|SNOMEDCT_US|Pleomorphic hyalinizing angiectatic tumor|8802/1
C1261358|T191|PT|271494|MEDCIN|giant cell sarcoma|8802/3
C1261358|T191|OP|C66759|NCI|Giant Cell Sarcoma|8802/3
C1261358|T191|PT|C66759|NCI|Giant Cell Sarcoma|8802/3
C1261358|T191|PT|Xa99h|RCD|Giant cell sarcoma|8802/3
C1261358|T191|SY|Xa99h|RCD|Pleomorphic cell sarcoma|8802/3
C0334452|T191|OA|BBF4.|RCDSY|Giant cell sarcoma-not bone|8802/3
C1261358|T191|PT|302840001|SNOMEDCT_US|Giant cell sarcoma|8802/3
C1261358|T191|SY|87992000|SNOMEDCT_US|Pleomorphic cell sarcoma|8802/3
C1261358|T191|SY|302840001|SNOMEDCT_US|Pleomorphic cell sarcoma|8802/3
C0334452|T191|SY|87992000|SNOMEDCT_US|Undifferentiated pleomorphic cell sarcoma|8802/3
C0553581|T191|PT|0000039090|CHV|round cell sarcoma|8803/3
C0206652|T191|PT|0000020996|CHV|small cell sarcoma|8803/3
C0553581|T191|PT|MTHU065046|ICPC2ICD10ENG|round cell; sarcoma|8803/3
C0553581|T191|PT|MTHU065931|ICPC2ICD10ENG|sarcoma; round cell|8803/3
C0206652|T191|PT|MTHU065916|ICPC2ICD10ENG|sarcoma; small cell|8803/3
C0206652|T191|PT|MTHU041514|ICPC2ICD10ENG|small cell; sarcoma|8803/3
C0206652|T191|PT|271495|MEDCIN|small cell sarcoma|8803/3
C0206652|T191|PM|D018228|MSH|Cell Sarcoma, Small|8803/3
C0206652|T191|PM|D018228|MSH|Cell Sarcomas, Small|8803/3
C0206652|T191|MH|D018228|MSH|Sarcoma, Small Cell|8803/3
C0206652|T191|PM|D018228|MSH|Sarcomas, Small Cell|8803/3
C0206652|T191|PM|D018228|MSH|Small Cell Sarcoma|8803/3
C0206652|T191|PM|D018228|MSH|Small Cell Sarcomas|8803/3
C0206652|T191|PT|C3746|NCI|Small Cell Sarcoma|8803/3
C0206652|T191|SY|C3746|NCI|Small Cell Sarcomas|8803/3
C0206652|T191|PT|C3746|NCI_CPTAC|Small Cell Sarcoma|8803/3
C0553581|T191|PT|X77oT|RCD|Round cell sarcoma|8803/3
C0206652|T191|PT|BBF5.|RCD|Small cell sarcoma|8803/3
C0553581|T191|SY|73506006|SNOMEDCT_US|Round cell sarcoma|8803/3
C0553581|T191|PT|253039003|SNOMEDCT_US|Round cell sarcoma|8803/3
C0206652|T191|PT|73506006|SNOMEDCT_US|Small cell sarcoma|8803/3
C0205944|T191|PT|MTHU026833|ICPC2ICD10ENG|epithelioid; sarcoma|8804/3
C0205944|T191|PT|MTHU065897|ICPC2ICD10ENG|sarcoma; epithelioid|8804/3
C0205944|T191|PT|10015099|MDR|Epithelioid sarcoma|8804/3
C0205944|T191|LLT|10015099|MDR|Epithelioid sarcoma|8804/3
C0205944|T191|LLT|10015103|MDR|Epithelioid sarcoma NOS|8804/3
C0205944|T191|HT|10015100|MDR|Epithelioid sarcomas|8804/3
C0205944|T191|PT|271496|MEDCIN|epithelioid sarcoma|8804/3
C0205944|T191|PM|D012509|MSH|Epithelioid Sarcoma|8804/3
C0205944|T191|PM|D012509|MSH|Epithelioid Sarcomas|8804/3
C0205944|T191|PEP|D012509|MSH|Sarcoma, Epithelioid|8804/3
C0205944|T191|PM|D012509|MSH|Sarcomas, Epithelioid|8804/3
C0205944|T191|PN|NOCODE|MTH|Sarcoma, Epithelioid|8804/3
C0205944|T191|SY|C3714|NCI|Epithelioid Cell Sarcoma|8804/3
C0205944|T191|PT|C3714|NCI|Epithelioid Sarcoma|8804/3
C0205944|T191|AB|C3714|NCI|ES|8804/3
C0205944|T191|SY|BBF6.|RCD|Epithelioid cell sarcoma|8804/3
C0205944|T191|PT|BBF6.|RCD|Epithelioid sarcoma|8804/3
C0205944|T191|SY|59238007|SNOMEDCT_US|Epithelioid cell sarcoma|8804/3
C0205944|T191|PT|782827000|SNOMEDCT_US|Epithelioid sarcoma|8804/3
C0205944|T191|PT|59238007|SNOMEDCT_US|Epithelioid sarcoma|8804/3
C0855073|T191|PT|0000050298|CHV|undifferentiated sarcoma|8805/3
C0855073|T191|PT|MTHU025481|ICPC2ICD10ENG|embryonal; sarcoma|8805/3
C0855073|T191|PT|MTHU065894|ICPC2ICD10ENG|sarcoma; embryonal|8805/3
C0855073|T191|LLT|10045515|MDR|Undifferentiated sarcoma|8805/3
C0855073|T191|PT|10045515|MDR|Undifferentiated sarcoma|8805/3
C0855073|T191|PT|271500|MEDCIN|embryonal sarcoma|8805/3
C0855073|T191|PT|271497|MEDCIN|undifferentiated sarcoma|8805/3
C0855073|T191|SY|C27096|NCI|Embryonal Sarcoma|8805/3
C0855073|T191|AB|C27096|NCI|UES|8805/3
C0855073|T191|SY|C27096|NCI|Undifferentiated Sarcoma|8805/3
C0855073|T191|SY|C27096|NCI_CDISC|Embryonal Sarcoma, Undifferentiated|8805/3
C0855073|T191|PT|C27096|NCI_CDISC|SARCOMA, UNDIFFERENTIATED, MALIGNANT|8805/3
C0855073|T191|PT|BBLD.|RCD|Embryonal sarcoma|8805/3
C0855073|T191|PT|59583009|SNOMEDCT_US|Embryonal sarcoma|8805/3
C0855073|T191|PT|128734000|SNOMEDCT_US|Undifferentiated sarcoma|8805/3
C0281508|T191|LLT|10064587|MDR|Desmoplastic small round cell tumor|8806/3
C0281508|T191|MTH_PT|10064581|MDR|Desmoplastic small round cell tumor|8806/3
C0281508|T191|LLT|10064581|MDR|Desmoplastic small round cell tumour|8806/3
C0281508|T191|PT|10064581|MDR|Desmoplastic small round cell tumour|8806/3
C0281508|T191|ET|D058405|MSH|Desmoplastic Small Cell Tumor|8806/3
C0281508|T191|MH|D058405|MSH|Desmoplastic Small Round Cell Tumor|8806/3
C0281508|T191|ET|D058405|MSH|Desmoplastic Small Round-Cell Tumor|8806/3
C0281508|T191|ET|D058405|MSH|Desmoplastic Small-Cell Tumor|8806/3
C0281508|T191|PM|D058405|MSH|Desmoplastic Small-Cell Tumors|8806/3
C0281508|T191|PM|D058405|MSH|Small-Cell Tumor, Desmoplastic|8806/3
C0281508|T191|PM|D058405|MSH|Small-Cell Tumors, Desmoplastic|8806/3
C0281508|T191|PM|D058405|MSH|Tumor, Desmoplastic Small-Cell|8806/3
C0281508|T191|PM|D058405|MSH|Tumors, Desmoplastic Small-Cell|8806/3
C0281508|T191|PN|NOCODE|MTH|Desmoplastic Small Round Cell Tumor|8806/3
C0281508|T191|PT|C8300|NCI|Desmoplastic Small Round Cell Tumor|8806/3
C0281508|T191|SY|C8300|NCI|Desmoplastic Small Round-Cell Neoplasm|8806/3
C0281508|T191|SY|C8300|NCI|Desmoplastic Small Round-Cell Tumor|8806/3
C0281508|T191|AB|C8300|NCI|DSRCT|8806/3
C0281508|T191|SY|C8300|NCI|Polyphenotypic Small Round Cell Tumor|8806/3
C0281508|T191|SY|10064587|NCI_CTEP-SDC|Desmoplas. small round cell tumor|8806/3
C0281508|T191|PT|10064587|NCI_CTEP-SDC|Desmoplastic small round cell tumor|8806/3
C0281508|T191|DN|C8300|NCI_CTRP|Desmoplastic Small Round Cell Tumor|8806/3
C0281508|T191|PT|CDR0000044495|NCI_NCI-GLOSS|desmoplastic small round cell tumor|8806/3
C0281508|T191|PT|128735004|SNOMEDCT_US|Desmoplastic small round cell tumor|8806/3
C0281508|T191|PTGB|128735004|SNOMEDCT_US|Desmoplastic small round cell tumour|8806/3
C0016045|T191|ET|0000004538|AOD|fibroma|8810/0
C0334067|T191|PT|0056523|CCPSS|BONE FIBROUS CORTICAL DEFECT|8810/0
C0016045|T191|PT|0011062|CCPSS|FIBROMA|8810/0
C0553647|T191|PT|0000039099|CHV|aponeurotic fibroma|8810/0
C0553647|T191|SY|0000039099|CHV|calcified fibroma|8810/0
C1300346|T191|PT|0000057622|CHV|collagenous fibroma|8810/0
C1300346|T191|SY|0000057622|CHV|desmoplastic fibroblastoma|8810/0
C0016045|T191|SY|0000005030|CHV|fibroma|8810/0
C0334067|T191|SY|0000029903|CHV|fibroma non ossifying|8810/0
C0016045|T191|SY|0000005030|CHV|fibromas|8810/0
C0334067|T191|SY|0000029903|CHV|fibromas non ossifying|8810/0
C0016045|T191|PT|0000005030|CHV|fibrous tissue tumor|8810/0
C0334067|T191|SY|0000029903|CHV|metaphyseal fibrous defect|8810/0
C0334067|T191|PT|0000029903|CHV|non-ossifying fibroma|8810/0
C0016045|T191|PT|2000-6014|CSP|fibroma|8810/0
C0016045|T191|PT|HP:0010614|HPO|Fibroma|8810/0
C0016045|T191|PT|S79001|ICPC2P|Fibroma|8810/0
C0016045|T191|PTN|S79001|ICPC2P|fibroma|8810/0
C0016045|T191|PT|U001784|LCH|Fibromas|8810/0
C0016045|T191|PT|sh85048035|LCH_NW|Fibromas|8810/0
C1300346|T191|LLT|10081841|MDR|Desmoplastic fibroblastoma|8810/0
C1300346|T191|PT|10081841|MDR|Desmoplastic fibroblastoma|8810/0
C0016045|T191|LLT|10016629|MDR|Fibroma|8810/0
C0016045|T191|PT|10016629|MDR|Fibroma|8810/0
C0016045|T191|LLT|10016630|MDR|Fibroma NOS|8810/0
C0334067|T191|LLT|10057717|MDR|Non-ossifying fibroma|8810/0
C0334067|T191|OL|10029649|MDR|Nonossifying fibroma|8810/0
C0016045|T191|LLT|10045154|MDR|Tumor of fibrous tissue NOS|8810/0
C0553647|T191|NM|C000625499|MSH|calcifying aponeurotic fibroma|8810/0
C0016045|T191|MH|D005350|MSH|Fibroma|8810/0
C0016045|T191|PM|D005350|MSH|Fibromas|8810/0
C1300346|T191|PN|NOCODE|MTH|Desmoplastic fibroblastoma|8810/0
C0016045|T191|PN|NOCODE|MTH|fibroma|8810/0
C1708187|T191|PN|NOCODE|MTH|Gardner Fibroma|8810/0
C0334067|T191|PN|NOCODE|MTH|Non-Ossifying Fibroma|8810/0
C1275237|T191|PN|NOCODE|MTH|Storiform collagenoma|8810/0
C0553647|T191|PT|C4818|NCI|Calcifying Aponeurotic Fibroma|8810/0
C1300346|T191|SY|C27515|NCI|Collagenous Fibroma|8810/0
C1708187|T191|SY|C49017|NCI|Desmoid Precursor Lesion|8810/0
C1300346|T191|PT|C27515|NCI|Desmoplastic Fibroblastoma|8810/0
C0016045|T191|PT|C3041|NCI|Fibroma|8810/0
C1708187|T191|PT|C49017|NCI|Gardner Fibroma|8810/0
C1708187|T191|SY|C49017|NCI|Gardner's Fibroma|8810/0
C0553647|T191|SY|C4818|NCI|Juvenile Aponeurotic Fibroma|8810/0
C0553647|T191|SY|C4818|NCI|Juvenile Aponeurotic Fibrosis|8810/0
C0334067|T191|AB|C121929|NCI|NOF|8810/0
C0334067|T191|PT|C121929|NCI|Non-Ossifying Fibroma|8810/0
C1532393|T191|SY|C6486|NCI|Nuchal Fibroma|8810/0
C1532393|T191|PT|C6486|NCI|Nuchal-Type Fibroma|8810/0
C1300346|T191|SY|C27515|NCI|Sclerotic Fibroma|8810/0
C1708187|T191|SY|C49017|NCI|Soft Fibroma|8810/0
C0016045|T191|PT|C3041|NCI_CDISC|FIBROMA, BENIGN|8810/0
C0553647|T191|SY|X50DL|RCD|Calcifying aponeurotic fibroma|8810/0
C0016045|T191|PT|Xa99j|RCD|Fibroma|8810/0
C0016045|T191|SY|Xa99j|RCD|Fibroma durum|8810/0
C0553647|T191|AB|X50DL|RCD|Juv palmo-plantar fibromatosis|8810/0
C0553647|T191|PT|X50DL|RCD|Juvenile aponeurotic fibroma|8810/0
C0553647|T191|SY|X50DL|RCD|Juvenile palmo-plantar fibromatosis|8810/0
C0016045|T191|OP|BBG0.|RCDSY|Fibroma NOS|8810/0
C0553647|T191|IS|133856002|SNOMEDCT_US|Aponeurotic fibroma|8810/0
C0553647|T191|OP|133856002|SNOMEDCT_US|Calcifying aponeurotic fibroma|8810/0
C0553647|T191|OP|238862009|SNOMEDCT_US|Calcifying aponeurotic fibroma|8810/0
C0553647|T191|PT|703612005|SNOMEDCT_US|Calcifying aponeurotic fibroma|8810/0
C0553647|T191|PT|703614006|SNOMEDCT_US|Calcifying aponeurotic fibroma|8810/0
C1300346|T191|SY|388984008|SNOMEDCT_US|Collagenous fibroma|8810/0
C1300346|T191|PT|388984008|SNOMEDCT_US|Desmoplastic fibroblastoma|8810/0
C0016045|T191|PT|424568000|SNOMEDCT_US|Fibroma|8810/0
C0016045|T191|OAS|154627003|SNOMEDCT_US|Fibroma|8810/0
C0016045|T191|OAS|269648000|SNOMEDCT_US|Fibroma|8810/0
C0016045|T191|PT|112682009|SNOMEDCT_US|Fibroma|8810/0
C0016045|T191|IS|112682009|SNOMEDCT_US|Fibroma durum|8810/0
C0016045|T191|SY|112682009|SNOMEDCT_US|Fibroma, no ICD-O subtype|8810/0
C0016045|T191|SY|112682009|SNOMEDCT_US|Fibroma, no International Classification of Diseases for Oncology subtype|8810/0
C0016045|T191|IS|112682009|SNOMEDCT_US|Fibroma, NOS|8810/0
C0334067|T191|SY|80415005|SNOMEDCT_US|Fibrous cortical defect of bone|8810/0
C1708187|T191|PT|703607009|SNOMEDCT_US|Gardner fibroma|8810/0
C0553647|T191|PT|238862009|SNOMEDCT_US|Juvenile aponeurotic fibroma|8810/0
C0553647|T191|PT|133856002|SNOMEDCT_US|Juvenile aponeurotic fibroma|8810/0
C0553647|T191|SY|238862009|SNOMEDCT_US|Juvenile palmo-plantar fibromatosis|8810/0
C0553647|T191|SY|133856002|SNOMEDCT_US|Keasbey tumor|8810/0
C0553647|T191|SYGB|133856002|SNOMEDCT_US|Keasbey tumour|8810/0
C0553647|T191|SY|133856002|SNOMEDCT_US|Keasbey's tumor|8810/0
C0553647|T191|SYGB|133856002|SNOMEDCT_US|Keasbey's tumour|8810/0
C0334067|T191|PT|80415005|SNOMEDCT_US|Metaphyseal fibrous defect|8810/0
C0334067|T191|SY|80415005|SNOMEDCT_US|Non-ossifying fibroma|8810/0
C1532393|T191|PT|403987004|SNOMEDCT_US|Nuchal fibroma|8810/0
C1532393|T191|SY|414881000|SNOMEDCT_US|Nuchal fibroma|8810/0
C1532393|T191|PT|414881000|SNOMEDCT_US|Nuchal-type fibroma|8810/0
C5230986|T191|PT|817948000|SNOMEDCT_US|Plaque-like CD34 positive dermal fibroma|8810/0
C1275237|T191|PT|709002005|SNOMEDCT_US|Sclerotic fibroma|8810/0
C1275237|T191|PT|403993007|SNOMEDCT_US|Storiform collagenoma|8810/0
C1275237|T191|SY|709002005|SNOMEDCT_US|Storiform collagenoma|8810/0
C1266118|T191|PT|C6892|NCI|Cellular Fibroma|8810/1
C1266118|T191|PT|128882001|SNOMEDCT_US|Cellular fibroma|8810/1
C0016057|T191|ET|0000004531|AOD|fibrosarcoma|8810/3
C0016057|T191|PT|0056525|CCPSS|FIBROSARCOMA|8810/3
C0016057|T191|PT|0000005036|CHV|fibrosarcoma|8810/3
C0016057|T191|SY|0000005036|CHV|fibrosarcomas|8810/3
C0016057|T191|PT|U000290|COSTAR|FIBROSARCOMA|8810/3
C0016057|T191|PT|2000-6227|CSP|fibrosarcoma|8810/3
C0016057|T191|DI|U000648|DXP|FIBROSARCOMA|8810/3
C0016057|T191|PT|HP:0100244|HPO|Fibrosarcoma|8810/3
C0016057|T191|PTN|L71017|ICPC2P|fibrosarcoma|8810/3
C0016057|T191|PT|L71017|ICPC2P|Fibrosarcoma|8810/3
C0016057|T191|LLT|10016632|MDR|Fibrosarcoma|8810/3
C0016057|T191|PT|10016632|MDR|Fibrosarcoma|8810/3
C0016057|T191|LLT|10016637|MDR|Fibrosarcoma NOS|8810/3
C0016057|T191|HT|10016634|MDR|Fibrosarcomas malignant|8810/3
C0016057|T191|PT|271507|MEDCIN|fibrosarcoma|8810/3
C0016057|T191|MH|D005354|MSH|Fibrosarcoma|8810/3
C0016057|T191|PM|D005354|MSH|Fibrosarcomas|8810/3
C0016057|T191|PN|NOCODE|MTH|Fibrosarcoma|8810/3
C0016057|T191|PT|C3043|NCI|Fibrosarcoma|8810/3
C0016057|T191|PT|C3043|NCI_CDISC|FIBROSARCOMA, MALIGNANT|8810/3
C0016057|T191|PT|C3043|NCI_CPTAC|Fibrosarcoma|8810/3
C0016057|T191|SY|10016637|NCI_CTEP-SDC|Fibrosarcoma - not infantile|8810/3
C0016057|T191|PT|CDR0000046403|NCI_NCI-GLOSS|fibrosarcoma|8810/3
C0016057|T191|PT|C3043|NCI_NICHD|Fibrosarcoma|8810/3
C0016057|T191|SY|C3043|NCI_NICHD|Malignant Fibromatous Neoplasm|8810/3
C0016057|T191|SY|BBG1.|RCD|Fibrosarcoma|8810/3
C0016057|T191|PT|BBG1.|RCDSY|Fibrosarcoma NOS|8810/3
C0016057|T191|SY|443250000|SNOMEDCT_US|Fibrosarcoma|8810/3
C0016057|T191|PT|53654007|SNOMEDCT_US|Fibrosarcoma|8810/3
C0016057|T191|IS|53654007|SNOMEDCT_US|Fibrosarcoma, NOS|8810/3
C0205766|T191|SY|0000020711|CHV|fibromyxoma|8811/0
C0205766|T191|PT|0000020711|CHV|myxofibroma|8811/0
C0205766|T191|ET|2000-6014|CSP|fibromyxoma|8811/0
C0205766|T191|ET|2000-6014|CSP|myxofibroma|8811/0
C0205766|T191|ET|D005350|MSH|Fibromyxoma|8811/0
C0205766|T191|PM|D005350|MSH|Fibromyxomas|8811/0
C0205766|T191|PEP|D005350|MSH|Myxofibroma|8811/0
C0205766|T191|PM|D005350|MSH|Myxofibromas|8811/0
C0205766|T191|SY|C66760|NCI|Fibromyxoid Neoplasm|8811/0
C0205766|T191|PT|C66760|NCI|Fibromyxoid Tumor|8811/0
C0205766|T191|SY|C66760|NCI|Fibromyxoma|8811/0
C3272426|T191|PT|C95902|NCI|Gastric Plexiform Fibromyxoma|8811/0
C0205766|T191|SY|C66760|NCI_CDISC|Fibromyxoma|8811/0
C0205766|T191|PT|C66760|NCI_CDISC|FIBROMYXOMA, BENIGN|8811/0
C0205766|T191|PT|BBG2.|RCD|Fibromyxoma|8811/0
C0205766|T191|SY|BBG2.|RCD|Myxofibroma|8811/0
C0205766|T191|SY|BBG2.|RCD|Myxoid fibroma|8811/0
C0205766|T191|PT|8664001|SNOMEDCT_US|Fibromyxoma|8811/0
C0205766|T191|SY|8664001|SNOMEDCT_US|Myxofibroma|8811/0
C0205766|T191|IS|8664001|SNOMEDCT_US|Myxofibroma, NOS|8811/0
C0205766|T191|SY|8664001|SNOMEDCT_US|Myxoid fibroma|8811/0
C1709103|T191|SY|C49025|NCI|Acral Myxoinflammatory Fibroblastic Sarcoma|8811/1
C1709103|T191|SY|C49025|NCI|Atypical Myxoinflammatory Fibroblastic Tumor|8811/1
C1709103|T191|SY|C49025|NCI|Inflammatory Myxohyaline Tumor of the Distal Extremities with Virocyte/Reed-Sternberg-Like Cells|8811/1
C1709103|T191|SY|C49025|NCI|Inflammatory Myxoid Tumor of the Soft Parts with Bizarre Giant Cells|8811/1
C1709103|T191|PT|C49025|NCI|Myxoinflammatory Fibroblastic Sarcoma|8811/1
C1709103|T191|SY|703608004|SNOMEDCT_US|Atypical myxoinflammatory fibroblastic tumor|8811/1
C1709103|T191|SYGB|703608004|SNOMEDCT_US|Atypical myxoinflammatory fibroblastic tumour|8811/1
C1709103|T191|PT|703608004|SNOMEDCT_US|Myxoinflammatory fibroblastic sarcoma|8811/1
C3714524|T191|SY|0000029984|CHV|fibromyxosarcoma|8811/3
C3714524|T191|PT|0000029984|CHV|myxofibrosarcoma|8811/3
C3714524|T191|LLT|10066948|MDR|Myxofibrosarcoma|8811/3
C3714524|T191|PT|10066948|MDR|Myxofibrosarcoma|8811/3
C3714524|T191|PT|271508|MEDCIN|fibromyxosarcoma|8811/3
C3714524|T191|PN|NOCODE|MTH|Fibromyxosarcoma|8811/3
C3714524|T191|PT|C6496|NCI|Myxofibrosarcoma|8811/3
C3714524|T191|OP|C6496|NCI|Myxoid Fibrous Histiocytoma|8811/3
C3714524|T191|OP|C6496|NCI|Myxoid Malignant Fibrous Histiocytoma|8811/3
C3714524|T191|OP|C6496|NCI|Myxoid MFH|8811/3
C3714524|T191|PT|CDR0000776765|PDQ|myxofibrosarcoma|8811/3
C3714524|T191|SY|CDR0000776765|PDQ|myxoid fibrous histiocytoma|8811/3
C3714524|T191|SY|CDR0000776765|PDQ|myxoid malignant fibrous histiocytoma|8811/3
C3714524|T191|SY|CDR0000776765|PDQ|myxoid MFH|8811/3
C3714524|T191|PT|BBG3.|RCD|Fibromyxosarcoma|8811/3
C3714524|T191|PT|6250003|SNOMEDCT_US|Fibromyxosarcoma|8811/3
C3714524|T191|IS|6250003|SNOMEDCT_US|Myxofibrosarcoma|8811/3
C3714524|T191|PT|703609007|SNOMEDCT_US|Myxofibrosarcoma|8811/3
C3714524|T191|IS|6250003|SNOMEDCT_US|Myxoid malignant fibrous histiocytoma|8811/3
C3714524|T191|SY|703609007|SNOMEDCT_US|Myxoid malignant fibrous histiocytoma|8811/3
C0334455|T191|PT|C66761|NCI|Periosteal Fibroma|8812/0
C0334455|T191|PT|BBG4.|RCD|Periosteal fibroma|8812/0
C0334455|T191|PT|53305005|SNOMEDCT_US|Periosteal fibroma|8812/0
C0334456|T191|OP|C66763|NCI|Periosteal Fibrosarcoma|8812/3
C0334456|T191|PT|C66763|NCI|Periosteal Fibrosarcoma|8812/3
C0334456|T191|PT|BBG5.|RCD|Periosteal fibrosarcoma|8812/3
C0334456|T191|SY|BBG5.|RCD|Periosteal sarcoma|8812/3
C0334456|T191|PT|65140001|SNOMEDCT_US|Periosteal fibrosarcoma|8812/3
C0334456|T191|SY|65140001|SNOMEDCT_US|Periosteal sarcoma|8812/3
C0334456|T191|IS|65140001|SNOMEDCT_US|Periosteal sarcoma, NOS|8812/3
C1275236|T191|PT|0000056964|CHV|fibroma of tendon sheath|8813/0
C0334457|T191|PT|C66764|NCI|Fascial Fibroma|8813/0
C1275236|T191|SY|C6485|NCI|Fibroma of Tendon Sheath|8813/0
C1275236|T191|SY|C6485|NCI|Fibroma of the Tendon Sheath|8813/0
C1275236|T191|PT|C6485|NCI|Tendon Sheath Fibroma|8813/0
C0334457|T191|PT|BBG6.|RCD|Fascial fibroma|8813/0
C0334457|T191|PT|52399003|SNOMEDCT_US|Fascial fibroma|8813/0
C1275236|T191|PT|703610002|SNOMEDCT_US|Fibroma of tendon sheath|8813/0
C1275236|T191|PT|403992002|SNOMEDCT_US|Fibroma of tendon sheath|8813/0
C3839308|T191|PT|703611003|SNOMEDCT_US|Palmar/plantar type fibromatosis|8813/1
C0334458|T191|PT|271509|MEDCIN|fascial fibrosarcoma|8813/3
C0334458|T191|PT|C66765|NCI|Fascial Fibrosarcoma|8813/3
C0334458|T191|PT|BBG7.|RCD|Fascial fibrosarcoma|8813/3
C0334458|T191|PT|19134004|SNOMEDCT_US|Fascial fibrosarcoma|8813/3
C0334459|T191|SY|0000029985|CHV|congenital fibrosarcoma|8814/3
C0334459|T191|PT|0000029985|CHV|infantile fibrosarcoma|8814/3
C0334459|T191|PT|MTHU018545|ICPC2ICD10ENG|congenital; fibrosarcoma|8814/3
C0334459|T191|PT|MTHU028228|ICPC2ICD10ENG|fibrosarcoma; congenital|8814/3
C0334459|T191|PT|MTHU028230|ICPC2ICD10ENG|fibrosarcoma; infantile|8814/3
C0334459|T191|PT|MTHU037878|ICPC2ICD10ENG|infantile; fibrosarcoma|8814/3
C0334459|T191|LLT|10065859|MDR|Congenital fibrosarcoma|8814/3
C0334459|T191|PT|10065859|MDR|Congenital fibrosarcoma|8814/3
C0334459|T191|PT|271510|MEDCIN|infantile fibrosarcoma|8814/3
C0334459|T191|PN|NOCODE|MTH|Infantile fibrosarcoma|8814/3
C0334459|T191|SY|C4244|NCI|Congenital Fibrosarcoma|8814/3
C0334459|T191|PT|C4244|NCI|Infantile Fibrosarcoma|8814/3
C0334459|T191|SY|10065859|NCI_CTEP-SDC|Infantile fibrosarcoma|8814/3
C0334459|T191|PT|C4244|NCI_NICHD|Infantile Fibrosarcoma|8814/3
C0334459|T191|SY|BBG8.|RCD|Congenital fibrosarcoma|8814/3
C0334459|T191|PT|BBG8.|RCD|Infantile fibrosarcoma|8814/3
C0334459|T191|SY|52040006|SNOMEDCT_US|Congenital fibrosarcoma|8814/3
C0334459|T191|PT|52040006|SNOMEDCT_US|Infantile fibrosarcoma|8814/3
C0334459|T191|PT|403996004|SNOMEDCT_US|Infantile fibrosarcoma|8814/3
C1266119|T191|PT|0000056686|CHV|solitary fibrous tumor|8815/0
C1266119|T191|SY|0000056686|CHV|solitary fibrous tumour|8815/0
C1266119|T191|LLT|10024773|MDR|Localised fibrous mesothelioma|8815/0
C1266119|T191|LLT|10062468|MDR|Localized fibrous mesothelioma|8815/0
C1266119|T191|LLT|10082807|MDR|Solitary fibrous tumor|8815/0
C1266119|T191|MTH_PT|10082804|MDR|Solitary fibrous tumor|8815/0
C1266119|T191|LLT|10082804|MDR|Solitary fibrous tumour|8815/0
C1266119|T191|PT|10082804|MDR|Solitary fibrous tumour|8815/0
C1266119|T191|PM|D054364|MSH|Fibrous Tumor, Solitary|8815/0
C1266119|T191|PM|D054364|MSH|Fibrous Tumors, Solitary|8815/0
C1266119|T191|PM|D054364|MSH|Solitary Fibrous Tumor|8815/0
C1266119|T191|MH|D054364|MSH|Solitary Fibrous Tumors|8815/0
C1266119|T191|PM|D054364|MSH|Tumor, Solitary Fibrous|8815/0
C1266119|T191|PM|D054364|MSH|Tumors, Solitary Fibrous|8815/0
C1266119|T191|PN|NOCODE|MTH|Solitary fibrous tumor|8815/0
C1266119|T191|OP|C7634|NCI|Hemangiopericytoma|8815/0
C1266119|T191|OP|C7634|NCI|Localized Fibrous Mesothelioma|8815/0
C1266119|T191|SY|C7634|NCI|Localized Fibrous Tumor|8815/0
C1266119|T191|AB|C7634|NCI|SFT|8815/0
C1266119|T191|PT|C7634|NCI|Solitary Fibrous Tumor|8815/0
C1266119|T191|OP|C7634|NCI|Submesothelial Fibroma|8815/0
C1266119|T191|SYGB|128736003|SNOMEDCT_US|Localised fibrous tumour|8815/0
C1266119|T191|SY|128736003|SNOMEDCT_US|Localized fibrous tumor|8815/0
C1266119|T191|PT|128736003|SNOMEDCT_US|Solitary fibrous tumor|8815/0
C4518377|T191|PT|734080003|SNOMEDCT_US|Solitary fibrous tumor and hemangiopericytoma grade 1|8815/0
C4518377|T191|SY|734080003|SNOMEDCT_US|Solitary fibrous tumor/hemangiopericytoma grade 1|8815/0
C1266119|T191|PTGB|128736003|SNOMEDCT_US|Solitary fibrous tumour|8815/0
C4518377|T191|PTGB|734080003|SNOMEDCT_US|Solitary fibrous tumour and haemangiopericytoma grade 1|8815/0
C4518377|T191|SYGB|734080003|SNOMEDCT_US|Solitary fibrous tumour/haemangiopericytoma grade 1|8815/0
C1266119|T191|PT|0000056686|CHV|solitary fibrous tumor|8815/1
C1266119|T191|SY|0000056686|CHV|solitary fibrous tumour|8815/1
C1266119|T191|LLT|10024773|MDR|Localised fibrous mesothelioma|8815/1
C1266119|T191|LLT|10062468|MDR|Localized fibrous mesothelioma|8815/1
C1266119|T191|LLT|10082807|MDR|Solitary fibrous tumor|8815/1
C1266119|T191|MTH_PT|10082804|MDR|Solitary fibrous tumor|8815/1
C1266119|T191|LLT|10082804|MDR|Solitary fibrous tumour|8815/1
C1266119|T191|PT|10082804|MDR|Solitary fibrous tumour|8815/1
C1266119|T191|PM|D054364|MSH|Fibrous Tumor, Solitary|8815/1
C1266119|T191|PM|D054364|MSH|Fibrous Tumors, Solitary|8815/1
C1266119|T191|PM|D054364|MSH|Solitary Fibrous Tumor|8815/1
C1266119|T191|MH|D054364|MSH|Solitary Fibrous Tumors|8815/1
C1266119|T191|PM|D054364|MSH|Tumor, Solitary Fibrous|8815/1
C1266119|T191|PM|D054364|MSH|Tumors, Solitary Fibrous|8815/1
C1266119|T191|PN|NOCODE|MTH|Solitary fibrous tumor|8815/1
C1266119|T191|OP|C7634|NCI|Hemangiopericytoma|8815/1
C1266119|T191|OP|C7634|NCI|Localized Fibrous Mesothelioma|8815/1
C1266119|T191|SY|C7634|NCI|Localized Fibrous Tumor|8815/1
C1266119|T191|AB|C7634|NCI|SFT|8815/1
C1266119|T191|PT|C7634|NCI|Solitary Fibrous Tumor|8815/1
C1266119|T191|OP|C7634|NCI|Submesothelial Fibroma|8815/1
C1266119|T191|SYGB|128736003|SNOMEDCT_US|Localised fibrous tumour|8815/1
C1266119|T191|SY|128736003|SNOMEDCT_US|Localized fibrous tumor|8815/1
C1266119|T191|PT|128736003|SNOMEDCT_US|Solitary fibrous tumor|8815/1
C1266119|T191|PTGB|128736003|SNOMEDCT_US|Solitary fibrous tumour|8815/1
C1266120|T191|PT|271511|MEDCIN|malignant solitary fibrous tumor|8815/3
C1266120|T191|PN|NOCODE|MTH|Malignant Solitary Fibrous Tumor|8815/3
C1266120|T191|OP|C6894|NCI|Malignant Hemangiopericytoma|8815/3
C1266120|T191|PT|C6894|NCI|Malignant Solitary Fibrous Tumor|8815/3
C1266120|T191|PT|C6894|NCI_CPTAC|Malignant Solitary Fibrous Tumor|8815/3
C4518379|T191|PT|734082006|SNOMEDCT_US|Solitary fibrous tumor and hemangiopericytoma grade 3|8815/3
C1266120|T191|PT|128737007|SNOMEDCT_US|Solitary fibrous tumor, malignant|8815/3
C4518379|T191|SY|734082006|SNOMEDCT_US|Solitary fibrous tumor/hemangiopericytoma grade 3|8815/3
C4518379|T191|PTGB|734082006|SNOMEDCT_US|Solitary fibrous tumour and haemangiopericytoma grade 3|8815/3
C1266120|T191|PTGB|128737007|SNOMEDCT_US|Solitary fibrous tumour, malignant|8815/3
C4518379|T191|SYGB|734082006|SNOMEDCT_US|Solitary fibrous tumour/haemangiopericytoma grade 3|8815/3
C0553647|T191|PT|0000039099|CHV|aponeurotic fibroma|8816/0
C0553647|T191|SY|0000039099|CHV|calcified fibroma|8816/0
C0553647|T191|NM|C000625499|MSH|calcifying aponeurotic fibroma|8816/0
C0553647|T191|PT|C4818|NCI|Calcifying Aponeurotic Fibroma|8816/0
C0553647|T191|SY|C4818|NCI|Juvenile Aponeurotic Fibroma|8816/0
C0553647|T191|SY|C4818|NCI|Juvenile Aponeurotic Fibrosis|8816/0
C0553647|T191|SY|X50DL|RCD|Calcifying aponeurotic fibroma|8816/0
C0553647|T191|AB|X50DL|RCD|Juv palmo-plantar fibromatosis|8816/0
C0553647|T191|PT|X50DL|RCD|Juvenile aponeurotic fibroma|8816/0
C0553647|T191|SY|X50DL|RCD|Juvenile palmo-plantar fibromatosis|8816/0
C0553647|T191|IS|133856002|SNOMEDCT_US|Aponeurotic fibroma|8816/0
C0553647|T191|OP|133856002|SNOMEDCT_US|Calcifying aponeurotic fibroma|8816/0
C0553647|T191|OP|238862009|SNOMEDCT_US|Calcifying aponeurotic fibroma|8816/0
C0553647|T191|PT|703612005|SNOMEDCT_US|Calcifying aponeurotic fibroma|8816/0
C0553647|T191|PT|703614006|SNOMEDCT_US|Calcifying aponeurotic fibroma|8816/0
C0553647|T191|PT|238862009|SNOMEDCT_US|Juvenile aponeurotic fibroma|8816/0
C0553647|T191|PT|133856002|SNOMEDCT_US|Juvenile aponeurotic fibroma|8816/0
C0553647|T191|SY|238862009|SNOMEDCT_US|Juvenile palmo-plantar fibromatosis|8816/0
C0553647|T191|SY|133856002|SNOMEDCT_US|Keasbey tumor|8816/0
C0553647|T191|SYGB|133856002|SNOMEDCT_US|Keasbey tumour|8816/0
C0553647|T191|SY|133856002|SNOMEDCT_US|Keasbey's tumor|8816/0
C0553647|T191|SYGB|133856002|SNOMEDCT_US|Keasbey's tumour|8816/0
C1332833|T191|MTH_PT|10064280|MDR|Calcifying fibrous pseudotumor|8817/0
C1332833|T191|LLT|10064284|MDR|Calcifying fibrous pseudotumor|8817/0
C1332833|T191|LLT|10064280|MDR|Calcifying fibrous pseudotumour|8817/0
C1332833|T191|PT|10064280|MDR|Calcifying fibrous pseudotumour|8817/0
C1332833|T191|PN|NOCODE|MTH|Calcifying Fibrous Pseudotumor|8817/0
C1332833|T191|SY|C6488|NCI|Calcifying Fibrous Pseudotumor|8817/0
C1332833|T191|PT|C6488|NCI|Calcifying Fibrous Tumor|8817/0
C1332833|T191|AB|C6488|NCI|CFT|8817/0
C1332833|T191|PT|703613000|SNOMEDCT_US|Calcifying fibrous tumor|8817/0
C1332833|T191|PTGB|703613000|SNOMEDCT_US|Calcifying fibrous tumour|8817/0
C0334460|T191|PT|0000029986|CHV|elastofibroma|8820/0
C0334460|T191|SY|0000029986|CHV|elastofibromas|8820/0
C0334460|T191|LLT|10079215|MDR|Elastofibroma|8820/0
C0334460|T191|PT|10079215|MDR|Elastofibroma|8820/0
C0334460|T191|PT|C4245|NCI|Elastofibroma|8820/0
C0334460|T191|SY|C4245|NCI|Elastofibroma Dorsi|8820/0
C0334460|T191|PT|BBG9.|RCD|Elastofibroma|8820/0
C0334460|T191|PT|9671003|SNOMEDCT_US|Elastofibroma|8820/0
C0079218|T191|SY|0000015129|CHV|aggressive fibromatoses|8821/1
C0079218|T191|SY|0000015129|CHV|aggressive fibromatosis|8821/1
C0079218|T191|PT|0000015129|CHV|desmoid|8821/1
C0079218|T191|PT|0000057703|CHV|desmoid fibromatosis|8821/1
C0079218|T191|SY|0000015129|CHV|desmoid tumor|8821/1
C0079218|T191|SY|0000015129|CHV|desmoid tumors|8821/1
C0079218|T191|SY|0000015129|CHV|desmoid tumour|8821/1
C0079218|T191|SY|0000015129|CHV|desmoid tumours|8821/1
C0079218|T191|SY|0000015129|CHV|desmoids|8821/1
C0079218|T191|SY|0000057703|CHV|fibromatosis desmoid|8821/1
C0079218|T191|SY|0000015129|CHV|musculoaponeurotic fibromatosis|8821/1
C0079218|T191|PT|HP:0100245|HPO|Desmoid tumors|8821/1
C0079218|T191|PT|MTHU022670|ICPC2ICD10ENG|desmoid|8821/1
C0079218|T191|LLT|10059353|MDR|Desmoid tumor|8821/1
C0079218|T191|MTH_PT|10059352|MDR|Desmoid tumor|8821/1
C0079218|T191|LLT|10059352|MDR|Desmoid tumour|8821/1
C0079218|T191|PT|10059352|MDR|Desmoid tumour|8821/1
C0079218|T191|PT|356604|MEDCIN|Deep fibromatosis|8821/1
C0079218|T191|PT|31704|MEDCIN|desmoid tumor|8821/1
C0079218|T191|SY|356604|MEDCIN|soft tissue neoplasm benign - deep fibromatosis|8821/1
C0079218|T191|PM|D018222|MSH|Aggressive Fibromatoses|8821/1
C0079218|T191|PM|D018222|MSH|Aggressive Fibromatosis|8821/1
C0079218|T191|ET|D018222|MSH|Desmoid|8821/1
C0079218|T191|PM|D018222|MSH|Desmoids|8821/1
C0079218|T191|PM|D018222|MSH|Fibromatoses, Aggressive|8821/1
C0079218|T191|MH|D018222|MSH|Fibromatosis, Aggressive|8821/1
C0079218|T191|SY|C9182|NCI|Aggressive Fibromatosis|8821/1
C0079218|T191|SY|C9182|NCI|Deep Fibromatosis|8821/1
C0079218|T191|SY|C9182|NCI|Deep Fibromatosis/Desmoid Tumor|8821/1
C0079218|T191|SY|C9182|NCI|Desmoid Fibromatosis|8821/1
C0079218|T191|SY|C9182|NCI|Desmoid Tumor|8821/1
C0079218|T191|PT|C9182|NCI|Desmoid-Type Fibromatosis|8821/1
C0079218|T191|DN|C9182|NCI_CTRP|Deep Fibromatosis/Desmoid Tumor|8821/1
C0079218|T191|PT|CDR0000045390|NCI_NCI-GLOSS|desmoid tumor|8821/1
C0079218|T191|SY|CDR0000041704|PDQ|aggressive fibromatosis|8821/1
C0079218|T191|PSC|CDR0000041704|PDQ|desmoid tumor|8821/1
C0079218|T191|SY|CDR0000041704|PDQ|musculoaponeurotic fibromatosis|8821/1
C0079218|T191|PT|BBGA.|RCD|Aggressive fibromatosis|8821/1
C0079218|T191|SY|BBGA.|RCD|Desmoid|8821/1
C0079218|T191|SY|BBGA.|RCD|Extra-abdominal desmoid|8821/1
C0079218|T191|SY|BBGA.|RCD|Invasive fibroma|8821/1
C0079218|T191|PT|725049005|SNOMEDCT_US|Aggressive fibromatosis|8821/1
C0079218|T191|PT|47284001|SNOMEDCT_US|Aggressive fibromatosis|8821/1
C0079218|T191|OAP|400055004|SNOMEDCT_US|Deep fibromatosis|8821/1
C0079218|T191|SY|725049005|SNOMEDCT_US|Deep fibromatosis|8821/1
C0079218|T191|SY|47284001|SNOMEDCT_US|Desmoid|8821/1
C0079218|T191|OAP|399994005|SNOMEDCT_US|Desmoid fibromatosis|8821/1
C0079218|T191|SY|725049005|SNOMEDCT_US|Desmoid fibromatosis|8821/1
C0079218|T191|SY|725049005|SNOMEDCT_US|Desmoid tumor|8821/1
C0079218|T191|SY|47284001|SNOMEDCT_US|Desmoid tumor|8821/1
C0079218|T191|SYGB|725049005|SNOMEDCT_US|Desmoid tumour|8821/1
C0079218|T191|SYGB|47284001|SNOMEDCT_US|Desmoid tumour|8821/1
C0079218|T191|SY|725049005|SNOMEDCT_US|Desmoid type fibromatosis|8821/1
C0079218|T191|SY|47284001|SNOMEDCT_US|Desmoid-type fibromatosis|8821/1
C0079218|T191|IS|47284001|SNOMEDCT_US|Desmoid, NOS|8821/1
C0079218|T191|IS|47284001|SNOMEDCT_US|Extra-abdominal desmoid|8821/1
C0079218|T191|SY|47284001|SNOMEDCT_US|Invasive fibroma|8821/1
C0206646|T191|SY|0000020992|CHV|abdominal desmoid|8822/1
C0206646|T191|SY|0000020992|CHV|abdominal fibromatosis|8822/1
C0206646|T191|SY|0000020992|CHV|fibromatosis abdominal|8822/1
C0206646|T191|PT|0000020992|CHV|mesenteric fibromatosis|8822/1
C0206646|T191|SY|0000020992|CHV|retroperitoneal fibromatosis|8822/1
C0206646|T191|PT|MTHU002229|ICPC2ICD10ENG|abdominal; desmoid|8822/1
C0206646|T191|PT|MTHU002230|ICPC2ICD10ENG|abdominal; desmoid tumor|8822/1
C0206646|T191|PT|MTHU002243|ICPC2ICD10ENG|abdominal; tumor, desmoid|8822/1
C0206646|T191|PT|MTHU022671|ICPC2ICD10ENG|desmoid; abdominal|8822/1
C0206646|T191|PT|MTHU022672|ICPC2ICD10ENG|desmoid; tumor, abdominal|8822/1
C0206646|T191|PT|MTHU028198|ICPC2ICD10ENG|fibromatosis; retroperitoneal|8822/1
C0206646|T191|PT|MTHU064571|ICPC2ICD10ENG|retroperitoneal; fibromatosis|8822/1
C0206646|T191|PT|MTHU077007|ICPC2ICD10ENG|tumor; abdominal, desmoid|8822/1
C0206646|T191|PT|MTHU077044|ICPC2ICD10ENG|tumor; desmoid, abdominal|8822/1
C0206646|T191|LLT|10059354|MDR|Abdominal fibromatosis|8822/1
C0206646|T191|PT|339773|MEDCIN|Abdominal fibromatosis|8822/1
C0206646|T191|PM|D018221|MSH|Abdominal Fibromatoses|8822/1
C0206646|T191|PM|D018221|MSH|Abdominal Fibromatosis|8822/1
C0206646|T191|PM|D018221|MSH|Fibromatoses, Abdominal|8822/1
C0206646|T191|MH|D018221|MSH|Fibromatosis, Abdominal|8822/1
C0206646|T191|SY|C3741|NCI|Abdominal Desmoid|8822/1
C0206646|T191|SY|C3741|NCI|Abdominal Desmoid Tumor|8822/1
C0206646|T191|SY|C3741|NCI|Abdominal Fibromatosis|8822/1
C0206646|T191|SY|C3741|NCI|Intraabdominal Desmoid|8822/1
C0206646|T191|SY|C3741|NCI|Intraabdominal Desmoid Tumor|8822/1
C0206646|T191|SY|C3741|NCI|Intraabdominal Fibromatosis|8822/1
C0206646|T191|SY|C3741|NCI|Mesenteric Desmoid|8822/1
C0206646|T191|SY|C3741|NCI|Mesenteric Desmoid Tumor|8822/1
C0206646|T191|SY|C3741|NCI|Mesenteric Fibromatosis|8822/1
C0206646|T191|SY|BBGB.|RCD|Abdominal desmoid|8822/1
C0206646|T191|PT|BBGB.|RCD|Abdominal fibromatosis|8822/1
C0206646|T191|SY|BBGB.|RCD|Mesenteric fibromatosis|8822/1
C0206646|T191|SY|BBGB.|RCD|Retroperitoneal fibromatosis|8822/1
C0206646|T191|OAS|45187003|SNOMEDCT_US|Abdominal desmoid|8822/1
C0206646|T191|SY|400153009|SNOMEDCT_US|Abdominal desmoid tumor|8822/1
C0206646|T191|SYGB|400153009|SNOMEDCT_US|Abdominal desmoid tumour|8822/1
C0206646|T191|PT|400153009|SNOMEDCT_US|Abdominal fibromatosis|8822/1
C0206646|T191|OAP|45187003|SNOMEDCT_US|Abdominal fibromatosis|8822/1
C0206646|T191|OAS|45187003|SNOMEDCT_US|Mesenteric fibromatosis|8822/1
C0206646|T191|OAS|45187003|SNOMEDCT_US|Retroperitoneal fibromatosis|8822/1
C0206645|T191|PT|39816|MEDCIN|desmoplastic fibroma of bone|8823/0
C0206645|T191|ET|D018220|MSH|Collagenous Fibroma|8823/0
C0206645|T191|PM|D018220|MSH|Collagenous Fibromas|8823/0
C0206645|T191|ET|D018220|MSH|Desmoplastic Fibroblastoma|8823/0
C0206645|T191|PM|D018220|MSH|Desmoplastic Fibroblastomas|8823/0
C0206645|T191|PM|D018220|MSH|Desmoplastic Fibroma|8823/0
C0206645|T191|PM|D018220|MSH|Desmoplastic Fibromas|8823/0
C0206645|T191|PM|D018220|MSH|Fibroblastoma, Desmoplastic|8823/0
C0206645|T191|PM|D018220|MSH|Fibroma, Collagenous|8823/0
C0206645|T191|MH|D018220|MSH|Fibroma, Desmoplastic|8823/0
C0206645|T191|PN|NOCODE|MTH|Desmoplastic fibroma|8823/0
C0206645|T191|PT|C3740|NCI|Bone Desmoplastic Fibroma|8823/0
C0206645|T191|SY|C3740|NCI|Desmoid Tumor of Bone|8823/0
C0206645|T191|SY|C3740|NCI|Desmoplastic Fibroma|8823/0
C0206645|T191|SY|C3740|NCI|Desmoplastic Fibroma of Bone|8823/0
C0206645|T191|SY|C3740|NCI|Desmoplastic Fibroma of the Bone|8823/0
C0206645|T191|SY|C3740|NCI|Osseous Desmoplastic Fibroma|8823/0
C0206645|T191|SY|C3740|NCI_CDISC|Desmoid Tumor of Bone|8823/0
C0206645|T191|SY|C3740|NCI_CDISC|Desmoplastic Fibroma|8823/0
C0206645|T191|SY|C3740|NCI_CDISC|Desmoplastic Fibroma of Bone|8823/0
C0206645|T191|SY|C3740|NCI_CDISC|Desmoplastic Fibroma of the Bone|8823/0
C0206645|T191|SY|C3740|NCI_CDISC|Osseous Desmoplastic Fibroma|8823/0
C0206645|T191|PT|C3740|NCI_CDISC|OSTEOFIBROMA, BENIGN|8823/0
C0206645|T191|PT|BBGC.|RCD|Desmoplastic fibroma|8823/0
C0206645|T191|OAP|128861007|SNOMEDCT_US|Desmoplastic fibroma|8823/0
C0206645|T191|PT|6842002|SNOMEDCT_US|Desmoplastic fibroma|8823/0
C0206645|T191|IS|6842002|SNOMEDCT_US|Desmoplastic fibroma -RETIRED-|8823/0
C0206645|T191|OF|6842002|SNOMEDCT_US|Desmoplastic fibroma -RETIRED-|8823/0
C0206645|T191|PT|39816|MEDCIN|desmoplastic fibroma of bone|8823/1
C0206645|T191|ET|D018220|MSH|Collagenous Fibroma|8823/1
C0206645|T191|PM|D018220|MSH|Collagenous Fibromas|8823/1
C0206645|T191|ET|D018220|MSH|Desmoplastic Fibroblastoma|8823/1
C0206645|T191|PM|D018220|MSH|Desmoplastic Fibroblastomas|8823/1
C0206645|T191|PM|D018220|MSH|Desmoplastic Fibroma|8823/1
C0206645|T191|PM|D018220|MSH|Desmoplastic Fibromas|8823/1
C0206645|T191|PM|D018220|MSH|Fibroblastoma, Desmoplastic|8823/1
C0206645|T191|PM|D018220|MSH|Fibroma, Collagenous|8823/1
C0206645|T191|MH|D018220|MSH|Fibroma, Desmoplastic|8823/1
C0206645|T191|PN|NOCODE|MTH|Desmoplastic fibroma|8823/1
C0206645|T191|PT|C3740|NCI|Bone Desmoplastic Fibroma|8823/1
C0206645|T191|SY|C3740|NCI|Desmoid Tumor of Bone|8823/1
C0206645|T191|SY|C3740|NCI|Desmoplastic Fibroma|8823/1
C0206645|T191|SY|C3740|NCI|Desmoplastic Fibroma of Bone|8823/1
C0206645|T191|SY|C3740|NCI|Desmoplastic Fibroma of the Bone|8823/1
C0206645|T191|SY|C3740|NCI|Osseous Desmoplastic Fibroma|8823/1
C0206645|T191|SY|C3740|NCI_CDISC|Desmoid Tumor of Bone|8823/1
C0206645|T191|SY|C3740|NCI_CDISC|Desmoplastic Fibroma|8823/1
C0206645|T191|SY|C3740|NCI_CDISC|Desmoplastic Fibroma of Bone|8823/1
C0206645|T191|SY|C3740|NCI_CDISC|Desmoplastic Fibroma of the Bone|8823/1
C0206645|T191|SY|C3740|NCI_CDISC|Osseous Desmoplastic Fibroma|8823/1
C0206645|T191|PT|C3740|NCI_CDISC|OSTEOFIBROMA, BENIGN|8823/1
C0206645|T191|PT|BBGC.|RCD|Desmoplastic fibroma|8823/1
C0206645|T191|PT|6842002|SNOMEDCT_US|Desmoplastic fibroma|8823/1
C0206645|T191|OAP|128861007|SNOMEDCT_US|Desmoplastic fibroma|8823/1
C0206645|T191|IS|6842002|SNOMEDCT_US|Desmoplastic fibroma -RETIRED-|8823/1
C0206645|T191|OF|6842002|SNOMEDCT_US|Desmoplastic fibroma -RETIRED-|8823/1
C1266121|T191|PT|0000056687|CHV|myofibroma|8824/0
C1266121|T191|LLT|10075377|MDR|Myofibroma|8824/0
C1266121|T191|MH|D047708|MSH|Myofibroma|8824/0
C1266121|T191|PM|D047708|MSH|Myofibromas|8824/0
C1368237|T191|PN|NOCODE|MTH|Solitary Myofibromatosis|8824/0
C1368237|T191|OP|C7052|NCI|Infantile Hemangiopericytoma|8824/0
C1368237|T191|PT|C7052|NCI|Myofibroma|8824/0
C1266121|T191|SY|Xa99u|RCD|Myofibroma|8824/0
C1266121|T191|SY|44598004|SNOMEDCT_US|Lipoleiomyoma|8824/0
C1266121|T191|PT|128917003|SNOMEDCT_US|Myofibroma|8824/0
C1266121|T191|IS|44598004|SNOMEDCT_US|Myofibroma|8824/0
C0206648|T191|SY|0000020994|CHV|juvenile fibromatosis|8824/1
C0206648|T191|PT|0000020994|CHV|myofibromatosis|8824/1
C0206648|T191|PT|HP:0020135|HPO|Myofibromatosis|8824/1
C0206648|T191|PT|MTHU051117|ICPC2ICD10ENG|myofibromatosis|8824/1
C0206648|T191|PM|D018224|MSH|Myofibromatoses|8824/1
C0206648|T191|MH|D018224|MSH|Myofibromatosis|8824/1
C0206648|T191|PN|NOCODE|MTH|Myofibromatosis|8824/1
C0206648|T191|OP|C3742|NCI|Infantile Hemangiopericytoma|8824/1
C0206648|T191|SY|C3742|NCI|Infantile Myofibromatosis|8824/1
C0206648|T191|SY|C3742|NCI|Multicentric Myofibromatosis|8824/1
C0206648|T191|PT|C3742|NCI|Myofibromatosis|8824/1
C0206648|T191|PT|X77oZ|RCD|Myofibromatosis|8824/1
C0206648|T191|OP|BBGN.|RCDSY|Myofibromatosis|8824/1
C0206648|T191|OAP|253043004|SNOMEDCT_US|Myofibromatosis|8824/1
C0206648|T191|OAP|238860001|SNOMEDCT_US|Myofibromatosis|8824/1
C0206648|T191|OF|238860001|SNOMEDCT_US|Myofibromatosis|8824/1
C0206648|T191|PT|73767002|SNOMEDCT_US|Myofibromatosis|8824/1
C0242404|T191|PEP|D009379|MSH|Myofibroblastoma|8825/0
C0242404|T191|PM|D009379|MSH|Myofibroblastomas|8825/0
C0242404|T191|PT|C49012|NCI|Myofibroblastoma|8825/0
C0242404|T191|PT|128738002|SNOMEDCT_US|Myofibroblastoma|8825/0
C3164851|T191|PT|449078000|SNOMEDCT_US|Palisaded myofibroblastoma|8825/0
C0334121|T191|PT|0000029918|CHV|inflammatory pseudotumor|8825/1
C0334121|T191|SY|0000029918|CHV|inflammatory pseudotumors|8825/1
C0334121|T191|SY|0000029918|CHV|inflammatory pseudotumour|8825/1
C0334121|T191|PT|0000056688|CHV|myofibroblastic tumor|8825/1
C0334121|T191|SY|0000056688|CHV|myofibroblastic tumors|8825/1
C0334121|T191|SY|0000056688|CHV|myofibroblastic tumour|8825/1
C0334121|T191|SY|0000029918|CHV|pseudotumor inflammatory|8825/1
C0334121|T191|LLT|10067918|MDR|Inflammatory myofibroblastic tumor|8825/1
C0334121|T191|MTH_PT|10067917|MDR|Inflammatory myofibroblastic tumor|8825/1
C0334121|T191|LLT|10067917|MDR|Inflammatory myofibroblastic tumour|8825/1
C0334121|T191|PT|10067917|MDR|Inflammatory myofibroblastic tumour|8825/1
C0334121|T191|LLT|10068332|MDR|Inflammatory pseudotumor|8825/1
C0334121|T191|MTH_PT|10068331|MDR|Inflammatory pseudotumor|8825/1
C0334121|T191|LLT|10068331|MDR|Inflammatory pseudotumour|8825/1
C0334121|T191|PT|10068331|MDR|Inflammatory pseudotumour|8825/1
C0334121|T191|LLT|10067746|MDR|Myofibroblastic tumor|8825/1
C0334121|T191|LLT|10067839|MDR|Myofibroblastic tumour|8825/1
C0334121|T191|DEV|D006104|MSH|INFLAMM PSEUDOTUMOR|8825/1
C0334121|T191|PEP|D006104|MSH|Inflammatory Pseudotumor|8825/1
C0334121|T191|PM|D006104|MSH|Inflammatory Pseudotumors|8825/1
C0334121|T191|DEV|D006104|MSH|PSEUDOTUMOR INFLAMM|8825/1
C0334121|T191|ET|D006104|MSH|Pseudotumor, Inflammatory|8825/1
C0334121|T191|PM|D006104|MSH|Pseudotumors, Inflammatory|8825/1
C0334121|T191|PN|NOCODE|MTH|Inflammatory Myofibroblastic Tumor|8825/1
C0334121|T191|AB|C6481|NCI|IMT|8825/1
C0334121|T191|SY|C6481|NCI|Inflammatory Fibrosarcoma|8825/1
C0334121|T191|SY|C6481|NCI|Inflammatory Myofibroblastic Neoplasm|8825/1
C0334121|T191|PT|C6481|NCI|Inflammatory Myofibroblastic Tumor|8825/1
C0334121|T191|SY|C6481|NCI|Inflammatory Pseudotumor|8825/1
C0334121|T191|PT|771233008|SNOMEDCT_US|Inflammatory myofibroblastic tumor|8825/1
C0334121|T191|SY|116064009|SNOMEDCT_US|Inflammatory myofibroblastic tumor|8825/1
C0334121|T191|PTGB|771233008|SNOMEDCT_US|Inflammatory myofibroblastic tumour|8825/1
C0334121|T191|SYGB|116064009|SNOMEDCT_US|Inflammatory myofibroblastic tumour|8825/1
C0334121|T191|PT|35073002|SNOMEDCT_US|Inflammatory pseudotumor|8825/1
C0334121|T191|PTGB|35073002|SNOMEDCT_US|Inflammatory pseudotumour|8825/1
C0334121|T191|PT|116064009|SNOMEDCT_US|Myofibroblastic tumor|8825/1
C0334121|T191|PTGB|116064009|SNOMEDCT_US|Myofibroblastic tumour|8825/1
C1708751|T191|PN|NOCODE|MTH|Low grade myofibroblastic sarcoma|8825/3
C1708751|T191|PT|C49024|NCI|Low Grade Myofibroblastic Sarcoma|8825/3
C1708751|T191|SY|C49024|NCI|Myofibrosarcoma|8825/3
C1708751|T191|PT|703615007|SNOMEDCT_US|Low grade myofibroblastic sarcoma|8825/3
C1266123|T191|LLT|10074730|MDR|Angiomyofibroblastoma|8826/0
C1266123|T191|PT|10074730|MDR|Angiomyofibroblastoma|8826/0
C1266123|T191|PT|C49016|NCI|Angiomyofibroblastoma|8826/0
C1266123|T191|PT|128739005|SNOMEDCT_US|Angiomyofibroblastoma|8826/0
C1266124|T191|PN|NOCODE|MTH|tumor miofibroblástico peribronquial congénito|8827/1
C1266124|T191|SY|C142823|NCI|Congenital Bronchopulmonary Leiomyosarcoma|8827/1
C1266124|T191|SY|C142823|NCI|Congenital Fibrosarcoma|8827/1
C1266124|T191|SY|C142823|NCI|Congenital Mesenchymal Malformation of Lung|8827/1
C1266124|T191|PT|C142823|NCI|Congenital Peribronchial Myofibroblastic Tumor|8827/1
C1266124|T191|SY|C142823|NCI|Congenital Pulmonary Myofibroblastic Tumor|8827/1
C1518038|T191|PT|C39740|NCI|Lung Inflammatory Myofibroblastic Tumor|8827/1
C1266124|T191|SY|C142823|NCI|Neonatal Pulmonary Hamartoma|8827/1
C1266124|T191|SY|128740007|SNOMEDCT_US|Congenital peribronchial myofibroblastic tumor|8827/1
C1266124|T191|SYGB|128740007|SNOMEDCT_US|Congenital peribronchial myofibroblastic tumour|8827/1
C1266124|T191|PT|128740007|SNOMEDCT_US|Myofibroblastic tumor, peribronchial|8827/1
C1266124|T191|PTGB|128740007|SNOMEDCT_US|Myofibroblastic tumour, peribronchial|8827/1
C0410005|T047|SY|0000021377|CHV|fasciitis nodular|8828/0
C0410005|T047|PT|0000021377|CHV|nodular fasciitis|8828/0
C0410005|T047|SY|0000021377|CHV|pseudosarcomatous fibromatosis|8828/0
C0410005|T047|DI|U000635|DXP|FASCIITIS, NODULAR|8828/0
C0410005|T047|PT|M72.3|ICD10|Nodular fasciitis|8828/0
C0410005|T047|PT|M72.4|ICD10|Pseudosarcomatous fibromatosis|8828/0
C0410005|T047|ET|M72.4|ICD10CM|Nodular fasciitis|8828/0
C0410005|T047|PT|M72.4|ICD10CM|Pseudosarcomatous fibromatosis|8828/0
C0410005|T047|AB|M72.4|ICD10CM|Pseudosarcomatous fibromatosis|8828/0
C0410005|T047|PT|MTHU027939|ICPC2ICD10ENG|fasciitis; nodular|8828/0
C0410005|T047|PT|MTHU028197|ICPC2ICD10ENG|fibromatosis; pseudosarcomatous|8828/0
C0410005|T047|PT|MTHU053407|ICPC2ICD10ENG|nodular; fasciitis|8828/0
C0410005|T047|PT|MTHU062327|ICPC2ICD10ENG|pseudosarcomatous; fibromatosis|8828/0
C0410005|T047|PT|10065988|MDR|Nodular fasciitis|8828/0
C0410005|T047|LLT|10065988|MDR|Nodular fasciitis|8828/0
C0410005|T047|PT|96818|MEDCIN|nodular fasciitis|8828/0
C0410005|T047|ET|728.79|MTHICD9|Nodular fasciitis|8828/0
C0410005|T047|ET|728.79|MTHICD9|Pseudosarcomatous Fibromatosis|8828/0
C0410005|T047|PT|C3827|NCI|Nodular Fasciitis|8828/0
C0410005|T047|SY|C3827|NCI|Pseudosarcomatous Fasciitis|8828/0
C0410005|T047|PT|N2372|RCD|Nodular fasciitis|8828/0
C0410005|T047|OP|N2373|RCD|Pseudosarcomatous fibromatosis|8828/0
C0410005|T047|OAS|268106003|SNOMEDCT_US|Fasciitis - nodular|8828/0
C0410005|T047|OAS|156729009|SNOMEDCT_US|Fasciitis - nodular|8828/0
C0410005|T047|OAS|35548007|SNOMEDCT_US|Infiltrative fasciitis|8828/0
C0410005|T047|SY|400138001|SNOMEDCT_US|Infiltrative fasciitis|8828/0
C0410005|T047|PT|703616008|SNOMEDCT_US|Nodular fasciitis|8828/0
C0410005|T047|PT|400138001|SNOMEDCT_US|Nodular fasciitis|8828/0
C0410005|T047|OAP|35548007|SNOMEDCT_US|Nodular fasciitis|8828/0
C0410005|T047|OAS|268106003|SNOMEDCT_US|Nodular fasciitis|8828/0
C0410005|T047|OAS|156729009|SNOMEDCT_US|Nodular fasciitis|8828/0
C0410005|T047|OAS|35548007|SNOMEDCT_US|Pseudosarcomatous fasciitis|8828/0
C0410005|T047|SY|400138001|SNOMEDCT_US|Pseudosarcomatous fasciitis|8828/0
C0410005|T047|IS|47284001|SNOMEDCT_US|Pseudosarcomatous fibromatosis|8828/0
C0410005|T047|OAP|203057005|SNOMEDCT_US|Pseudosarcomatous fibromatosis|8828/0
C0410005|T047|OAS|35548007|SNOMEDCT_US|Pseudosarcomatous fibromatosis|8828/0
C0410005|T047|SY|400138001|SNOMEDCT_US|Pseudosarcomatous fibromatosis|8828/0
C0206644|T191|PT|0056519|CCPSS|FIBROUS HISTIOCYTOMA|8830/0
C0206644|T191|SY|0000020991|CHV|benign fibrous histiocytoma|8830/0
C0206644|T191|PT|0000020991|CHV|fibrous histiocytoma|8830/0
C0206644|T191|SY|0000020991|CHV|fibrous histiocytomas|8830/0
C0206644|T191|SY|0000020991|CHV|fibroxanthoma|8830/0
C0206644|T191|SY|0000020991|CHV|xanthofibroma|8830/0
C0206644|T191|SY|NOCODE|DXP|FIBROXANTHOMA|8830/0
C0206644|T191|LLT|10053717|MDR|Fibrous histiocytoma|8830/0
C0206644|T191|PT|10053717|MDR|Fibrous histiocytoma|8830/0
C0206644|T191|LLT|10069780|MDR|Fibroxanthoma|8830/0
C0206644|T191|ET|D018219|MSH|Benign Fibrous Histiocytoma|8830/0
C0206644|T191|PM|D018219|MSH|Benign Fibrous Histiocytomas|8830/0
C0206644|T191|PM|D018219|MSH|Fibrous Histiocytoma|8830/0
C0206644|T191|PM|D018219|MSH|Fibrous Histiocytoma, Benign|8830/0
C0206644|T191|PM|D018219|MSH|Fibrous Histiocytomas|8830/0
C0206644|T191|PM|D018219|MSH|Fibrous Histiocytomas, Benign|8830/0
C0206644|T191|MH|D018219|MSH|Histiocytoma, Benign Fibrous|8830/0
C0206644|T191|ET|D018219|MSH|Histiocytoma, Fibrous|8830/0
C0206644|T191|PM|D018219|MSH|Histiocytomas, Benign Fibrous|8830/0
C0206644|T191|PM|D018219|MSH|Histiocytomas, Fibrous|8830/0
C0206644|T191|PN|NOCODE|MTH|Histiocytoma, Benign Fibrous|8830/0
C0206644|T191|PT|C3739|NCI|Benign Fibrous Histiocytoma|8830/0
C1707544|T191|SY|C49079|NCI|Cutaneous Epithelioid Fibrous Histiocytoma|8830/0
C1707544|T191|PT|C49079|NCI|Cutaneous Fibrous Histiocytoma, Epithelioid Variant|8830/0
C1707544|T191|SY|C49079|NCI|Epithelioid Fibrous Histiocytoma|8830/0
C0206644|T191|SY|C3739|NCI|Fibrous Histiocytoma|8830/0
C0206644|T191|SY|C3739|NCI_CDISC|Fibrous Histiocytoma|8830/0
C0206644|T191|PT|C3739|NCI_CDISC|HISTIOCYTOMA, FIBROUS, BENIGN|8830/0
C0206644|T191|PT|Xa99m|RCD|Fibrous histiocytoma|8830/0
C0206644|T191|SY|Xa99m|RCD|Fibroxanthoma|8830/0
C0206644|T191|SY|Xa99m|RCD|Xanthofibroma|8830/0
C0206644|T191|OP|BBGD.|RCDSY|Fibrous histiocytoma NOS|8830/0
C0206644|T191|OP|BBGG.|RCDSY|Fibroxanthoma NOS|8830/0
C0206644|T191|IS|BBGG.|RCDSY|Xanthofibroma|8830/0
C0206644|T191|PT|25889007|SNOMEDCT_US|Benign fibrous histiocytoma|8830/0
C1707544|T191|PT|816970007|SNOMEDCT_US|Epithelioid fibrous histiocytoma|8830/0
C0206644|T191|SY|25889007|SNOMEDCT_US|Fibrous histiocytoma|8830/0
C0206644|T191|IS|25889007|SNOMEDCT_US|Fibrous histiocytoma, NOS|8830/0
C0206644|T191|SY|25889007|SNOMEDCT_US|Fibroxanthoma|8830/0
C0206644|T191|IS|25889007|SNOMEDCT_US|Fibroxanthoma, NOS|8830/0
C0206644|T191|SY|25889007|SNOMEDCT_US|Xanthofibroma|8830/0
C0346053|T191|SY|0000029987|CHV|atypical fibrous histiocytoma|8830/1
C0346053|T191|PT|0000029987|CHV|atypical fibroxanthoma|8830/1
C0346053|T191|SY|0000029987|CHV|fibroxanthoma atypical|8830/1
C0346053|T191|LLT|10064755|MDR|Atypical fibroxanthoma|8830/1
C0346053|T191|PT|10064755|MDR|Atypical fibroxanthoma|8830/1
C0346053|T191|PT|355139|MEDCIN|skin neoplasm malignant fibrohistiocytic atypical fibroxanthoma|8830/1
C0346053|T191|PN|NOCODE|MTH|Atypical fibroxanthoma of skin|8830/1
C0346053|T191|SY|C4246|NCI|Atypical Cutaneous Fibroxanthoma|8830/1
C0346053|T191|SY|C4246|NCI|Atypical Fibrous Histiocytoma|8830/1
C0346053|T191|PT|C4246|NCI|Atypical Fibroxanthoma|8830/1
C0346053|T191|SY|C4246|NCI|Atypical Fibroxanthoma of Skin|8830/1
C0346053|T191|SY|C4246|NCI|Atypical Fibroxanthoma of the Skin|8830/1
C0346053|T191|SY|C4246|NCI|Atypical Skin Fibroxanthoma|8830/1
C0346053|T191|OP|C4246|NCI|Superficial Malignant Fibrous Histiocytoma|8830/1
C0346053|T191|PT|BBGE.|RCD|Atypical fibrous histiocytoma|8830/1
C0346053|T191|SY|BBGE.|RCD|Atypical fibroxanthoma|8830/1
C0346053|T191|PT|X78Tm|RCD|Atypical fibroxanthoma of skin|8830/1
C0346053|T191|SY|X78Tm|RCD|Fibroxanthosarcoma of skin|8830/1
C0346053|T191|PT|26496005|SNOMEDCT_US|Atypical fibrous histiocytoma|8830/1
C0346053|T191|OAP|189771003|SNOMEDCT_US|Atypical fibrous histiocytoma|8830/1
C0346053|T191|OF|189771003|SNOMEDCT_US|Atypical fibrous histiocytoma|8830/1
C0346053|T191|SY|26496005|SNOMEDCT_US|Atypical fibroxanthoma|8830/1
C0346053|T191|PT|254754005|SNOMEDCT_US|Atypical fibroxanthoma of skin|8830/1
C0346053|T191|OAP|254755006|SNOMEDCT_US|Atypical fibroxanthoma of skin|8830/1
C0346053|T191|OF|254755006|SNOMEDCT_US|Atypical fibroxanthoma of skin|8830/1
C0346053|T191|SY|254754005|SNOMEDCT_US|Fibroxanthosarcoma of skin|8830/1
C0334463|T191|PT|0025244|CCPSS|HISTIOCYTOMA MALIGNANT FIBROUS|8830/3
C0334463|T191|SY|0000029988|CHV|fibrous histiocytoma malignant|8830/3
C0334463|T191|PT|0000029988|CHV|malignant fibrous histiocytoma|8830/3
C0334463|T191|LLT|10016665|MDR|Fibrous histiocytoma malignant|8830/3
C0334463|T191|HT|10025553|MDR|Fibrous histiocytomas malignant|8830/3
C0334463|T191|LLT|10025552|MDR|Malignant fibrous histiocytoma|8830/3
C0334463|T191|PT|10025552|MDR|Malignant fibrous histiocytoma|8830/3
C0334463|T191|LLT|10025556|MDR|Malignant fibrous histiocytoma NOS|8830/3
C0334463|T191|LLT|10025562|MDR|Malignant fibrous histiocytoma stage unspecified|8830/3
C0334463|T191|PT|271533|MEDCIN|malignant fibrous histiocytoma|8830/3
C0334463|T191|PM|D051677|MSH|Fibrohistiocytic Tumor, Malignant|8830/3
C0334463|T191|PM|D051677|MSH|Fibrohistiocytic Tumors, Malignant|8830/3
C0334463|T191|PM|D051677|MSH|Fibrous Histiocytoma, Malignant|8830/3
C0334463|T191|PM|D051677|MSH|Fibrous Histiocytomas, Malignant|8830/3
C0334463|T191|MH|D051677|MSH|Histiocytoma, Malignant Fibrous|8830/3
C0334463|T191|PM|D051677|MSH|Histiocytomas, Malignant Fibrous|8830/3
C0334463|T191|PM|D051677|MSH|Malignant Fibrohistiocytic Tumor|8830/3
C0334463|T191|ET|D051677|MSH|Malignant Fibrohistiocytic Tumors|8830/3
C0334463|T191|ET|D051677|MSH|Malignant Fibrous Histiocytoma|8830/3
C0334463|T191|PM|D051677|MSH|Malignant Fibrous Histiocytomas|8830/3
C0334463|T191|PM|D051677|MSH|Tumor, Malignant Fibrohistiocytic|8830/3
C0334463|T191|PM|D051677|MSH|Tumors, Malignant Fibrohistiocytic|8830/3
C0334463|T191|PN|NOCODE|MTH|Malignant Fibrous Histiocytoma|8830/3
C0334463|T191|OP|C4247|NCI|Fibroxanthosarcoma|8830/3
C0334463|T191|OP|C4247|NCI|Malignant Fibrous Histiocytoma|8830/3
C0334463|T191|OP|C4247|NCI|Malignant Fibroxanthoma|8830/3
C0334463|T191|AB|C4247|NCI|MFH|8830/3
C0334463|T191|OP|C4247|NCI|Storiform-Pleomorphic Fibrous Histiocytoma|8830/3
C0334463|T191|SY|C4247|NCI|Storiform-Pleomorphic Malignant Fibrous Histiocytoma|8830/3
C0334463|T191|OP|C4247|NCI|Storiform-Pleomorphic MFH|8830/3
C0334463|T191|SY|C4247|NCI|Unclassified Pleomorphic Sarcoma|8830/3
C0334463|T191|PT|C4247|NCI|Undifferentiated Pleomorphic Sarcoma|8830/3
C0334463|T191|SY|C4247|NCI|Undifferentiated Pleomorphic Soft Tissue Sarcoma|8830/3
C0334463|T191|AB|C4247|NCI|UPS|8830/3
C0334463|T191|PT|C4247|NCI_CDISC|FIBROSARCOMA, PLEOMORPHIC, MALIGNANT|8830/3
C0334463|T191|SY|C4247|NCI_CDISC|Fibroxanthosarcoma|8830/3
C0334463|T191|SY|C4247|NCI_CDISC|Histiocytoma, Fibrous, Malignant|8830/3
C0334463|T191|SY|C4247|NCI_CDISC|Malignant Fibrous Histiocytoma of Soft Tissue and Bone|8830/3
C0334463|T191|SY|C4247|NCI_CDISC|Malignant Fibrous Histiocytoma of the Soft Tissue and Bone|8830/3
C0334463|T191|SY|C4247|NCI_CDISC|Malignant Fibroxanthoma|8830/3
C0334463|T191|SY|C4247|NCI_CDISC|MFH|8830/3
C0334463|T191|PT|10025556|NCI_CTEP-SDC|Malignant fibrous histiocytoma|8830/3
C0334463|T191|PT|CDR0000349461|NCI_NCI-GLOSS|malignant fibrous cytoma|8830/3
C0334463|T191|PT|CDR0000046174|NCI_NCI-GLOSS|malignant fibrous histiocytoma|8830/3
C0334463|T191|PT|BBGF.|RCD|Malignant fibrous histiocytoma|8830/3
C0334463|T191|IS|X77oV|RCD|Malignant fibroxanthoma|8830/3
C0334463|T191|OP|X77oV|RCDSY|Fibroxanthosarcoma|8830/3
C0334463|T191|PT|34360000|SNOMEDCT_US|Fibrous histiocytoma, malignant|8830/3
C0334463|T191|SY|34360000|SNOMEDCT_US|Fibroxanthoma, malignant|8830/3
C0334463|T191|SY|34360000|SNOMEDCT_US|Malignant fibrous histiocytoma|8830/3
C0334463|T191|PT|443439001|SNOMEDCT_US|Malignant fibrous histiocytoma|8830/3
C0334463|T191|SY|34360000|SNOMEDCT_US|Malignant fibroxanthoma|8830/3
C0334463|T191|SY|34360000|SNOMEDCT_US|Undifferentiated high grade pleomorphic sarcoma|8830/3
C1509147|T191|ET|0000004543|AOD|histiocytoma|8831/0
C1509147|T191|PT|0028796|CCPSS|HISTIOCYTOMA|8831/0
C1509147|T191|PT|0000057998|CHV|histiocytoma|8831/0
C1509147|T191|PT|NOCODE|COSTAR|Histiocytoma|8831/0
C1509147|T191|PT|2004-1029|CSP|histiocytoma|8831/0
C1509147|T191|PT|HP:0012315|HPO|Histiocytoma|8831/0
C1509147|T191|LLT|10020115|MDR|Histiocytoma|8831/0
C1509147|T191|MH|D051642|MSH|Histiocytoma|8831/0
C1509147|T191|PM|D051642|MSH|Histiocytomas|8831/0
C1266125|T191|PN|NOCODE|MTH|Deep histiocytoma|8831/0
C1509147|T191|PN|NOCODE|MTH|Histiocytoma|8831/0
C1266125|T191|SY|C6492|NCI|Benign Deep Fibrous Histiocytoma|8831/0
C1266125|T191|PT|C6492|NCI|Deep Benign Fibrous Histiocytoma|8831/0
C1509147|T191|PT|C35765|NCI|Histiocytoma|8831/0
C1509147|T191|PT|Xa99o|RCD|Histiocytoma|8831/0
C1266125|T191|SY|128741006|SNOMEDCT_US|Deep benign fibrous histiocytoma|8831/0
C1266125|T191|PT|128741006|SNOMEDCT_US|Deep histiocytoma|8831/0
C1509147|T191|SY|128741006|SNOMEDCT_US|Histiocytoma|8831/0
C1509147|T191|OAP|154614002|SNOMEDCT_US|Histiocytoma|8831/0
C1509147|T191|PT|302843004|SNOMEDCT_US|Histiocytoma|8831/0
C1509147|T191|OAP|189773000|SNOMEDCT_US|Histiocytoma|8831/0
C1509147|T191|OF|154614002|SNOMEDCT_US|Histiocytoma|8831/0
C1509147|T191|OF|189773000|SNOMEDCT_US|Histiocytoma|8831/0
C1509147|T191|IS|72079004|SNOMEDCT_US|Histiocytoma, NOS|8831/0
C1266125|T191|SY|128741006|SNOMEDCT_US|Juvenile histiocytoma|8831/0
C0002991|T191|PT|0058687|CCPSS|DERMATOFIBROMA|8832/0
C0002991|T191|SY|0000001175|CHV|cutaneous histiocytoma|8832/0
C0002991|T191|SY|0000001175|CHV|dermatofibroma|8832/0
C0002991|T191|SY|0000001175|CHV|dermatofibromas|8832/0
C0002991|T191|PT|0000001175|CHV|histiocytoma|8832/0
C0002991|T191|SY|0000001175|CHV|histiocytomas|8832/0
C0002991|T191|SY|0000001175|CHV|pleomorphic fibroma|8832/0
C0002991|T191|SY|0000001175|CHV|sclerosing hemangioma|8832/0
C0002991|T191|PT|U000182|COSTAR|DERMATOFIBROMA|8832/0
C0002991|T191|ET|2004-1029|CSP|dermatofibroma|8832/0
C0002991|T191|PTN|S79005|ICPC2P|dermatofibroma|8832/0
C0002991|T191|PT|S79005|ICPC2P|Dermatofibroma|8832/0
C0002991|T191|PT|sh89006247|LCH_NW|Dermatofibroma|8832/0
C0002991|T191|LLT|10012494|MDR|Dermatofibroma|8832/0
C1334455|T191|LLT|10081106|MDR|Sclerosing pneumocytoma|8832/0
C1334455|T191|PT|10081106|MDR|Sclerosing pneumocytoma|8832/0
C0002991|T191|ET|D018219|MSH|Angioma, Sclerosing|8832/0
C0002991|T191|PM|D018219|MSH|Angiomas, Sclerosing|8832/0
C0002991|T191|PM|D018219|MSH|Cutaneous Histiocytoma|8832/0
C0002991|T191|PM|D018219|MSH|Cutaneous Histiocytomas|8832/0
C0002991|T191|PEP|D018219|MSH|Dermatofibroma|8832/0
C0002991|T191|PM|D018219|MSH|Dermatofibromas|8832/0
C1334455|T191|DEV|D047868|MSH|HEMANGIOMA SCLEROSING PULM|8832/0
C0002991|T191|ET|D018219|MSH|Hemangioma, Sclerosing|8832/0
C1334455|T191|ET|D047868|MSH|Hemangioma, Sclerosing, Pulmonary|8832/0
C0002991|T191|PM|D018219|MSH|Hemangiomas, Sclerosing|8832/0
C0002991|T191|ET|D018219|MSH|Histiocytoma, Cutaneous|8832/0
C0002991|T191|PM|D018219|MSH|Histiocytomas, Cutaneous|8832/0
C1334455|T191|ET|D047868|MSH|Lung Sclerosing Hemangioma|8832/0
C1334455|T191|PM|D047868|MSH|Lung Sclerosing Hemangiomas|8832/0
C1334455|T191|DEV|D047868|MSH|PULM SCLEROSING HEMANGIOMA|8832/0
C1334455|T191|MH|D047868|MSH|Pulmonary Sclerosing Hemangioma|8832/0
C1334455|T191|PM|D047868|MSH|Pulmonary Sclerosing Hemangiomas|8832/0
C0002991|T191|PM|D018219|MSH|Sclerosing Angioma|8832/0
C0002991|T191|PM|D018219|MSH|Sclerosing Angiomas|8832/0
C0002991|T191|PM|D018219|MSH|Sclerosing Hemangioma|8832/0
C1334455|T191|ET|D047868|MSH|Sclerosing Hemangioma of the Lung|8832/0
C1334455|T191|ET|D047868|MSH|Sclerosing Hemangioma, Lung|8832/0
C1334455|T191|PM|D047868|MSH|Sclerosing Hemangioma, Pulmonary|8832/0
C0002991|T191|PM|D018219|MSH|Sclerosing Hemangiomas|8832/0
C1334455|T191|PM|D047868|MSH|Sclerosing Hemangiomas, Lung|8832/0
C1334455|T191|PM|D047868|MSH|Sclerosing Hemangiomas, Pulmonary|8832/0
C0002991|T191|PN|NOCODE|MTH|Cutaneous Fibrous Histiocytoma|8832/0
C0002991|T191|SY|C6801|NCI|Benign Cutaneous Fibrous Histiocytoma|8832/0
C0002991|T191|SY|C6801|NCI|Benign Fibrous Cutaneous Histiocytoma|8832/0
C0002991|T191|SY|C6801|NCI|Benign Fibrous Histiocytoma of Skin|8832/0
C0002991|T191|SY|C6801|NCI|Benign Fibrous Histiocytoma of the Skin|8832/0
C0002991|T191|SY|C6801|NCI|Benign Skin Fibrous Histiocytoma|8832/0
C0002991|T191|PT|C6801|NCI|Cutaneous Fibrous Histiocytoma|8832/0
C0002991|T191|SY|C6801|NCI|Dermatofibroma|8832/0
C0002991|T191|SY|C6801|NCI|Fibrous Histiocytoma of Skin|8832/0
C0002991|T191|SY|C6801|NCI|Fibrous Histiocytoma of the Skin|8832/0
C1334455|T191|SY|C5656|NCI|Lung Sclerosing Angioma|8832/0
C1334455|T191|SY|C5656|NCI|Lung Sclerosing Hemangioma|8832/0
C1334455|T191|SY|C5656|NCI|Pneumocytoma|8832/0
C1334455|T191|SY|C5656|NCI|Sclerosing Angioma of Lung|8832/0
C1334455|T191|SY|C5656|NCI|Sclerosing Angioma of the Lung|8832/0
C1334455|T191|SY|C5656|NCI|Sclerosing Hemangioma of Lung|8832/0
C1334455|T191|SY|C5656|NCI|Sclerosing Hemangioma of the Lung|8832/0
C1334455|T191|PT|C5656|NCI|Sclerosing Pneumocytoma|8832/0
C0002991|T191|SY|Xa99o|RCD|Dermatofibroma|8832/0
C0002991|T191|SY|X50K5|RCD|Dermatofibroma lenticulare|8832/0
C0002991|T191|PT|X78Tj|RCD|Fibrous histiocytoma of skin|8832/0
C0002991|T191|OP|X78Tl|RCD|Fibrous xanthoma of skin|8832/0
C0002991|T191|PT|Xa0DA|RCD|Sclerosing angioma|8832/0
C0002991|T191|SY|Xa99o|RCDSY|Dermatofibroma NOS|8832/0
C0002991|T191|SY|254750001|SNOMEDCT_US|Benign fibrous histiocytoma of skin|8832/0
C0002991|T191|OAP|403997008|SNOMEDCT_US|Cutaneous histiocytoma|8832/0
C0002991|T191|SY|427186000|SNOMEDCT_US|Cutaneous histiocytoma|8832/0
C0002991|T191|SY|72079004|SNOMEDCT_US|Cutaneous histiocytoma|8832/0
C0002991|T191|PT|72079004|SNOMEDCT_US|Dermatofibroma|8832/0
C0002991|T191|OAS|189051001|SNOMEDCT_US|Dermatofibroma|8832/0
C0002991|T191|SY|302843004|SNOMEDCT_US|Dermatofibroma|8832/0
C0002991|T191|PT|427186000|SNOMEDCT_US|Dermatofibroma|8832/0
C0002991|T191|SY|72079004|SNOMEDCT_US|Dermatofibroma lenticulare|8832/0
C3164179|T191|PT|448295005|SNOMEDCT_US|Dermatofibroma with monster cells|8832/0
C0002991|T191|SY|72079004|SNOMEDCT_US|Dermatofibroma, no ICD-O subtype|8832/0
C0002991|T191|SY|72079004|SNOMEDCT_US|Dermatofibroma, no International Classification of Diseases for Oncology subtype|8832/0
C0002991|T191|IS|72079004|SNOMEDCT_US|Dermatofibroma, NOS|8832/0
C0002991|T191|PT|254750001|SNOMEDCT_US|Fibrous histiocytoma of skin|8832/0
C0002991|T191|OAP|254753004|SNOMEDCT_US|Fibrous xanthoma of skin|8832/0
C0002991|T191|SY|254750001|SNOMEDCT_US|Fibrous xanthoma of skin|8832/0
C0002991|T191|IS|403997008|SNOMEDCT_US|Pleomorphic fibroma|8832/0
C0002991|T191|PT|448015002|SNOMEDCT_US|Pleomorphic fibroma|8832/0
C1334455|T191|SYGB|707365008|SNOMEDCT_US|Pulmonary sclerosing haemangioma|8832/0
C1334455|T191|SY|707365008|SNOMEDCT_US|Pulmonary sclerosing hemangioma|8832/0
C0002991|T191|PT|134302009|SNOMEDCT_US|Sclerosing angioma|8832/0
C0002991|T191|SY|403999006|SNOMEDCT_US|Sclerosing angioma|8832/0
C0002991|T191|PT|403999006|SNOMEDCT_US|Sclerosing angioma of skin|8832/0
C1334455|T191|PTGB|707365008|SNOMEDCT_US|Sclerosing haemangioma of lung|8832/0
C1334455|T191|PT|707365008|SNOMEDCT_US|Sclerosing hemangioma of lung|8832/0
C1334455|T191|PT|725967000|SNOMEDCT_US|Sclerosing pneumocytoma|8832/0
C0002991|T191|SY|427186000|SNOMEDCT_US|Subepidermal nodular fibrosis|8832/0
C0392784|T191|PT|0000032172|CHV|dermatofibrosarcoma protuberans|8832/1
C0392784|T191|SY|0000032172|CHV|dermatofibrosarcomas protuberans|8832/1
C0392784|T191|PT|MTHU022575|ICPC2ICD10ENG|dermatofibrosarcoma; protuberans|8832/1
C0392784|T191|PT|MTHU062206|ICPC2ICD10ENG|protuberans; dermatofibrosarcoma|8832/1
C0392784|T191|PT|10057070|MDR|Dermatofibrosarcoma protuberans|8832/1
C0392784|T191|LLT|10057070|MDR|Dermatofibrosarcoma protuberans|8832/1
C0392784|T191|PT|355123|MEDCIN|Dermatofibrosarcoma protuberans|8832/1
C0392784|T191|SY|355123|MEDCIN|soft tissue malignant neoplasm dermatofibrosarcoma protuberans|8832/1
C0392784|T191|PN|NOCODE|MTH|Dermatofibrosarcoma Protuberans|8832/1
C0392784|T191|SY|C4683|NCI|Dermatofibrosarcoma|8832/1
C0392784|T191|PT|C4683|NCI|Dermatofibrosarcoma Protuberans|8832/1
C0392784|T191|AB|C4683|NCI|DFSP|8832/1
C0392784|T191|PT|10057043|NCI_CTEP-SDC|Dermatofibrosarcoma|8832/1
C0392784|T191|DN|C4683|NCI_CTRP|Dermatofibrosarcoma Protuberans|8832/1
C0392784|T191|PT|CDR0000044276|NCI_NCI-GLOSS|dermatofibrosarcoma protuberans|8832/1
C0392784|T191|PT|CDR0000474442|PDQ|dermatofibrosarcoma protuberans|8832/1
C0392784|T191|AB|CDR0000474442|PDQ|DFSP|8832/1
C0392784|T191|AB|Xa0D9|RCD|Dermatofibrosarcom protuberans|8832/1
C0392784|T191|PT|Xa0D9|RCD|Dermatofibrosarcoma protuberans|8832/1
C0392784|T191|AB|Xa0D9|RCD|DFSP - Dermatofibrosarc protru|8832/1
C0392784|T191|SY|Xa0D9|RCD|DFSP - Dermatofibrosarcoma protruberans|8832/1
C0392784|T191|OP|BBGL.|RCDSY|Dermatofibroma protuberans|8832/1
C0392784|T191|SY|276799004|SNOMEDCT_US|Dermatofibrosarcoma|8832/1
C0392784|T191|SY|76594008|SNOMEDCT_US|Dermatofibrosarcoma|8832/1
C0392784|T191|PT|76594008|SNOMEDCT_US|Dermatofibrosarcoma protuberans|8832/1
C0392784|T191|OAP|188140006|SNOMEDCT_US|Dermatofibrosarcoma protuberans|8832/1
C0392784|T191|PT|276799004|SNOMEDCT_US|Dermatofibrosarcoma protuberans|8832/1
C0392784|T191|OF|188140006|SNOMEDCT_US|Dermatofibrosarcoma protuberans|8832/1
C0392784|T191|IS|76594008|SNOMEDCT_US|Dermatofibrosarcoma protuberans, NOS|8832/1
C0392784|T191|SY|76594008|SNOMEDCT_US|Dermatofibrosarcoma, no ICD-O subtype|8832/1
C0392784|T191|SY|76594008|SNOMEDCT_US|Dermatofibrosarcoma, no International Classification of Diseases for Oncology subtype|8832/1
C0392784|T191|IS|76594008|SNOMEDCT_US|Dermatofibrosarcoma, NOS|8832/1
C0392784|T191|IS|276799004|SNOMEDCT_US|DFSP - Dermatofibrosarcoma protruberans|8832/1
C0392784|T191|SY|276799004|SNOMEDCT_US|DFSP - dermatofibrosarcoma protuberans|8832/1
C0392784|T191|PT|0000032172|CHV|dermatofibrosarcoma protuberans|8832/3
C0392784|T191|SY|0000032172|CHV|dermatofibrosarcomas protuberans|8832/3
C0392784|T191|PT|MTHU022575|ICPC2ICD10ENG|dermatofibrosarcoma; protuberans|8832/3
C0392784|T191|PT|MTHU062206|ICPC2ICD10ENG|protuberans; dermatofibrosarcoma|8832/3
C0392784|T191|PT|10057070|MDR|Dermatofibrosarcoma protuberans|8832/3
C0392784|T191|LLT|10057070|MDR|Dermatofibrosarcoma protuberans|8832/3
C3665732|T191|LLT|10073574|MDR|Dermatofibrosarcoma protuberans metastatic|8832/3
C3665732|T191|PT|10073574|MDR|Dermatofibrosarcoma protuberans metastatic|8832/3
C0392784|T191|PT|355123|MEDCIN|Dermatofibrosarcoma protuberans|8832/3
C0392784|T191|SY|355123|MEDCIN|soft tissue malignant neoplasm dermatofibrosarcoma protuberans|8832/3
C3665732|T191|PM|D018223|MSH|Dermatofibrosarcoma Protuberan, Fibrosarcomatous|8832/3
C3665732|T191|PM|D018223|MSH|Dermatofibrosarcoma Protuberan, Metastatic|8832/3
C3665732|T191|ET|D018223|MSH|Dermatofibrosarcoma Protuberans, Fibrosarcomatous|8832/3
C3665732|T191|PM|D018223|MSH|Dermatofibrosarcoma Protuberans, Metastatic|8832/3
C3665732|T191|ET|D018223|MSH|DFSP, Fibrosarcomatous|8832/3
C3665732|T191|PM|D018223|MSH|DFSPs, Fibrosarcomatous|8832/3
C3665732|T191|PM|D018223|MSH|Fibrosarcomatous Dermatofibrosarcoma Protuberan|8832/3
C3665732|T191|ET|D018223|MSH|Fibrosarcomatous Dermatofibrosarcoma Protuberans|8832/3
C3665732|T191|PM|D018223|MSH|Fibrosarcomatous DFSP|8832/3
C3665732|T191|PM|D018223|MSH|Fibrosarcomatous DFSPs|8832/3
C3665732|T191|ET|D018223|MSH|FS-DFSP|8832/3
C3665732|T191|PM|D018223|MSH|Metastatic Dermatofibrosarcoma Protuberan|8832/3
C3665732|T191|PEP|D018223|MSH|Metastatic Dermatofibrosarcoma Protuberans|8832/3
C3665732|T191|PM|D018223|MSH|Protuberan, Fibrosarcomatous Dermatofibrosarcoma|8832/3
C3665732|T191|PM|D018223|MSH|Protuberan, Metastatic Dermatofibrosarcoma|8832/3
C3665732|T191|PM|D018223|MSH|Protuberans, Fibrosarcomatous Dermatofibrosarcoma|8832/3
C3665732|T191|PM|D018223|MSH|Protuberans, Metastatic Dermatofibrosarcoma|8832/3
C0392784|T191|PN|NOCODE|MTH|Dermatofibrosarcoma Protuberans|8832/3
C0392784|T191|SY|C4683|NCI|Dermatofibrosarcoma|8832/3
C0392784|T191|PT|C4683|NCI|Dermatofibrosarcoma Protuberans|8832/3
C0392784|T191|AB|C4683|NCI|DFSP|8832/3
C3665732|T191|PT|C27547|NCI|Fibrosarcomatous Dermatofibrosarcoma Protuberans|8832/3
C0392784|T191|PT|10057043|NCI_CTEP-SDC|Dermatofibrosarcoma|8832/3
C0392784|T191|DN|C4683|NCI_CTRP|Dermatofibrosarcoma Protuberans|8832/3
C0392784|T191|PT|CDR0000044276|NCI_NCI-GLOSS|dermatofibrosarcoma protuberans|8832/3
C0392784|T191|PT|CDR0000474442|PDQ|dermatofibrosarcoma protuberans|8832/3
C0392784|T191|AB|CDR0000474442|PDQ|DFSP|8832/3
C0392784|T191|AB|Xa0D9|RCD|Dermatofibrosarcom protuberans|8832/3
C0392784|T191|PT|Xa0D9|RCD|Dermatofibrosarcoma protuberans|8832/3
C0392784|T191|AB|Xa0D9|RCD|DFSP - Dermatofibrosarc protru|8832/3
C0392784|T191|SY|Xa0D9|RCD|DFSP - Dermatofibrosarcoma protruberans|8832/3
C0392784|T191|OP|BBGL.|RCDSY|Dermatofibroma protuberans|8832/3
C0392784|T191|SY|276799004|SNOMEDCT_US|Dermatofibrosarcoma|8832/3
C0392784|T191|SY|76594008|SNOMEDCT_US|Dermatofibrosarcoma|8832/3
C0392784|T191|PT|76594008|SNOMEDCT_US|Dermatofibrosarcoma protuberans|8832/3
C0392784|T191|OAP|188140006|SNOMEDCT_US|Dermatofibrosarcoma protuberans|8832/3
C0392784|T191|PT|276799004|SNOMEDCT_US|Dermatofibrosarcoma protuberans|8832/3
C0392784|T191|OF|188140006|SNOMEDCT_US|Dermatofibrosarcoma protuberans|8832/3
C0392784|T191|IS|76594008|SNOMEDCT_US|Dermatofibrosarcoma protuberans, NOS|8832/3
C0392784|T191|SY|76594008|SNOMEDCT_US|Dermatofibrosarcoma, no ICD-O subtype|8832/3
C0392784|T191|SY|76594008|SNOMEDCT_US|Dermatofibrosarcoma, no International Classification of Diseases for Oncology subtype|8832/3
C0392784|T191|IS|76594008|SNOMEDCT_US|Dermatofibrosarcoma, NOS|8832/3
C0392784|T191|IS|276799004|SNOMEDCT_US|DFSP - Dermatofibrosarcoma protruberans|8832/3
C0392784|T191|SY|276799004|SNOMEDCT_US|DFSP - dermatofibrosarcoma protuberans|8832/3
C3665732|T191|PT|733859002|SNOMEDCT_US|Fibrosarcomatous dermatofibrosarcoma protuberans|8832/3
C0334464|T191|PT|MTHU022576|ICPC2ICD10ENG|dermatofibrosarcoma; protuberans, pigmented|8833/1
C0334464|T191|PT|MTHU062207|ICPC2ICD10ENG|protuberans; dermatofibrosarcoma, pigmented|8833/1
C0334464|T191|PT|231676|MEDCIN|pigmented dermatofibrosarcoma protuberans of skin|8833/1
C0334464|T191|ET|D018223|MSH|Bednar Tumor|8833/1
C0334464|T191|ET|D018223|MSH|Bednar's Tumor|8833/1
C0334464|T191|PM|D018223|MSH|Bednars Tumor|8833/1
C0334464|T191|PM|D018223|MSH|Dermatofibrosarcoma Protuberan, Pigmented|8833/1
C0334464|T191|PEP|D018223|MSH|Dermatofibrosarcoma Protuberans, Pigmented|8833/1
C0334464|T191|ET|D018223|MSH|DFSP, Pigmented|8833/1
C0334464|T191|PM|D018223|MSH|DFSPs, Pigmented|8833/1
C0334464|T191|PM|D018223|MSH|Pigmented Dermatofibrosarcoma Protuberan|8833/1
C0334464|T191|PM|D018223|MSH|Pigmented Dermatofibrosarcoma Protuberans|8833/1
C0334464|T191|PM|D018223|MSH|Pigmented DFSP|8833/1
C0334464|T191|PM|D018223|MSH|Pigmented DFSPs|8833/1
C0334464|T191|PM|D018223|MSH|Protuberan, Pigmented Dermatofibrosarcoma|8833/1
C0334464|T191|PM|D018223|MSH|Protuberans, Pigmented Dermatofibrosarcoma|8833/1
C0334464|T191|PM|D018223|MSH|Tumor, Bednar|8833/1
C0334464|T191|PM|D018223|MSH|Tumor, Bednar's|8833/1
C0334464|T191|SY|C9430|NCI|Bednar Tumor|8833/1
C0334464|T191|PT|C9430|NCI|Pigmented Dermatofibrosarcoma Protuberans|8833/1
C0334464|T191|SY|X77oW|RCD|Bednar tumour|8833/1
C0334464|T191|AB|X77oW|RCD|Pigm dermatofibrosarc protub|8833/1
C0334464|T191|SY|X77oW|RCD|Pigmented dermatofibrosarcoma|8833/1
C0334464|T191|PT|X77oW|RCD|Pigmented dermatofibrosarcoma protuberans|8833/1
C0334464|T191|AB|X77oW|RCD|Pigmented storif neurofibroma|8833/1
C0334464|T191|SY|X77oW|RCD|Pigmented storiform neurofibroma|8833/1
C0334464|T191|SY|X77oW|RCDAE|Bednar tumor|8833/1
C0334464|T191|OA|BBGP.|RCDSY|Pigmen dermatfibsarc protub|8833/1
C0334464|T191|OP|BBGP.|RCDSY|Pigmented dermatofibrosarcoma protuberans|8833/1
C0334464|T191|SY|398670003|SNOMEDCT_US|Bednar tumor|8833/1
C0334464|T191|OAS|253041002|SNOMEDCT_US|Bednar tumor|8833/1
C0334464|T191|SY|62621002|SNOMEDCT_US|Bednar tumor|8833/1
C0334464|T191|OAS|253041002|SNOMEDCT_US|Bednar tumour|8833/1
C0334464|T191|SYGB|62621002|SNOMEDCT_US|Bednar tumour|8833/1
C0334464|T191|SYGB|398670003|SNOMEDCT_US|Bednar tumour|8833/1
C0334464|T191|SY|398670003|SNOMEDCT_US|Pigmented dermatofibrosarcoma|8833/1
C0334464|T191|OAS|253041002|SNOMEDCT_US|Pigmented dermatofibrosarcoma|8833/1
C0334464|T191|OAP|253041002|SNOMEDCT_US|Pigmented dermatofibrosarcoma protuberans|8833/1
C0334464|T191|PT|62621002|SNOMEDCT_US|Pigmented dermatofibrosarcoma protuberans|8833/1
C0334464|T191|PT|398670003|SNOMEDCT_US|Pigmented dermatofibrosarcoma protuberans of skin|8833/1
C0334464|T191|OAS|253041002|SNOMEDCT_US|Pigmented storiform neurofibroma|8833/1
C0334464|T191|SY|398670003|SNOMEDCT_US|Pigmented storiform neurofibroma|8833/1
C0334464|T191|PT|MTHU022576|ICPC2ICD10ENG|dermatofibrosarcoma; protuberans, pigmented|8833/3
C0334464|T191|PT|MTHU062207|ICPC2ICD10ENG|protuberans; dermatofibrosarcoma, pigmented|8833/3
C0334464|T191|PT|231676|MEDCIN|pigmented dermatofibrosarcoma protuberans of skin|8833/3
C0334464|T191|ET|D018223|MSH|Bednar Tumor|8833/3
C0334464|T191|ET|D018223|MSH|Bednar's Tumor|8833/3
C0334464|T191|PM|D018223|MSH|Bednars Tumor|8833/3
C0334464|T191|PM|D018223|MSH|Dermatofibrosarcoma Protuberan, Pigmented|8833/3
C0334464|T191|PEP|D018223|MSH|Dermatofibrosarcoma Protuberans, Pigmented|8833/3
C0334464|T191|ET|D018223|MSH|DFSP, Pigmented|8833/3
C0334464|T191|PM|D018223|MSH|DFSPs, Pigmented|8833/3
C0334464|T191|PM|D018223|MSH|Pigmented Dermatofibrosarcoma Protuberan|8833/3
C0334464|T191|PM|D018223|MSH|Pigmented Dermatofibrosarcoma Protuberans|8833/3
C0334464|T191|PM|D018223|MSH|Pigmented DFSP|8833/3
C0334464|T191|PM|D018223|MSH|Pigmented DFSPs|8833/3
C0334464|T191|PM|D018223|MSH|Protuberan, Pigmented Dermatofibrosarcoma|8833/3
C0334464|T191|PM|D018223|MSH|Protuberans, Pigmented Dermatofibrosarcoma|8833/3
C0334464|T191|PM|D018223|MSH|Tumor, Bednar|8833/3
C0334464|T191|PM|D018223|MSH|Tumor, Bednar's|8833/3
C0334464|T191|SY|C9430|NCI|Bednar Tumor|8833/3
C0334464|T191|PT|C9430|NCI|Pigmented Dermatofibrosarcoma Protuberans|8833/3
C0334464|T191|SY|X77oW|RCD|Bednar tumour|8833/3
C0334464|T191|AB|X77oW|RCD|Pigm dermatofibrosarc protub|8833/3
C0334464|T191|SY|X77oW|RCD|Pigmented dermatofibrosarcoma|8833/3
C0334464|T191|PT|X77oW|RCD|Pigmented dermatofibrosarcoma protuberans|8833/3
C0334464|T191|AB|X77oW|RCD|Pigmented storif neurofibroma|8833/3
C0334464|T191|SY|X77oW|RCD|Pigmented storiform neurofibroma|8833/3
C0334464|T191|SY|X77oW|RCDAE|Bednar tumor|8833/3
C0334464|T191|OA|BBGP.|RCDSY|Pigmen dermatfibsarc protub|8833/3
C0334464|T191|OP|BBGP.|RCDSY|Pigmented dermatofibrosarcoma protuberans|8833/3
C0334464|T191|OAS|253041002|SNOMEDCT_US|Bednar tumor|8833/3
C0334464|T191|SY|62621002|SNOMEDCT_US|Bednar tumor|8833/3
C0334464|T191|SY|398670003|SNOMEDCT_US|Bednar tumor|8833/3
C0334464|T191|SYGB|62621002|SNOMEDCT_US|Bednar tumour|8833/3
C0334464|T191|SYGB|398670003|SNOMEDCT_US|Bednar tumour|8833/3
C0334464|T191|OAS|253041002|SNOMEDCT_US|Bednar tumour|8833/3
C0334464|T191|OAS|253041002|SNOMEDCT_US|Pigmented dermatofibrosarcoma|8833/3
C0334464|T191|SY|398670003|SNOMEDCT_US|Pigmented dermatofibrosarcoma|8833/3
C0334464|T191|PT|62621002|SNOMEDCT_US|Pigmented dermatofibrosarcoma protuberans|8833/3
C0334464|T191|OAP|253041002|SNOMEDCT_US|Pigmented dermatofibrosarcoma protuberans|8833/3
C0334464|T191|PT|398670003|SNOMEDCT_US|Pigmented dermatofibrosarcoma protuberans of skin|8833/3
C0334464|T191|OAS|253041002|SNOMEDCT_US|Pigmented storiform neurofibroma|8833/3
C0334464|T191|SY|398670003|SNOMEDCT_US|Pigmented storiform neurofibroma|8833/3
C3693482|T191|PT|355131|MEDCIN|Giant cell fibroblastoma of skin|8834/1
C3693482|T191|SY|355131|MEDCIN|skin neoplasm giant cell fibroblastoma|8834/1
C3693482|T191|PM|D018223|MSH|Cell Fibroblastoma, Giant|8834/1
C3693482|T191|PM|D018223|MSH|Cell Fibroblastomas, Giant|8834/1
C3693482|T191|PM|D018223|MSH|Dermatofibrosarcoma Protuberan, Familial|8834/1
C3693482|T191|PM|D018223|MSH|Dermatofibrosarcoma Protuberan, Giant|8834/1
C3693482|T191|ET|D018223|MSH|Dermatofibrosarcoma Protuberans, Familial|8834/1
C3693482|T191|PM|D018223|MSH|Dermatofibrosarcoma Protuberans, Giant|8834/1
C3693482|T191|ET|D018223|MSH|Dermatofibrosarcoma Protuberans, Giant Cell|8834/1
C3693482|T191|ET|D018223|MSH|DFSP, Juvenile|8834/1
C3693482|T191|PM|D018223|MSH|DFSPs, Juvenile|8834/1
C3693482|T191|PM|D018223|MSH|Familial Dermatofibrosarcoma Protuberan|8834/1
C3693482|T191|ET|D018223|MSH|Familial Dermatofibrosarcoma Protuberans|8834/1
C3693482|T191|PM|D018223|MSH|Fibroblastoma, Giant Cell|8834/1
C3693482|T191|PM|D018223|MSH|Fibroblastomas, Giant Cell|8834/1
C3693482|T191|PEP|D018223|MSH|Giant Cell Fibroblastoma|8834/1
C3693482|T191|PM|D018223|MSH|Giant Cell Fibroblastomas|8834/1
C3693482|T191|PM|D018223|MSH|Giant Dermatofibrosarcoma Protuberan|8834/1
C3693482|T191|ET|D018223|MSH|Giant Dermatofibrosarcoma Protuberans|8834/1
C3693482|T191|PM|D018223|MSH|Juvenile DFSP|8834/1
C3693482|T191|PM|D018223|MSH|Juvenile DFSPs|8834/1
C3693482|T191|PM|D018223|MSH|Protuberan, Familial Dermatofibrosarcoma|8834/1
C3693482|T191|PM|D018223|MSH|Protuberan, Giant Dermatofibrosarcoma|8834/1
C3693482|T191|PM|D018223|MSH|Protuberans, Familial Dermatofibrosarcoma|8834/1
C3693482|T191|PM|D018223|MSH|Protuberans, Giant Dermatofibrosarcoma|8834/1
C3693482|T191|PN|NOCODE|MTH|Giant Cell Fibroblastoma|8834/1
C3693482|T191|AB|C4700|NCI|GCF|8834/1
C3693482|T191|PT|C4700|NCI|Giant Cell Fibroblastoma|8834/1
C3693482|T191|PT|CDR0000390282|NCI_NCI-GLOSS|giant cell fibroblastoma|8834/1
C3693482|T191|PT|X50DM|RCD|Giant cell fibroblastoma|8834/1
C3693482|T191|SY|238863004|SNOMEDCT_US|Giant cell fibroblastoma|8834/1
C3693482|T191|PT|128742004|SNOMEDCT_US|Giant cell fibroblastoma|8834/1
C3693482|T191|PT|238863004|SNOMEDCT_US|Giant cell fibroblastoma of skin|8834/1
C1266126|T191|AB|C6493|NCI|PFHT|8835/1
C1266126|T191|SY|C6493|NCI|Plexiform Fibrohistiocytic Neoplasm|8835/1
C1266126|T191|PT|C6493|NCI|Plexiform Fibrohistiocytic Tumor|8835/1
C1266126|T191|PT|128743009|SNOMEDCT_US|Plexiform fibrohistiocytic tumor|8835/1
C1266126|T191|PTGB|128743009|SNOMEDCT_US|Plexiform fibrohistiocytic tumour|8835/1
C1266127|T191|PT|0000056689|CHV|angiomatoid fibrous histiocytoma|8836/1
C1266127|T191|NM|C563181|MSH|Histiocytoma, Angiomatoid Fibrous|8836/1
C1266127|T191|AB|C6494|NCI|AFH|8836/1
C1266127|T191|PT|C6494|NCI|Angiomatoid Fibrous Histiocytoma|8836/1
C1266127|T191|SY|C6494|NCI|Angiomatoid Malignant Fibrous Histiocytoma|8836/1
C1266127|T191|PT|128744003|SNOMEDCT_US|Angiomatoid fibrous histiocytoma|8836/1
C0027149|T191|PT|0024763|CCPSS|MYXOMA|8840/0
C0027149|T191|PT|0000057855|CHV|angiomyxoma|8840/0
C0027149|T191|PT|0000008451|CHV|myxoma|8840/0
C0027149|T191|SY|0000008451|CHV|myxomas|8840/0
C0027149|T191|PT|U003112|LCH|Myxoma|8840/0
C0027149|T191|PT|sh85089453|LCH_NW|Myxoma|8840/0
C0027149|T191|LLT|10076892|MDR|Angiomyxoma|8840/0
C0027149|T191|PT|10076892|MDR|Angiomyxoma|8840/0
C0027149|T191|PT|355060|MEDCIN|Angiomyxoma|8840/0
C0027149|T191|SY|355060|MEDCIN|neoplasm of uncertain behavior angiomyxoma|8840/0
C0027149|T191|ET|D009232|MSH|Angiomyxoma|8840/0
C0027149|T191|PM|D009232|MSH|Angiomyxomas|8840/0
C0027149|T191|MH|D009232|MSH|Myxoma|8840/0
C0027149|T191|PM|D009232|MSH|Myxomas|8840/0
C0027149|T191|PT|C3254|NCI|Angiomyxoma|8840/0
C0027149|T191|PT|C6577|NCI|Myxoma|8840/0
C0027149|T191|PT|C6577|NCI_CDISC|MYXOMA, BENIGN|8840/0
C0027149|T191|OP|BBHZ.|RCDSY|Angiomyxoma|8840/0
C0027149|T191|OP|BBH0.|RCDSY|Myxoma NOS|8840/0
C0027149|T191|PT|404083008|SNOMEDCT_US|Angiomyxoma|8840/0
C0027149|T191|PT|57723004|SNOMEDCT_US|Angiomyxoma|8840/0
C0027149|T191|PT|404082003|SNOMEDCT_US|Myxoma|8840/0
C0027149|T191|PT|39143003|SNOMEDCT_US|Myxoma|8840/0
C0027149|T191|IS|39143003|SNOMEDCT_US|Myxoma, NOS|8840/0
C0027155|T191|ET|0000004532|AOD|myxosarcoma|8840/3
C1275282|T191|PT|355173|MEDCIN|Low-grade fibromyxoid sarcoma|8840/3
C1275282|T191|SY|355173|MEDCIN|malignant neoplasm sarcoma low-grade fibromyxoid|8840/3
C0027155|T191|PT|215623|MEDCIN|myxosarcoma|8840/3
C0027155|T191|MH|D009236|MSH|Myxosarcoma|8840/3
C0027155|T191|PM|D009236|MSH|Myxosarcomas|8840/3
C1710026|T191|PN|NOCODE|MTH|Sclerosing Epithelioid Fibrosarcoma|8840/3
C1275282|T191|PT|C45202|NCI|Low Grade Fibromyxoid Sarcoma|8840/3
C0027155|T191|PT|C3255|NCI|Myxosarcoma|8840/3
C1710026|T191|PT|C49027|NCI|Sclerosing Epithelioid Fibrosarcoma|8840/3
C1710026|T191|AB|C49027|NCI|SEF|8840/3
C0027155|T191|PT|C3255|NCI_CDISC|MYXOSARCOMA, MALIGNANT|8840/3
C0027155|T191|OP|BBH1.|RCDSY|Myxosarcoma|8840/3
C1275282|T191|PT|703617004|SNOMEDCT_US|Low grade fibromyxoid sarcoma|8840/3
C1275282|T191|PT|404088004|SNOMEDCT_US|Low-grade fibromyxoid sarcoma|8840/3
C0027155|T191|PT|28351005|SNOMEDCT_US|Myxosarcoma|8840/3
C1710026|T191|PT|703618009|SNOMEDCT_US|Sclerosing epithelioid fibrosarcoma|8840/3
C0027149|T191|PT|0024763|CCPSS|MYXOMA|8841/0
C0027149|T191|PT|0000057855|CHV|angiomyxoma|8841/0
C0027149|T191|PT|0000008451|CHV|myxoma|8841/0
C0027149|T191|SY|0000008451|CHV|myxomas|8841/0
C0027149|T191|PT|U003112|LCH|Myxoma|8841/0
C0027149|T191|PT|sh85089453|LCH_NW|Myxoma|8841/0
C0027149|T191|LLT|10076892|MDR|Angiomyxoma|8841/0
C0027149|T191|PT|10076892|MDR|Angiomyxoma|8841/0
C0027149|T191|PT|355060|MEDCIN|Angiomyxoma|8841/0
C0027149|T191|SY|355060|MEDCIN|neoplasm of uncertain behavior angiomyxoma|8841/0
C0027149|T191|ET|D009232|MSH|Angiomyxoma|8841/0
C0027149|T191|PM|D009232|MSH|Angiomyxomas|8841/0
C0027149|T191|MH|D009232|MSH|Myxoma|8841/0
C0027149|T191|PM|D009232|MSH|Myxomas|8841/0
C0027149|T191|PT|C3254|NCI|Angiomyxoma|8841/0
C0027149|T191|PT|C6577|NCI|Myxoma|8841/0
C0027149|T191|PT|C6577|NCI_CDISC|MYXOMA, BENIGN|8841/0
C0027149|T191|OP|BBHZ.|RCDSY|Angiomyxoma|8841/0
C0027149|T191|OP|BBH0.|RCDSY|Myxoma NOS|8841/0
C0027149|T191|PT|57723004|SNOMEDCT_US|Angiomyxoma|8841/0
C0027149|T191|PT|404083008|SNOMEDCT_US|Angiomyxoma|8841/0
C0027149|T191|PT|404082003|SNOMEDCT_US|Myxoma|8841/0
C0027149|T191|PT|39143003|SNOMEDCT_US|Myxoma|8841/0
C0027149|T191|IS|39143003|SNOMEDCT_US|Myxoma, NOS|8841/0
C0027149|T191|PT|0024763|CCPSS|MYXOMA|8841/1
C0027149|T191|PT|0000057855|CHV|angiomyxoma|8841/1
C0027149|T191|PT|0000008451|CHV|myxoma|8841/1
C0027149|T191|SY|0000008451|CHV|myxomas|8841/1
C0027149|T191|PT|U003112|LCH|Myxoma|8841/1
C0027149|T191|PT|sh85089453|LCH_NW|Myxoma|8841/1
C0027149|T191|LLT|10076892|MDR|Angiomyxoma|8841/1
C0027149|T191|PT|10076892|MDR|Angiomyxoma|8841/1
C0027149|T191|PT|355060|MEDCIN|Angiomyxoma|8841/1
C0027149|T191|SY|355060|MEDCIN|neoplasm of uncertain behavior angiomyxoma|8841/1
C0027149|T191|ET|D009232|MSH|Angiomyxoma|8841/1
C0027149|T191|PM|D009232|MSH|Angiomyxomas|8841/1
C0027149|T191|MH|D009232|MSH|Myxoma|8841/1
C0027149|T191|PM|D009232|MSH|Myxomas|8841/1
C0027149|T191|PT|C3254|NCI|Angiomyxoma|8841/1
C0027149|T191|PT|C6577|NCI|Myxoma|8841/1
C0027149|T191|PT|C6577|NCI_CDISC|MYXOMA, BENIGN|8841/1
C0027149|T191|OP|BBHZ.|RCDSY|Angiomyxoma|8841/1
C0027149|T191|OP|BBH0.|RCDSY|Myxoma NOS|8841/1
C0027149|T191|PT|404083008|SNOMEDCT_US|Angiomyxoma|8841/1
C0027149|T191|PT|57723004|SNOMEDCT_US|Angiomyxoma|8841/1
C0027149|T191|PT|404082003|SNOMEDCT_US|Myxoma|8841/1
C0027149|T191|PT|39143003|SNOMEDCT_US|Myxoma|8841/1
C0027149|T191|IS|39143003|SNOMEDCT_US|Myxoma, NOS|8841/1
C1266128|T191|AB|C6582|NCI|OFMT|8842/0
C1266128|T191|SY|C6582|NCI|Ossifying Fibromyxoid Neoplasm|8842/0
C1266128|T191|PT|C6582|NCI|Ossifying Fibromyxoid Tumor|8842/0
C1266128|T191|SY|C6582|NCI|Ossifying Fibromyxoma|8842/0
C1266128|T191|PT|128745002|SNOMEDCT_US|Ossifying fibromyxoid tumor|8842/0
C1266128|T191|PT|404076001|SNOMEDCT_US|Ossifying fibromyxoid tumor|8842/0
C1266128|T191|PTGB|404076001|SNOMEDCT_US|Ossifying fibromyxoid tumour|8842/0
C1266128|T191|PTGB|128745002|SNOMEDCT_US|Ossifying fibromyxoid tumour|8842/0
C3839955|T191|PT|C121774|NCI|Malignant Ossifying Fibromyxoid Tumor|8842/3
C3839955|T191|PT|703631004|SNOMEDCT_US|Ossifying fibromyxoid tumor, malignant|8842/3
C3839955|T191|PTGB|703631004|SNOMEDCT_US|Ossifying fibromyxoid tumour, malignant|8842/3
C0023798|T191|PT|BI00600|BI|lipoma|8850/0
C0023798|T191|PT|1011468|CCPSS|LIPOMA|8850/0
C0023798|T191|PT|0000007464|CHV|fatty tumor|8850/0
C0023798|T191|SY|0000007464|CHV|fatty tumors|8850/0
C0023798|T191|SY|0000007464|CHV|lipoma|8850/0
C0023798|T191|SY|0000007464|CHV|lipoma nos|8850/0
C0023798|T191|SY|0000007464|CHV|lipomas|8850/0
C0023798|T191|SY|0000007464|CHV|lipomata|8850/0
C0023798|T191|PT|454|COSTAR|LIPOMA|8850/0
C0023798|T191|ET|0729-5644|CSP|lipoma|8850/0
C0023798|T191|ET|2008-3809|CSP|lipoma|8850/0
C0023798|T191|GT|NEOPL|CST|LIPOMA|8850/0
C0023798|T191|SY|HP:0012032|HPO|Fatty lump|8850/0
C0023798|T191|PT|HP:0012032|HPO|Lipoma|8850/0
C0023798|T191|ET|HP:0001012|HPO|Lipomas|8850/0
C0023798|T191|SY|HP:0012032|HPO|Noncancerous fatty lump|8850/0
C0023798|T191|ET|D17.9|ICD10CM|Lipoma NOS|8850/0
C0023798|T191|HT|214|ICD9CM|Lipoma|8850/0
C0023798|T191|AB|214.9|ICD9CM|Lipoma NOS|8850/0
C0023798|T191|PT|214.9|ICD9CM|Lipoma, unspecified site|8850/0
C0023798|T191|PT|S78|ICPC|Lipoma|8850/0
C0023798|T191|AB|S78|ICPC2EENG|Lipoma|8850/0
C0023798|T191|PT|S78|ICPC2EENG|Lipoma|8850/0
C0023798|T191|PT|MTHU045584|ICPC2ICD10ENG|lipoma|8850/0
C0023798|T191|LA|LA26514-2|LNC|Lipoma, NOS|8850/0
C0023798|T191|LLT|10024612|MDR|Lipoma|8850/0
C0023798|T191|PT|10024612|MDR|Lipoma|8850/0
C0023798|T191|LLT|10024615|MDR|Lipoma NOS|8850/0
C0023798|T191|LLT|10024623|MDR|Lipoma, unspecified site|8850/0
C0023798|T191|ET|D008067|MSH|Fatty Tumor|8850/0
C0023798|T191|PM|D008067|MSH|Fatty Tumors|8850/0
C0023798|T191|MH|D008067|MSH|Lipoma|8850/0
C0023798|T191|PM|D008067|MSH|Lipomas|8850/0
C0023798|T191|ET|D008067|MSH|Lipomata|8850/0
C0023798|T191|PM|D008067|MSH|Lipomatas|8850/0
C0023798|T191|PM|D008067|MSH|Tumor, Fatty|8850/0
C0023798|T191|PM|D008067|MSH|Tumors, Fatty|8850/0
C0023798|T191|PN|NOCODE|MTH|Lipoma|8850/0
C0023798|T191|PT|C3192|NCI|Lipoma|8850/0
C1336744|T191|PT|C6452|NCI|Thymolipoma|8850/0
C1336744|T191|SY|C6452|NCI|Thymolipomatous Hamartoma|8850/0
C0023798|T191|PT|C3192|NCI_CDISC|LIPOMA, BENIGN|8850/0
C0023798|T191|PT|C3192|NCI_CPTAC|Lipoma|8850/0
C0023798|T191|PT|CDR0000454795|NCI_NCI-GLOSS|lipoma|8850/0
C0023798|T191|PT|C3192|NCI_NICHD|Lipoma|8850/0
C0023798|T191|PT|B74..|RCD|Lipoma|8850/0
C0431102|T191|PT|Xa99q|RCD|Lipoma morphology|8850/0
C0023798|T191|OP|B74z.|RCD|Lipoma NOS|8850/0
C0023798|T191|OP|BBJ0.|RCDSY|Lipoma NOS|8850/0
C0023798|T191|OF|154612003|SNOMEDCT_US|Lipoma|8850/0
C0023798|T191|SY|93163002|SNOMEDCT_US|Lipoma|8850/0
C0023798|T191|OAP|154612003|SNOMEDCT_US|Lipoma|8850/0
C0023798|T191|PT|46720004|SNOMEDCT_US|Lipoma|8850/0
C0431102|T191|PT|134328007|SNOMEDCT_US|Lipoma morphology|8850/0
C0023798|T191|OAP|189018005|SNOMEDCT_US|Lipoma NOS|8850/0
C0023798|T191|IS|93163002|SNOMEDCT_US|Lipoma of unspecified body site|8850/0
C0023798|T191|SY|46720004|SNOMEDCT_US|Lipoma, no ICD-O subtype|8850/0
C0023798|T191|SY|46720004|SNOMEDCT_US|Lipoma, no International Classification of Diseases for Oncology subtype|8850/0
C0023798|T191|IS|46720004|SNOMEDCT_US|Lipoma, NOS|8850/0
C2959648|T191|PT|447061000|SNOMEDCT_US|Osteolipoma|8850/0
C1336744|T191|PT|447137005|SNOMEDCT_US|Thymolipoma|8850/0
C0023798|T191|PT|1067|WHO|LIPOMA|8850/0
C1266129|T191|PN|NOCODE|MTH|Atypical Lipoma|8850/1
C1266129|T191|AB|C6505|NCI|ALT|8850/1
C1266129|T191|SY|C6505|NCI|Atypical Lipoma|8850/1
C1266129|T191|PT|C6505|NCI|Atypical Lipomatous Tumor|8850/1
C1266129|T191|SY|C6505|NCI|Lipoma-Like Liposarcoma|8850/1
C1266129|T191|SY|C6505|NCI|Superficial Well Differentiated Liposarcoma|8850/1
C1266129|T191|SY|C6505|NCI|Well Differentiated Liposarcoma|8850/1
C1266129|T191|SY|C6505|NCI|Well Differentiated Liposarcoma of Superficial Soft Tissue|8850/1
C1266129|T191|SY|116063003|SNOMEDCT_US|Atypical lipoma|8850/1
C1266129|T191|PT|116063003|SNOMEDCT_US|Atypical lipomatous tumor|8850/1
C1266129|T191|PTGB|116063003|SNOMEDCT_US|Atypical lipomatous tumour|8850/1
C1266129|T191|SY|28655007|SNOMEDCT_US|Lipoma-like liposarcoma|8850/1
C1266129|T191|IS|116063003|SNOMEDCT_US|Superficial well differentated liposarcoma|8850/1
C1266129|T191|IS|116063003|SNOMEDCT_US|Superficial well differentiated liposarcoma|8850/1
C1266129|T191|IS|116063003|SNOMEDCT_US|Well differentiated liposarcoma of superficial soft tissue|8850/1
C0023827|T191|PT|0025508|CCPSS|LIPOSARCOMA|8850/3
C0023827|T191|PT|0000007477|CHV|liposarcoma|8850/3
C0023827|T191|SY|0000007477|CHV|liposarcomas|8850/3
C0023827|T191|PT|2000-7292|CSP|liposarcoma|8850/3
C0023827|T191|DI|U001066|DXP|LIPOSARCOMA|8850/3
C0023827|T191|PT|HP:0012034|HPO|Liposarcoma|8850/3
C0023827|T191|PT|sh88002663|LCH_NW|Liposarcoma|8850/3
C0023827|T191|LLT|10024627|MDR|Liposarcoma|8850/3
C0023827|T191|PT|10024627|MDR|Liposarcoma|8850/3
C0023827|T191|LLT|10024631|MDR|Liposarcoma NOS|8850/3
C0023827|T191|HT|10024628|MDR|Liposarcomas malignant|8850/3
C0023827|T191|PT|271512|MEDCIN|liposarcoma|8850/3
C0023827|T191|MH|D008080|MSH|Liposarcoma|8850/3
C0023827|T191|PM|D008080|MSH|Liposarcomas|8850/3
C0023827|T191|PN|NOCODE|MTH|liposarcoma|8850/3
C0023827|T191|PT|C3194|NCI|Liposarcoma|8850/3
C0023827|T191|SY|C3194|NCI|Liposarcoma Not Otherwise Specified|8850/3
C0023827|T191|PT|C3194|NCI_CDISC|LIPOSARCOMA, MALIGNANT|8850/3
C0023827|T191|PT|C3194|NCI_CPTAC|Liposarcoma|8850/3
C0023827|T191|PT|10024631|NCI_CTEP-SDC|Liposarcoma|8850/3
C0023827|T191|PT|C3194|NCI_CTRP|Liposarcoma|8850/3
C0023827|T191|DN|C3194|NCI_CTRP|Liposarcoma|8850/3
C0023827|T191|PT|CDR0000046028|NCI_NCI-GLOSS|liposarcoma|8850/3
C0023827|T191|SY|Xa99r|RCD|Fibroliposarcoma|8850/3
C0023827|T191|PT|X78Vj|RCD|Liposarcoma|8850/3
C0023827|T191|PT|Xa99r|RCD|Liposarcoma morphology|8850/3
C0023827|T191|OP|BBJ1.|RCDSY|Liposarcoma NOS|8850/3
C0023827|T191|SY|49430005|SNOMEDCT_US|Fibroliposarcoma|8850/3
C0023827|T191|PT|254829001|SNOMEDCT_US|Liposarcoma|8850/3
C0023827|T191|PT|49430005|SNOMEDCT_US|Liposarcoma|8850/3
C0023827|T191|SY|49430005|SNOMEDCT_US|Liposarcoma morphology|8850/3
C0023827|T191|SY|49430005|SNOMEDCT_US|Liposarcoma, no ICD-O subtype|8850/3
C0023827|T191|SY|49430005|SNOMEDCT_US|Liposarcoma, no International Classification of Diseases for Oncology subtype|8850/3
C0023827|T191|IS|49430005|SNOMEDCT_US|Liposarcoma, NOS|8850/3
C0334467|T191|PT|0000029990|CHV|fibrolipoma|8851/0
C0334467|T191|SY|273483|MEDCIN|adipose tissue fibrolipoma|8851/0
C0334467|T191|PT|273483|MEDCIN|fibrolipoma of fatty tissue|8851/0
C0334467|T191|PN|NOCODE|MTH|Fibrolipoma|8851/0
C0334467|T191|PT|C4249|NCI|Fibrolipoma|8851/0
C0334467|T191|PT|C4249|NCI_CDISC|FIBROLIPOMA, BENIGN|8851/0
C0334467|T191|PT|BBJ2.|RCD|Fibrolipoma|8851/0
C0334467|T191|PT|2710003|SNOMEDCT_US|Fibrolipoma|8851/0
C3274592|T191|SY|C99180|NCI|Infantile Fibromatosis, Non-Desmoid Type|8851/1
C3274592|T191|PT|C99180|NCI|Lipofibromatosis|8851/1
C3274592|T191|PT|703633001|SNOMEDCT_US|Lipofibromatosis|8851/1
C1370889|T191|PT|271513|MEDCIN|well differentiated liposarcoma|8851/3
C1370889|T191|ET|D008080|MSH|Atypical Lipomatous Tumor|8851/3
C1370889|T191|PM|D008080|MSH|Atypical Lipomatous Tumors|8851/3
C1370889|T191|PM|D008080|MSH|Lipomatous Tumor, Atypical|8851/3
C1370889|T191|ET|D008080|MSH|Liposarcoma, Well Differentiated|8851/3
C1370889|T191|PEP|D008080|MSH|Well Differentiated Liposarcoma|8851/3
C1370889|T191|PM|D008080|MSH|Well Differentiated Liposarcomas|8851/3
C1370889|T191|PN|NOCODE|MTH|Liposarcoma, well differentiated|8851/3
C1370889|T191|PT|C4250|NCI|Well Differentiated Liposarcoma|8851/3
C1370889|T191|SY|TCGA|NCI|Well Differentiated Liposarcoma|8851/3
C1370889|T191|SY|C4250|NCI|Well Differentiated Liposarcoma of Deep Soft Tissue|8851/3
C1370889|T191|SY|C4250|NCI|Well-Differentiated Liposarcoma|8851/3
C1370889|T191|SY|BBJ3.|RCD|Liposarcoma - differentiated|8851/3
C1370889|T191|AB|BBJ3.|RCD|Liposarcoma - well different|8851/3
C1370889|T191|PT|BBJ3.|RCD|Liposarcoma - well differentiated|8851/3
C1370889|T191|SY|28655007|SNOMEDCT_US|Liposarcoma - differentiated|8851/3
C1370889|T191|SY|28655007|SNOMEDCT_US|Liposarcoma - well differentiated|8851/3
C1370889|T191|SY|28655007|SNOMEDCT_US|Liposarcoma, differentiated|8851/3
C1370889|T191|PT|28655007|SNOMEDCT_US|Liposarcoma, well differentiated|8851/3
C0334470|T191|PT|MTHU028206|ICPC2ICD10ENG|fibromyxolipoma|8852/0
C0334470|T191|PT|MTHU051310|ICPC2ICD10ENG|myxolipoma|8852/0
C0334470|T191|SY|273491|MEDCIN|adipose tissue myxolipoma|8852/0
C0334470|T191|PT|273491|MEDCIN|myxolipoma of fatty tissue|8852/0
C0334470|T191|PT|C4251|NCI|Fibromyxolipoma|8852/0
C0334470|T191|SY|C4251|NCI|Myxolipoma|8852/0
C0334470|T191|PT|BBJ4.|RCD|Fibromyxolipoma|8852/0
C0334470|T191|SY|BBJ4.|RCD|Myxolipoma|8852/0
C0334470|T191|PT|58243007|SNOMEDCT_US|Fibromyxolipoma|8852/0
C0334470|T191|SY|58243007|SNOMEDCT_US|Myxolipoma|8852/0
C0206634|T191|SY|0000020983|CHV|liposarcoma myxoid|8852/3
C0206634|T191|PT|0000020983|CHV|myxoid liposarcoma|8852/3
C0206634|T191|SY|0000020983|CHV|myxoliposarcoma|8852/3
C0206634|T191|PT|HP:0012268|HPO|Myxoid liposarcoma|8852/3
C0206634|T191|PT|MTHU025479|ICPC2ICD10ENG|embryonal; liposarcoma|8852/3
C0206634|T191|PT|MTHU045619|ICPC2ICD10ENG|liposarcoma; embryonal|8852/3
C0545074|T191|PT|MTHU045621|ICPC2ICD10ENG|liposarcoma; mixed type|8852/3
C0206634|T191|PT|MTHU045623|ICPC2ICD10ENG|liposarcoma; myxoid|8852/3
C0334471|T191|PT|MTHU045625|ICPC2ICD10ENG|liposarcoma; round cell|8852/3
C0206634|T191|PT|MTHU051309|ICPC2ICD10ENG|myxoid; liposarcoma|8852/3
C0334471|T191|PT|MTHU065045|ICPC2ICD10ENG|round cell; liposarcoma|8852/3
C0206634|T191|LLT|10073137|MDR|Myxoid liposarcoma|8852/3
C0206634|T191|PT|10073137|MDR|Myxoid liposarcoma|8852/3
C0334471|T191|LLT|10073139|MDR|Round cell liposarcoma|8852/3
C0334471|T191|PT|10073139|MDR|Round cell liposarcoma|8852/3
C0545074|T191|PT|271517|MEDCIN|mixed type liposarcoma|8852/3
C0206634|T191|PT|271514|MEDCIN|myxoid liposarcoma|8852/3
C0334471|T191|PT|271515|MEDCIN|round cell liposarcoma|8852/3
C0206634|T191|MH|D018208|MSH|Liposarcoma, Myxoid|8852/3
C0206634|T191|PM|D018208|MSH|Liposarcoma, Round Cell|8852/3
C0206634|T191|PM|D018208|MSH|Liposarcomas, Myxoid|8852/3
C0206634|T191|ET|D018208|MSH|Myxoid Liposarcoma|8852/3
C0206634|T191|PM|D018208|MSH|Myxoid Liposarcomas|8852/3
C0206634|T191|ET|D018208|MSH|Round Cell Liposarcoma|8852/3
C0206634|T191|PM|D018208|MSH|Round Cell Liposarcomas|8852/3
C0206634|T191|PN|NOCODE|MTH|Liposarcoma, Myxoid|8852/3
C0545074|T191|PN|NOCODE|MTH|Myxoid/Round Cell Liposarcoma|8852/3
C0334471|T191|PN|NOCODE|MTH|Round Cell Liposarcoma|8852/3
C0334471|T191|OP|C4252|NCI|Cellular Myxoid Liposarcoma|8852/3
C0545074|T191|PT|C27781|NCI|Myxoid Liposarcoma|8852/3
C0545074|T191|SY|C27781|NCI|Myxoid/Round Cell Liposarcoma|8852/3
C0334471|T191|OP|C4252|NCI|Round Cell Liposarcoma|8852/3
C0334471|T191|PT|C4252|NCI|Round Cell Liposarcoma|8852/3
C0206634|T191|SY|CDR0000776766|PDQ|cellular myxoid liposarcoma|8852/3
C0545074|T191|PT|CDR0000776767|PDQ|myxoid liposarcoma|8852/3
C0545074|T191|SY|CDR0000776767|PDQ|myxoid/round cell liposarcoma|8852/3
C0334471|T191|PT|CDR0000776766|PDQ|round cell liposarcoma|8852/3
C0334471|T191|SY|BBJ6.|RCD|Lipoblastic liposarcoma|8852/3
C0206634|T191|PT|BBJ5.|RCD|Myxoid liposarcoma|8852/3
C0206634|T191|SY|BBJ5.|RCD|Myxoliposarcoma|8852/3
C0334471|T191|PT|BBJ6.|RCD|Round cell liposarcoma|8852/3
C0334471|T191|SY|404070007|SNOMEDCT_US|Lipoblastic liposarcoma|8852/3
C0334471|T191|SY|43296007|SNOMEDCT_US|Lipoblastic liposarcoma|8852/3
C0206634|T191|PT|404069006|SNOMEDCT_US|Myxoid liposarcoma|8852/3
C0206634|T191|PT|27849002|SNOMEDCT_US|Myxoid liposarcoma|8852/3
C0206634|T191|SY|27849002|SNOMEDCT_US|Myxoliposarcoma|8852/3
C0334471|T191|PT|43296007|SNOMEDCT_US|Round cell liposarcoma|8852/3
C0334471|T191|PT|404070007|SNOMEDCT_US|Round cell liposarcoma|8852/3
C0334471|T191|PT|MTHU045625|ICPC2ICD10ENG|liposarcoma; round cell|8853/3
C0334471|T191|PT|MTHU065045|ICPC2ICD10ENG|round cell; liposarcoma|8853/3
C0334471|T191|PT|10073139|MDR|Round cell liposarcoma|8853/3
C0334471|T191|LLT|10073139|MDR|Round cell liposarcoma|8853/3
C0334471|T191|PT|271515|MEDCIN|round cell liposarcoma|8853/3
C0334471|T191|PN|NOCODE|MTH|Round Cell Liposarcoma|8853/3
C0334471|T191|OP|C4252|NCI|Cellular Myxoid Liposarcoma|8853/3
C0334471|T191|OP|C4252|NCI|Round Cell Liposarcoma|8853/3
C0334471|T191|PT|C4252|NCI|Round Cell Liposarcoma|8853/3
C0334471|T191|PT|CDR0000776766|PDQ|round cell liposarcoma|8853/3
C0334471|T191|SY|BBJ6.|RCD|Lipoblastic liposarcoma|8853/3
C0334471|T191|PT|BBJ6.|RCD|Round cell liposarcoma|8853/3
C0334471|T191|SY|43296007|SNOMEDCT_US|Lipoblastic liposarcoma|8853/3
C0334471|T191|SY|404070007|SNOMEDCT_US|Lipoblastic liposarcoma|8853/3
C0334471|T191|PT|43296007|SNOMEDCT_US|Round cell liposarcoma|8853/3
C0334471|T191|PT|404070007|SNOMEDCT_US|Round cell liposarcoma|8853/3
C0205823|T191|SY|0000020723|CHV|lipoma pleomorphic|8854/0
C0205823|T191|PT|0000020723|CHV|pleomorphic lipoma|8854/0
C0205823|T191|PT|MTHU045604|ICPC2ICD10ENG|lipoma; pleomorphic|8854/0
C0205823|T191|PT|MTHU060028|ICPC2ICD10ENG|pleomorphic; lipoma|8854/0
C0205823|T191|ET|D008067|MSH|Atypical Lipoma|8854/0
C0205823|T191|PM|D008067|MSH|Atypical Lipomas|8854/0
C0205823|T191|PM|D008067|MSH|Lipoma, Atypical|8854/0
C0205823|T191|PEP|D008067|MSH|Lipoma, Pleomorphic|8854/0
C0205823|T191|PM|D008067|MSH|Lipomas, Atypical|8854/0
C0205823|T191|PM|D008067|MSH|Lipomas, Pleomorphic|8854/0
C0205823|T191|PM|D008067|MSH|Pleomorphic Lipoma|8854/0
C0205823|T191|PM|D008067|MSH|Pleomorphic Lipomas|8854/0
C0205823|T191|PN|NOCODE|MTH|Pleomorphic Lipoma|8854/0
C0205823|T191|PT|C3703|NCI|Pleomorphic Lipoma|8854/0
C0205823|T191|PT|X77od|RCD|Pleomorphic lipoma|8854/0
C0205823|T191|PT|404059000|SNOMEDCT_US|Pleomorphic lipoma|8854/0
C0205823|T191|PT|21396005|SNOMEDCT_US|Pleomorphic lipoma|8854/0
C0205823|T191|OAP|189783001|SNOMEDCT_US|Pleomorphic lipoma|8854/0
C0205823|T191|OF|189783001|SNOMEDCT_US|Pleomorphic lipoma|8854/0
C0205825|T191|PT|MTHU045624|ICPC2ICD10ENG|liposarcoma; pleomorphic|8854/3
C0205825|T191|PT|MTHU060029|ICPC2ICD10ENG|pleomorphic; liposarcoma|8854/3
C0205825|T191|PT|10073138|MDR|Pleomorphic liposarcoma|8854/3
C0205825|T191|LLT|10073138|MDR|Pleomorphic liposarcoma|8854/3
C0205825|T191|PT|271516|MEDCIN|pleomorphic liposarcoma|8854/3
C0205825|T191|PEP|D008080|MSH|Liposarcoma, Pleomorphic|8854/3
C0205825|T191|PM|D008080|MSH|Pleomorphic Liposarcoma|8854/3
C0205825|T191|PM|D008080|MSH|Pleomorphic Liposarcomas|8854/3
C0205825|T191|PT|C3705|NCI|Pleomorphic Liposarcoma|8854/3
C0205825|T191|PT|CDR0000776769|PDQ|pleomorphic liposarcoma|8854/3
C0205825|T191|PT|BBJ7.|RCD|Pleomorphic liposarcoma|8854/3
C0205825|T191|PT|404071006|SNOMEDCT_US|Pleomorphic liposarcoma|8854/3
C0205825|T191|PT|112683004|SNOMEDCT_US|Pleomorphic liposarcoma|8854/3
C0334472|T191|LLT|10073136|MDR|Mixed-type liposarcoma|8855/3
C0334472|T191|PT|10073136|MDR|Mixed-type liposarcoma|8855/3
C0334472|T191|PN|NOCODE|MTH|Mixed Liposarcoma|8855/3
C0334472|T191|PT|C4253|NCI|Mixed Liposarcoma|8855/3
C0334472|T191|PT|BBJ8.|RCD|Mixed liposarcoma|8855/3
C0334472|T191|PT|11073003|SNOMEDCT_US|Mixed liposarcoma|8855/3
C0334472|T191|SY|11073003|SNOMEDCT_US|Mixed-type liposarcoma|8855/3
C0334473|T191|SY|0000029991|CHV|infiltrating lipoma|8856/0
C0334473|T191|SY|0000029991|CHV|infiltrating lipomas|8856/0
C0334473|T191|PT|0000029991|CHV|intramuscular lipoma|8856/0
C0334473|T191|PT|MTHU039177|ICPC2ICD10ENG|infiltrating; lipoma|8856/0
C0334473|T191|PT|MTHU040073|ICPC2ICD10ENG|intramuscular; lipoma|8856/0
C0334473|T191|PT|MTHU045598|ICPC2ICD10ENG|lipoma; infiltrating|8856/0
C0334473|T191|PT|MTHU045600|ICPC2ICD10ENG|lipoma; intramuscular|8856/0
C0334473|T191|PT|C7451|NCI|Infiltrating Lipoma|8856/0
C0334473|T191|PT|C7450|NCI|Intramuscular Lipoma|8856/0
C0334473|T191|SY|BBJ9.|RCD|Infiltrating lipoma|8856/0
C0334473|T191|PT|BBJ9.|RCD|Intramuscular lipoma|8856/0
C0334473|T191|SY|24045002|SNOMEDCT_US|Infiltrating lipoma|8856/0
C0334473|T191|PT|24045002|SNOMEDCT_US|Intramuscular lipoma|8856/0
C0334474|T191|PT|MTHU045607|ICPC2ICD10ENG|lipoma; spindle cell|8857/0
C0334474|T191|PT|MTHU069006|ICPC2ICD10ENG|spindle cell; lipoma|8857/0
C0334474|T191|PT|C4254|NCI|Spindle Cell Lipoma|8857/0
C0334474|T191|PT|BBJA.|RCD|Spindle cell lipoma|8857/0
C0334474|T191|PT|404058008|SNOMEDCT_US|Spindle cell lipoma|8857/0
C0334474|T191|PT|27313007|SNOMEDCT_US|Spindle cell lipoma|8857/0
C1266130|T191|PT|271518|MEDCIN|fibroblastic liposarcoma|8857/3
C1266130|T191|PT|C6509|NCI|Fibroblastic Liposarcoma|8857/3
C1266130|T191|OP|C6509|NCI|Fibroblastic Liposarcoma|8857/3
C1266130|T191|PT|128883006|SNOMEDCT_US|Fibroblastic liposarcoma|8857/3
C0205824|T191|PT|MTHU030784|ICPC2ICD10ENG|dedifferentiated; liposarcoma|8858/3
C0205824|T191|PT|MTHU045620|ICPC2ICD10ENG|liposarcoma; dedifferentiated|8858/3
C0205824|T191|PT|10073135|MDR|Dedifferentiated liposarcoma|8858/3
C0205824|T191|LLT|10073135|MDR|Dedifferentiated liposarcoma|8858/3
C0205824|T191|PT|271519|MEDCIN|dedifferentiated liposarcoma|8858/3
C0205824|T191|PM|D008080|MSH|Dedifferentiated Liposarcoma|8858/3
C0205824|T191|PM|D008080|MSH|Dedifferentiated Liposarcomas|8858/3
C0205824|T191|PEP|D008080|MSH|Liposarcoma, Dedifferentiated|8858/3
C0205824|T191|SY|TCGA|NCI|Dedifferentiated Liposarcoma|8858/3
C0205824|T191|PT|C3704|NCI|Dedifferentiated Liposarcoma|8858/3
C0205824|T191|PT|CDR0000776768|PDQ|dedifferentiated liposarcoma|8858/3
C0205824|T191|PT|X77ob|RCD|Dedifferentiated liposarcoma|8858/3
C0205824|T191|AB|X77ob|RCDSY|Dedifferntiated liposarcoma|8858/3
C0205824|T191|OAP|189784007|SNOMEDCT_US|Dedifferentiated liposarcoma|8858/3
C0205824|T191|OF|189784007|SNOMEDCT_US|Dedifferentiated liposarcoma|8858/3
C0205824|T191|PT|67280001|SNOMEDCT_US|Dedifferentiated liposarcoma|8858/3
C0205824|T191|PT|404072004|SNOMEDCT_US|Dedifferentiated liposarcoma|8858/3
C0206633|T191|PT|0000020982|CHV|angiomyolipoma|8860/0
C0206633|T191|SY|0000020982|CHV|angiomyolipomas|8860/0
C0206633|T191|LLT|10051810|MDR|Angiomyolipoma|8860/0
C0206633|T191|PT|10051810|MDR|Angiomyolipoma|8860/0
C0206633|T191|MH|D018207|MSH|Angiomyolipoma|8860/0
C0206633|T191|PM|D018207|MSH|Angiomyolipomas|8860/0
C0206633|T191|PN|NOCODE|MTH|Angiomyolipoma|8860/0
C0206633|T191|PT|C3734|NCI|Angiomyolipoma|8860/0
C0206633|T191|DN|C3734|NCI_CTRP|Angiomyolipoma|8860/0
C0206633|T191|PT|CDR0000443027|NCI_NCI-GLOSS|angiomyolipoma|8860/0
C0206633|T191|PT|CDR0000441219|PDQ|angiomyolipoma|8860/0
C0206633|T191|PT|BBJB0|RCD|Angiomyolipoma|8860/0
C0206633|T191|PT|19929002|SNOMEDCT_US|Angiomyolipoma|8860/0
C2959647|T191|PT|447205003|SNOMEDCT_US|Angiomyomyelolipoma|8860/0
C0476076|T191|OP|BBJB1|RCDSY|Angiomyoliposarcoma|8860/3
C0476076|T191|PT|110457005|SNOMEDCT_US|Angiomyoliposarcoma|8860/3
C0206632|T191|PT|0000020981|CHV|angiolipoma|8861/0
C0206632|T191|SY|0000020981|CHV|angiolipomas|8861/0
C0206632|T191|PT|MTHU006368|ICPC2ICD10ENG|angiolipoma|8861/0
C0206632|T191|PT|10048945|MDR|Angiolipoma|8861/0
C0206632|T191|LLT|10048945|MDR|Angiolipoma|8861/0
C0206632|T191|SY|273479|MEDCIN|adipose tissue angiolipoma|8861/0
C0206632|T191|PT|273479|MEDCIN|angiolipoma of fatty tissue|8861/0
C0206632|T191|MH|D018206|MSH|Angiolipoma|8861/0
C0206632|T191|PM|D018206|MSH|Angiolipomas|8861/0
C0206632|T191|PT|C3733|NCI|Angiolipoma|8861/0
C0206632|T191|SY|C3733|NCI_CDISC|Angiolipoma|8861/0
C0206632|T191|PT|C3733|NCI_CDISC|ANGIOLIPOMA, BENIGN|8861/0
C0206632|T191|PT|Xa99s|RCD|Angiolipoma|8861/0
C0206632|T191|OP|BBJB2|RCDSY|Angiolipoma NOS|8861/0
C0206632|T191|PT|73219006|SNOMEDCT_US|Angiolipoma|8861/0
C0206632|T191|PT|404057003|SNOMEDCT_US|Angiolipoma|8861/0
C0206632|T191|IS|73219006|SNOMEDCT_US|Angiolipoma, NOS|8861/0
C1266131|T191|PT|C6503|NCI|Chondroid Lipoma|8862/0
C1266131|T191|PT|404065000|SNOMEDCT_US|Chondroid lipoma|8862/0
C1266131|T191|PT|128746001|SNOMEDCT_US|Chondroid lipoma|8862/0
C0206635|T191|PT|0000020984|CHV|myelolipoma|8870/0
C0206635|T191|SY|0000020984|CHV|myelolipomas|8870/0
C0206635|T191|PT|10077376|MDR|Myelolipoma|8870/0
C0206635|T191|LLT|10077376|MDR|Myelolipoma|8870/0
C0206635|T191|SY|273487|MEDCIN|adipose tissue myelolipoma|8870/0
C0206635|T191|PT|273487|MEDCIN|myelolipoma of fatty tissue|8870/0
C0206635|T191|MH|D018209|MSH|Myelolipoma|8870/0
C0206635|T191|PM|D018209|MSH|Myelolipomas|8870/0
C0206635|T191|PT|C3736|NCI|Adrenal Gland Myelolipoma|8870/0
C0206635|T191|SY|C3736|NCI|Myelolipoma|8870/0
C0206635|T191|SY|C3736|NCI_CDISC|Myelolipoma|8870/0
C0206635|T191|PT|C3736|NCI_CDISC|MYELOLIPOMA, BENIGN|8870/0
C0206635|T191|PT|BBJC.|RCD|Myelolipoma|8870/0
C0206635|T191|PT|20810002|SNOMEDCT_US|Myelolipoma|8870/0
C0205822|T191|PT|0000020722|CHV|hibernoma|8880/0
C0205822|T191|SY|0000020722|CHV|hibernomas|8880/0
C0205822|T191|PT|MTHU080728|ICPC2ICD10ENG|fat cells; fetal lipoma|8880/0
C0205822|T191|PT|MTHU080729|ICPC2ICD10ENG|fat cells; lipoma, fetal|8880/0
C0205822|T191|PT|MTHU029053|ICPC2ICD10ENG|fetal; lipoma, fat cells|8880/0
C0205822|T191|PT|MTHU045609|ICPC2ICD10ENG|lipoma; fat cells, fetal|8880/0
C0205822|T191|PT|MTHU045594|ICPC2ICD10ENG|lipoma; fetal, fat cells|8880/0
C0205822|T191|PEP|D008067|MSH|Hibernoma|8880/0
C0205822|T191|PM|D008067|MSH|Hibernomas|8880/0
C0205822|T191|PN|NOCODE|MTH|Hibernoma|8880/0
C0205822|T191|SY|C3702|NCI|Brown Fat Neoplasm|8880/0
C0205822|T191|SY|C3702|NCI|Brown Fat Tumor|8880/0
C0205822|T191|SY|C3702|NCI|Fetal Fat Cell Lipoma|8880/0
C0205822|T191|PT|C3702|NCI|Hibernoma|8880/0
C0205822|T191|SY|C3702|NCI_CDISC|Brown Fat Neoplasm|8880/0
C0205822|T191|SY|C3702|NCI_CDISC|Brown Fat Tumor|8880/0
C0205822|T191|SY|C3702|NCI_CDISC|Fetal Fat Cell Lipoma|8880/0
C0205822|T191|PT|C3702|NCI_CDISC|HIBERNOMA, BENIGN|8880/0
C0205822|T191|SY|BBJD.|RCD|Brown fat tumour|8880/0
C0205822|T191|SY|BBJD.|RCD|Fetal fat cell lipoma|8880/0
C0205822|T191|PT|BBJD.|RCD|Hibernoma|8880/0
C0205822|T191|SY|BBJD.|RCDAE|Brown fat tumor|8880/0
C0205822|T191|SY|77027006|SNOMEDCT_US|Brown fat tumor|8880/0
C0205822|T191|SYGB|77027006|SNOMEDCT_US|Brown fat tumour|8880/0
C0205822|T191|SY|77027006|SNOMEDCT_US|Fetal fat cell lipoma|8880/0
C0205822|T191|SYGB|77027006|SNOMEDCT_US|Foetal fat cell lipoma|8880/0
C0205822|T191|SY|404064001|SNOMEDCT_US|Granular cell lipoma|8880/0
C0205822|T191|PT|77027006|SNOMEDCT_US|Hibernoma|8880/0
C0205822|T191|PT|404064001|SNOMEDCT_US|Hibernoma|8880/0
C0334475|T191|LLT|10074548|MDR|Lipoblastomatosis|8881/0
C0334475|T191|PM|D062689|MSH|Lipoblastomatoses|8881/0
C0334475|T191|PEP|D062689|MSH|Lipoblastomatosis|8881/0
C0334475|T191|PN|NOCODE|MTH|Lipoblastomatosis|8881/0
C0334475|T191|SY|C4255|NCI|Fetal Lipomatosis|8881/0
C0334475|T191|PT|C4255|NCI|Lipoblastomatosis|8881/0
C0334475|T191|SY|XM1FN|RCD|Fetal lipomatosis|8881/0
C0334475|T191|PT|XM1FN|RCD|Lipoblastomatosis|8881/0
C0334475|T191|OP|BBJE.|RCDSY|Lipoblastomatosis|8881/0
C0334475|T191|OAS|274906009|SNOMEDCT_US|Fetal lipomatosis|8881/0
C0334475|T191|SY|63629005|SNOMEDCT_US|Fetal lipomatosis|8881/0
C0334475|T191|SY|400149007|SNOMEDCT_US|Fetal lipomatosis|8881/0
C0334475|T191|SY|63629005|SNOMEDCT_US|Foetal lipoma|8881/0
C0334475|T191|SY|63629005|SNOMEDCT_US|Foetal lipomatosis|8881/0
C0334475|T191|SY|400149007|SNOMEDCT_US|Foetal lipomatosis|8881/0
C0334475|T191|SY|63629005|SNOMEDCT_US|Lipoblastoma AND/OR lipoblastomatosis|8881/0
C1720179|T191|PT|420777000|SNOMEDCT_US|Lipoblastoma, circumscribed|8881/0
C1720128|T191|PT|421419001|SNOMEDCT_US|Lipoblastoma, diffuse|8881/0
C0334475|T191|PT|421098004|SNOMEDCT_US|Lipoblastoma/lipoblastomatosis|8881/0
C0334475|T191|PT|400149007|SNOMEDCT_US|Lipoblastomatosis|8881/0
C0334475|T191|PT|63629005|SNOMEDCT_US|Lipoblastomatosis|8881/0
C0334475|T191|OAP|274906009|SNOMEDCT_US|Lipoblastomatosis|8881/0
C0334475|T191|SY|421419001|SNOMEDCT_US|Lipoblastomatosis|8881/0
C0023267|T191|ET|0000004542|AOD|leiomyoma|8890/0
C0023267|T191|SY|BI00407|BI|fibroid|8890/0
C0042133|T191|SY|BI00407|BI|fibroid uterus|8890/0
C0042133|T191|PT|BI00407|BI|uterine fibroid|8890/0
C0023267|T191|PT|0037156|CCPSS|LEIOMYOMA|8890/0
C0042133|T191|PT|1017189|CCPSS|UTERINE LEIOMYOMA|8890/0
C0023267|T191|SY|0000007288|CHV|fibroid|8890/0
C0023267|T191|PT|0000007288|CHV|fibroid tumor|8890/0
C0023267|T191|SY|0000007288|CHV|fibroid tumors|8890/0
C0023267|T191|SY|0000007288|CHV|fibroids|8890/0
C0042133|T191|SY|0000012820|CHV|fibroids|8890/0
C0023267|T191|SY|0000007288|CHV|fibroids tumor|8890/0
C0023267|T191|SY|0000007288|CHV|fibroids tumors|8890/0
C0042133|T191|SY|0000012820|CHV|fibroleiomyoma|8890/0
C0042133|T191|SY|0000012820|CHV|fibromyoma|8890/0
C0023267|T191|SY|0000007288|CHV|fibromyoma|8890/0
C0023267|T191|SY|0000007288|CHV|fibromyomas|8890/0
C0023267|T191|SY|0000007288|CHV|leiomyofibroma|8890/0
C0042133|T191|SY|0000012820|CHV|leiomyofibroma|8890/0
C0042133|T191|SY|0000012820|CHV|leiomyoma|8890/0
C0023267|T191|SY|0000007288|CHV|leiomyoma|8890/0
C0042133|T191|SY|0000012820|CHV|leiomyoma of uterus|8890/0
C0042133|T191|SY|0000012820|CHV|leiomyomas|8890/0
C0023267|T191|SY|0000007288|CHV|leiomyomas|8890/0
C0042133|T191|SY|0000012820|CHV|myofibroma|8890/0
C0023267|T191|SY|0000007288|CHV|tumor fibroid|8890/0
C0042133|T191|PT|0000012820|CHV|tumor of uterine muscle|8890/0
C0042133|T191|SY|0000012820|CHV|uterine fibroid|8890/0
C0042133|T191|SY|0000012820|CHV|uterine fibroids|8890/0
C0042133|T191|SY|0000012820|CHV|uterine fibroma|8890/0
C0042133|T191|SY|0000012820|CHV|uterine fibromas|8890/0
C0042133|T191|SY|0000012820|CHV|uterine fibromyoma|8890/0
C0042133|T191|SY|0000012820|CHV|uterine leiomyoma|8890/0
C0042133|T191|SY|0000012820|CHV|uterine leiomyoma nos|8890/0
C0042133|T191|SY|0000012820|CHV|uterine myoma|8890/0
C0042133|T191|SY|0000012820|CHV|uterus fibroid|8890/0
C0042133|T191|SY|0000012820|CHV|uterus fibroids|8890/0
C0042133|T191|SY|0000012820|CHV|uterus fibroma|8890/0
C0042133|T191|SY|0000012820|CHV|uterus leiomyoma|8890/0
C0042133|T191|SY|0000012820|CHV|uterus myoma|8890/0
C0023267|T191|PT|NOCODE|COSTAR|Fibroids|8890/0
C0023267|T191|PT|449|COSTAR|LEIOMYOMA|8890/0
C0042133|T191|PT|NOCODE|COSTAR|Uterine Fibroid|8890/0
C0042133|T191|PT|769|COSTAR|UTERINE FIBROMA|8890/0
C0042133|T191|PT|NOCODE|COSTAR|Uterine Leiomyoma|8890/0
C0042133|T191|PT|NOCODE|COSTAR|Uterine Myoma|8890/0
C0023267|T191|SY|2011-3663|CSP|fibroid|8890/0
C0023267|T191|PT|2011-3663|CSP|leiomyoma|8890/0
C0042133|T191|GT|UTER FIBROID ENLARGE|CST|FIBROIDS|8890/0
C0042133|T191|GT|UTER FIBROID ENLARGE|CST|UTERINE FIBROID|8890/0
C0042133|T191|GT|UTER FIBROID ENLARGE|CST|UTERINE FIBROMYOMA|8890/0
C0042133|T191|SY|NOCODE|DXP|UTERUS, FIBROIDS|8890/0
C0042133|T191|SY|NOCODE|DXP|UTERUS, FIBROMYOMA|8890/0
C0042133|T191|DI|U001987|DXP|UTERUS, LEIOMYOMA|8890/0
C0042133|T191|SY|NOCODE|DXP|UTERUS, MYOMA|8890/0
C0042133|T191|SY|HP:0000131|HPO|Benign uterine leiomyomas|8890/0
C0042133|T191|SY|HP:0000131|HPO|Uterine fibroid|8890/0
C0042133|T191|PT|HP:0000131|HPO|Uterine leiomyoma|8890/0
C0042133|T191|HT|D25|ICD10|Leiomyoma of uterus|8890/0
C0042133|T191|PT|D25.9|ICD10|Leiomyoma of uterus, unspecified|8890/0
C0042133|T191|HT|D25|ICD10CM|Leiomyoma of uterus|8890/0
C0042133|T191|AB|D25|ICD10CM|Leiomyoma of uterus|8890/0
C0042133|T191|AB|D25.9|ICD10CM|Leiomyoma of uterus, unspecified|8890/0
C0042133|T191|PT|D25.9|ICD10CM|Leiomyoma of uterus, unspecified|8890/0
C0042133|T191|ET|D25|ICD10CM|uterine fibroid|8890/0
C0042133|T191|ET|D25|ICD10CM|uterine fibromyoma|8890/0
C0042133|T191|ET|D25|ICD10CM|uterine myoma|8890/0
C0042133|T191|PT|218.9|ICD9CM|Leiomyoma of uterus, unspecified|8890/0
C0042133|T191|HT|218|ICD9CM|Uterine leiomyoma|8890/0
C0042133|T191|AB|218.9|ICD9CM|Uterine leiomyoma NOS|8890/0
C0042133|T191|AB|X78|ICPC2EENG|Fibromyoma uterus|8890/0
C0042133|T191|PT|X78|ICPC2EENG|Fibromyoma uterus|8890/0
C0042133|T191|PT|MTHU028201|ICPC2ICD10ENG|fibromyoma; uterus|8890/0
C0042133|T191|PT|MTHU043162|ICPC2ICD10ENG|leiomyoma; uterus|8890/0
C0042133|T191|PT|MTHU078442|ICPC2ICD10ENG|uterus; fibromyoma|8890/0
C0042133|T191|PT|MTHU078496|ICPC2ICD10ENG|uterus; leiomyoma|8890/0
C0042133|T191|PT|X78001|ICPC2P|Fibroid;uterus|8890/0
C0042133|T191|PTN|X78005|ICPC2P|fibromyoma of the uterus|8890/0
C0042133|T191|PT|X78005|ICPC2P|Fibromyoma;uterus|8890/0
C0042133|T191|PT|X78002|ICPC2P|Myoma;uterus|8890/0
C0042133|T191|PTN|X78001|ICPC2P|uterine fibroid|8890/0
C0042133|T191|PTN|X78002|ICPC2P|uterine myoma|8890/0
C0042133|T191|PT|sh86005513|LCH_NW|Uterine fibroids|8890/0
C0023267|T191|LA|LA26513-4|LNC|Leiomyoma, NOS|8890/0
C0023267|T191|LLT|10016628|MDR|Fibroids|8890/0
C0023267|T191|PT|10024184|MDR|Leiomyoma|8890/0
C0023267|T191|LLT|10024184|MDR|Leiomyoma|8890/0
C0023267|T191|LLT|10024185|MDR|Leiomyoma NOS|8890/0
C0042133|T191|LLT|10024186|MDR|Leiomyoma of uterus, unspecified|8890/0
C0042133|T191|LLT|10046783|MDR|Uterine fibroid|8890/0
C0042133|T191|LLT|10046784|MDR|Uterine fibroids|8890/0
C0042133|T191|LLT|10081129|MDR|Uterine fibroma|8890/0
C0042133|T191|LLT|10046787|MDR|Uterine fibromyoma|8890/0
C0042133|T191|LLT|10046798|MDR|Uterine leiomyoma|8890/0
C0042133|T191|PT|10046798|MDR|Uterine leiomyoma|8890/0
C0042133|T191|LLT|10046801|MDR|Uterine myoma|8890/0
C0042133|T191|PT|31755|MEDCIN|benign leiomyoma of uterus|8890/0
C0042133|T191|ET|1222|MEDLINEPLUS|Fibroids|8890/0
C0042133|T191|SY|1222|MEDLINEPLUS|Fibroids|8890/0
C0042133|T191|PT|1222|MEDLINEPLUS|Uterine Fibroids|8890/0
C0042133|T191|ET|1222|MEDLINEPLUS|Uterine Leiomyomata|8890/0
C0042133|T191|SY|1222|MEDLINEPLUS|Uterine leiomyomata|8890/0
C0023267|T191|ET|D007889|MSH|Fibroid|8890/0
C0023267|T191|ET|D007889|MSH|Fibroid Tumor|8890/0
C0023267|T191|PM|D007889|MSH|Fibroid Tumors|8890/0
C0042133|T191|PEP|D007889|MSH|Fibroid Uterus|8890/0
C0042133|T191|PM|D007889|MSH|Fibroid, Uterine|8890/0
C0023267|T191|PM|D007889|MSH|Fibroids|8890/0
C0042133|T191|ET|D007889|MSH|Fibroids, Uterine|8890/0
C0042133|T191|ET|D007889|MSH|Fibroma, Uterine|8890/0
C0042133|T191|PM|D007889|MSH|Fibromas, Uterine|8890/0
C0023267|T191|ET|D007889|MSH|Fibromyoma|8890/0
C0023267|T191|PM|D007889|MSH|Fibromyomas|8890/0
C0023267|T191|MH|D007889|MSH|Leiomyoma|8890/0
C0042133|T191|ET|D007889|MSH|Leiomyoma, Uterine|8890/0
C0023267|T191|PM|D007889|MSH|Leiomyomas|8890/0
C0023267|T191|PM|D007889|MSH|Tumor, Fibroid|8890/0
C0023267|T191|PM|D007889|MSH|Tumors, Fibroid|8890/0
C0042133|T191|PM|D007889|MSH|Uterine Fibroid|8890/0
C0042133|T191|PM|D007889|MSH|Uterine Fibroids|8890/0
C0042133|T191|PM|D007889|MSH|Uterine Fibroma|8890/0
C0042133|T191|PM|D007889|MSH|Uterine Fibromas|8890/0
C0042133|T191|PM|D007889|MSH|Uterus, Fibroid|8890/0
C0023267|T191|PN|U002038|MTH|Fibroid Tumor|8890/0
C0042133|T191|PN|NOCODE|MTH|Uterine Fibroids|8890/0
C0042133|T191|PT|769|MTH|UTERUS FIBROMA|8890/0
C0042133|T191|SY|C3434|NCI|Body of Uterus Fibroid|8890/0
C0042133|T191|SY|C3434|NCI|Body of Uterus Leiomyoma|8890/0
C0042133|T191|SY|C3434|NCI|Corpus Uteri Fibroid|8890/0
C0042133|T191|SY|C3434|NCI|Corpus Uteri Leiomyoma|8890/0
C0023267|T191|SY|C3157|NCI|Fibroid|8890/0
C0042133|T191|SY|C3434|NCI|Fibroid of Body of Uterus|8890/0
C0042133|T191|SY|C3434|NCI|Fibroid of Corpus Uteri|8890/0
C0042133|T191|SY|C3434|NCI|Fibroid of the Body of Uterus|8890/0
C0042133|T191|SY|C3434|NCI|Fibroid of the Corpus Uteri|8890/0
C0042133|T191|SY|C3434|NCI|Fibroid of the Uterine Body|8890/0
C0042133|T191|SY|C3434|NCI|Fibroid of the Uterine Corpus|8890/0
C0042133|T191|SY|C3434|NCI|Fibroid of Uterine Body|8890/0
C0042133|T191|SY|C3434|NCI|Fibroid of Uterine Corpus|8890/0
C0023267|T191|PT|C3157|NCI|Leiomyoma|8890/0
C0042133|T191|SY|C3434|NCI|Leiomyoma of Body of Uterus|8890/0
C0042133|T191|SY|C3434|NCI|Leiomyoma of Corpus Uteri|8890/0
C0042133|T191|SY|C3434|NCI|Leiomyoma of the Body of Uterus|8890/0
C0042133|T191|SY|C3434|NCI|Leiomyoma of the Corpus Uteri|8890/0
C0042133|T191|SY|C3434|NCI|Leiomyoma of the Uterine Body|8890/0
C0042133|T191|SY|C3434|NCI|Leiomyoma of the Uterine Corpus|8890/0
C0042133|T191|SY|C3434|NCI|Leiomyoma of Uterine Body|8890/0
C0042133|T191|SY|C3434|NCI|Leiomyoma of Uterine Corpus|8890/0
C0023267|T191|SY|C3157|NCI|Leiomyomatous Tumor|8890/0
C0042133|T191|SY|C3434|NCI|Uterine Body Fibroid|8890/0
C0042133|T191|SY|C3434|NCI|Uterine Body Leiomyoma|8890/0
C0042133|T191|SY|C3434|NCI|Uterine Corpus Fibroid|8890/0
C0042133|T191|PT|C3434|NCI|Uterine Corpus Leiomyoma|8890/0
C0042133|T191|SY|C3434|NCI|Uterine Corpus Leiomyomata|8890/0
C0042133|T191|SY|C3434|NCI|Uterine Fibroid|8890/0
C0023267|T191|SY|C3157|NCI_CDISC|Fibroid|8890/0
C0023267|T191|SY|C3157|NCI_CDISC|Fibroid Neoplasm|8890/0
C0023267|T191|SY|C3157|NCI_CDISC|Fibroid Tumor|8890/0
C0023267|T191|PT|C3157|NCI_CDISC|LEIOMYOMA, BENIGN|8890/0
C0023267|T191|SY|C3157|NCI_CDISC|Leiomyomatous Neoplasm|8890/0
C0023267|T191|SY|C3157|NCI_CDISC|Leiomyomatous Tumor|8890/0
C0042133|T191|PT|C3434|NCI_CPTAC|Uterine Corpus Leiomyoma|8890/0
C0042133|T191|SY|C3434|NCI_CPTAC|Uterine Fibroids|8890/0
C0042133|T191|DN|C3434|NCI_CTRP|Uterine Corpus Leiomyoma|8890/0
C0023267|T191|PT|CDR0000046402|NCI_NCI-GLOSS|fibroid|8890/0
C0023267|T191|PT|CDR0000044870|NCI_NCI-GLOSS|leiomyoma|8890/0
C0042133|T191|OP|CDR0000279773|PDQ|uterine leiomyoma|8890/0
C0042133|T191|PT|CDR0000279978|PDQ|uterine leiomyomata|8890/0
C0042133|T191|SY|B78..|RCD|Fibroid uterus|8890/0
C0042133|T191|SY|B78..|RCD|Fibroids|8890/0
C0023267|T191|SY|Xa99u|RCD|Fibromyoma|8890/0
C0023267|T191|SY|Xa99u|RCD|Leiomyofibroma|8890/0
C0023267|T191|PT|Xa99u|RCD|Leiomyoma|8890/0
C0042133|T191|SY|B78..|RCD|Leiomyoma of body of uterus|8890/0
C0042133|T191|PT|B78..|RCD|Uterine fibroid|8890/0
C0042133|T191|SY|B78..|RCD|Uterine fibroids|8890/0
C0042133|T191|SY|B78..|RCD|Uterine leiomyoma - fibroids|8890/0
C0042133|T191|OP|B78z.|RCD|Uterine leiomyoma NOS|8890/0
C0023267|T191|OP|BBK00|RCDSY|Leiomyoma NOS|8890/0
C0023267|T191|OP|BBK0z|RCDSY|Leiomyomatous neoplasm NOS|8890/0
C0023267|T191|OP|BBK0.|RCDSY|Leiomyomatous neoplasms|8890/0
C4518207|T191|PT|733850003|SNOMEDCT_US|Apoplectic leiomyoma|8890/0
C1302861|T191|PT|400169002|SNOMEDCT_US|Benign leiomyomatous neoplasm - category|8890/0
C0042133|T191|SY|44598004|SNOMEDCT_US|Fibroid uterus|8890/0
C0042133|T191|SY|95315005|SNOMEDCT_US|Fibroid uterus|8890/0
C0042133|T191|SY|95315005|SNOMEDCT_US|Fibroids|8890/0
C0042133|T191|SY|44598004|SNOMEDCT_US|Fibroleiomyoma|8890/0
C0042133|T191|SY|44598004|SNOMEDCT_US|Fibromyoma|8890/0
C4518207|T191|SYGB|733850003|SNOMEDCT_US|Haemorrhagic cellular leiomyoma|8890/0
C4518207|T191|SY|733850003|SNOMEDCT_US|Hemorrhagic cellular leiomyoma|8890/0
C4542910|T191|PT|734305000|SNOMEDCT_US|Hydropic leiomyoma|8890/0
C0042133|T191|IS|44598004|SNOMEDCT_US|Leiomyofibroma|8890/0
C0023267|T191|PT|702978006|SNOMEDCT_US|Leiomyofibroma|8890/0
C0042133|T191|PT|146801000119103|SNOMEDCT_US|Leiomyoma|8890/0
C0042133|T191|PT|44598004|SNOMEDCT_US|Leiomyoma|8890/0
C0042133|T191|SY|95315005|SNOMEDCT_US|Leiomyoma of body of uterus|8890/0
C0042133|T191|SY|95315005|SNOMEDCT_US|Leiomyoma of uterus|8890/0
C0042133|T191|SY|44598004|SNOMEDCT_US|Leiomyoma, no ICD-O subtype|8890/0
C0042133|T191|SY|44598004|SNOMEDCT_US|Leiomyoma, no International Classification of Diseases for Oncology subtype|8890/0
C0042133|T191|IS|44598004|SNOMEDCT_US|Leiomyoma, NOS|8890/0
C4511806|T191|PT|726424006|SNOMEDCT_US|Mitotically active leiomyoma|8890/0
C0042133|T191|OAP|154616000|SNOMEDCT_US|Uterine fibroid|8890/0
C0042133|T191|OF|154616000|SNOMEDCT_US|Uterine fibroid|8890/0
C0042133|T191|SY|95315005|SNOMEDCT_US|Uterine fibroid|8890/0
C0042133|T191|SY|95315005|SNOMEDCT_US|Uterine fibroids|8890/0
C0042133|T191|SY|44598004|SNOMEDCT_US|Uterine fibroids|8890/0
C0042133|T191|PT|95315005|SNOMEDCT_US|Uterine leiomyoma|8890/0
C0042133|T191|SY|95315005|SNOMEDCT_US|Uterine leiomyoma - fibroids|8890/0
C0042133|T191|OAP|189106003|SNOMEDCT_US|Uterine leiomyoma NOS|8890/0
C0042133|T191|IS|95315005|SNOMEDCT_US|Uterine leiomyoma, NOS|8890/0
C0023267|T191|IT|0857|WHO|FIBROIDS|8890/0
C0042133|T191|PT|0857|WHO|UTERINE FIBROID|8890/0
C0042133|T191|IT|0857|WHO|UTERINE FIBROMYOMA|8890/0
C0206654|T191|PT|0050531|CCPSS|LEIOMYOMATOSIS|8890/1
C0206654|T191|PT|0000020998|CHV|leiomyomatosis|8890/1
C0206654|T191|PM|D018231|MSH|Leiomyomatoses|8890/1
C0206654|T191|MH|D018231|MSH|Leiomyomatosis|8890/1
C0206654|T191|PN|NOCODE|MTH|Leiomyomatosis|8890/1
C0267785|T191|SY|C3958|NCI|Diffuse Peritoneal Leiomyomatosis|8890/1
C0267785|T191|PT|C3958|NCI|Disseminated Peritoneal Leiomyomatosis|8890/1
C0206654|T191|PT|C3748|NCI|Leiomyomatosis|8890/1
C0267785|T191|SY|C3958|NCI|Leiomyomatosis Peritonealis Disseminata|8890/1
C0267785|T191|AB|Xa0Ej|RCD|Leiomyom perit disseminata|8890/1
C0206654|T191|PT|X77oh|RCD|Leiomyomatosis|8890/1
C0267785|T191|PT|Xa0Ej|RCD|Leiomyomatosis peritonealis disseminata|8890/1
C0206654|T191|OA|BBK01|RCDSY|Intravascul.leiomyomatosis|8890/1
C0206654|T191|OP|BBK01|RCDSY|Intravascular leiomyomatosis|8890/1
C0206654|T191|SY|75210008|SNOMEDCT_US|Intravascular leiomyomatosis|8890/1
C0206654|T191|SY|75210008|SNOMEDCT_US|Intravenous leiomyomatosis|8890/1
C0206654|T191|PT|75210008|SNOMEDCT_US|Leiomyomatosis|8890/1
C0267785|T191|PT|62557001|SNOMEDCT_US|Leiomyomatosis peritonealis disseminata|8890/1
C0206654|T191|SY|75210008|SNOMEDCT_US|Leiomyomatosis, no ICD-O subtype|8890/1
C0206654|T191|SY|75210008|SNOMEDCT_US|Leiomyomatosis, no International Classification of Diseases for Oncology subtype|8890/1
C0206654|T191|IS|75210008|SNOMEDCT_US|Leiomyomatosis, NOS|8890/1
C0267785|T191|PT|703634007|SNOMEDCT_US|Leiomyomatosis, peritonealis disseminata|8890/1
C0023269|T191|ET|0000004533|AOD|leiomyosarcoma|8890/3
C0023269|T191|PT|0047244|CCPSS|LEIOMYOSARCOMA|8890/3
C0023269|T191|PT|0000007289|CHV|leiomyosarcoma|8890/3
C0023269|T191|SY|0000007289|CHV|leiomyosarcomas|8890/3
C0023269|T191|PT|NOCODE|COSTAR|Leiomyosarcoma|8890/3
C0023269|T191|PT|2011-3842|CSP|leiomyosarcoma|8890/3
C0023269|T191|PT|HP:0100243|HPO|Leiomyosarcoma|8890/3
C0023269|T191|LA|LA26518-3|LNC|Leiomyosarcoma, NOS|8890/3
C0023269|T191|PT|10024189|MDR|Leiomyosarcoma|8890/3
C0023269|T191|LLT|10024189|MDR|Leiomyosarcoma|8890/3
C0023269|T191|LLT|10024193|MDR|Leiomyosarcoma NOS|8890/3
C0023269|T191|HT|10024190|MDR|Leiomyosarcomas|8890/3
C0023269|T191|PT|271521|MEDCIN|leiomyosarcoma|8890/3
C0023269|T191|MH|D007890|MSH|Leiomyosarcoma|8890/3
C0023269|T191|PM|D007890|MSH|Leiomyosarcomas|8890/3
C0023269|T191|PN|NOCODE|MTH|leiomyosarcoma|8890/3
C0023269|T191|PT|C3158|NCI|Leiomyosarcoma|8890/3
C0023269|T191|SY|TCGA|NCI|Leiomyosarcoma|8890/3
C0023269|T191|PT|C3158|NCI_CDISC|LEIOMYOSARCOMA, MALIGNANT|8890/3
C0023269|T191|SY|C3158|NCI_CDISC|Leiomyosarcomas|8890/3
C0023269|T191|PT|C3158|NCI_CPTAC|Leiomyosarcoma|8890/3
C0023269|T191|SY|10024193|NCI_CTEP-SDC|Leiomyosarcoma - not uterine|8890/3
C0023269|T191|PT|C3158|NCI_CTRP|Leiomyosarcoma|8890/3
C0023269|T191|DN|C3158|NCI_CTRP|Leiomyosarcoma|8890/3
C0023269|T191|PT|CDR0000046027|NCI_NCI-GLOSS|leiomyosarcoma|8890/3
C0023269|T191|PT|Xa99v|RCD|Leiomyosarcoma|8890/3
C0023269|T191|SY|Xa99v|RCD|LMS - Leiomyosarcoma|8890/3
C0023269|T191|OP|BBK02|RCDSY|Leiomyosarcoma NOS|8890/3
C0023269|T191|PT|51549004|SNOMEDCT_US|Leiomyosarcoma|8890/3
C0023269|T191|PT|443719001|SNOMEDCT_US|Leiomyosarcoma|8890/3
C0023269|T191|SY|51549004|SNOMEDCT_US|Leiomyosarcoma, no subtype|8890/3
C0023269|T191|IS|51549004|SNOMEDCT_US|Leiomyosarcoma, NOS|8890/3
C0023269|T191|SY|51549004|SNOMEDCT_US|LMS - Leiomyosarcoma|8890/3
C0086533|T191|LLT|10051431|MDR|Epithelioid leiomyoma|8891/0
C0086533|T191|LLT|10067401|MDR|Leiomyoblastoma|8891/0
C0086533|T191|PM|D018230|MSH|Epithelioid Leiomyoma|8891/0
C0086533|T191|PM|D018230|MSH|Epithelioid Leiomyomas|8891/0
C0086533|T191|ET|D018230|MSH|Leiomyoblastoma|8891/0
C0086533|T191|PM|D018230|MSH|Leiomyoblastomas|8891/0
C0086533|T191|MH|D018230|MSH|Leiomyoma, Epithelioid|8891/0
C0086533|T191|PM|D018230|MSH|Leiomyomas, Epithelioid|8891/0
C0086533|T191|PT|C3486|NCI|Epithelioid Cell Type Gastrointestinal Stromal Tumor|8891/0
C0086533|T191|SY|C3486|NCI|Epithelioid Cell Type GIST|8891/0
C0086533|T191|OP|C3486|NCI|Leiomyoblastoma|8891/0
C0086533|T191|OP|C3486|NCI|Stout's Leiomyoblastoma|8891/0
C0086533|T191|PT|BBK03|RCD|Epithelioid leiomyoma|8891/0
C0086533|T191|SY|BBK03|RCD|Leiomyoblastoma|8891/0
C0086533|T191|PT|19071004|SNOMEDCT_US|Epithelioid leiomyoma|8891/0
C0086533|T191|SY|19071004|SNOMEDCT_US|Leiomyoblastoma|8891/0
C0205815|T191|PT|271522|MEDCIN|epithelioid leiomyosarcoma|8891/3
C0205815|T191|PM|D007890|MSH|Epithelioid Leiomyosarcoma|8891/3
C0205815|T191|PM|D007890|MSH|Epithelioid Leiomyosarcomas|8891/3
C0205815|T191|PEP|D007890|MSH|Leiomyosarcoma, Epithelioid|8891/3
C0205815|T191|PM|D007890|MSH|Leiomyosarcomas, Epithelioid|8891/3
C0205815|T191|PT|C3700|NCI|Epithelioid Leiomyosarcoma|8891/3
C0205815|T191|PT|BBK04|RCD|Epithelioid leiomyosarcoma|8891/3
C0205815|T191|PT|42392001|SNOMEDCT_US|Epithelioid leiomyosarcoma|8891/3
C0334477|T191|PT|C4256|NCI|Cellular Leiomyoma|8892/0
C0334477|T191|PT|BBK05|RCD|Cellular leiomyoma|8892/0
C0334477|T191|PT|90955001|SNOMEDCT_US|Cellular leiomyoma|8892/0
C0334478|T191|SY|0000029992|CHV|atypical leiomyoma|8893/0
C0334478|T191|SY|0000029992|CHV|bizarre leiomyoma|8893/0
C0334478|T191|PT|0000029992|CHV|symplastic leiomyoma|8893/0
C0334478|T191|SY|C4257|NCI|Atypical Leiomyoma|8893/0
C0334478|T191|PT|C4257|NCI|Bizarre Leiomyoma|8893/0
C0334478|T191|SY|C4257|NCI|Pleomorphic Leiomyoma|8893/0
C0334478|T191|PT|BBK06|RCD|Bizarre leiomyoma|8893/0
C0334478|T191|SY|48897006|SNOMEDCT_US|Atypical leiomyoma|8893/0
C0334478|T191|PT|48897006|SNOMEDCT_US|Bizarre leiomyoma|8893/0
C0334478|T191|SY|48897006|SNOMEDCT_US|Pleomorphic leiomyoma|8893/0
C0334478|T191|IS|48897006|SNOMEDCT_US|Symplastic leiomyoma|8893/0
C0334478|T191|SY|48897006|SNOMEDCT_US|Symplastic leiomyoma|8893/0
C0206653|T191|PT|0000020997|CHV|angioleiomyoma|8894/0
C0206653|T191|SY|0000020997|CHV|angiomyoma|8894/0
C0206653|T191|LLT|10068762|MDR|Angioleiomyoma|8894/0
C0206653|T191|ET|D018229|MSH|Angioleiomyoma|8894/0
C0206653|T191|PM|D018229|MSH|Angioleiomyomas|8894/0
C0206653|T191|MH|D018229|MSH|Angiomyoma|8894/0
C0206653|T191|PM|D018229|MSH|Angiomyomas|8894/0
C0206653|T191|ET|D018229|MSH|Leiomyoma, Vascular|8894/0
C0206653|T191|PM|D018229|MSH|Leiomyomas, Vascular|8894/0
C0206653|T191|PM|D018229|MSH|Vascular Leiomyoma|8894/0
C0206653|T191|PM|D018229|MSH|Vascular Leiomyomas|8894/0
C0206653|T191|PT|C3747|NCI|Angioleiomyoma|8894/0
C0206653|T191|SY|C3747|NCI|Angiomyoma|8894/0
C0206653|T191|SY|C3747|NCI|Vascular Leiomyoma|8894/0
C0206653|T191|SY|BBK10|RCD|Angioleiomyoma|8894/0
C0206653|T191|PT|BBK10|RCD|Angiomyoma|8894/0
C0206653|T191|SY|BBK10|RCD|Vascular leiomyoma|8894/0
C0206653|T191|SY|86959002|SNOMEDCT_US|Angioleiomyoma|8894/0
C0206653|T191|PT|86959002|SNOMEDCT_US|Angiomyoma|8894/0
C0206653|T191|SY|86959002|SNOMEDCT_US|Vascular leiomyoma|8894/0
C0334479|T191|PT|271529|MEDCIN|angiomyosarcoma|8894/3
C0334479|T191|OP|C66771|NCI|Angiomyosarcoma|8894/3
C0334479|T191|PT|C66771|NCI|Angiomyosarcoma|8894/3
C0334479|T191|PT|BBK11|RCD|Angiomyosarcoma|8894/3
C0334479|T191|PT|28953002|SNOMEDCT_US|Angiomyosarcoma|8894/3
C0027086|T191|ET|0000004540|AOD|myoma|8895/0
C0027086|T191|PT|0000008435|CHV|myoma|8895/0
C0027086|T191|SY|0000008435|CHV|myomas|8895/0
C0027086|T191|PT|NOCODE|COSTAR|Myoma|8895/0
C0027086|T191|ET|2011-3484|CSP|myoma|8895/0
C0027086|T191|PT|HP:0031460|HPO|Benign muscle neoplasm|8895/0
C0027086|T191|ET|D21|ICD10CM|benign neoplasm of muscle|8895/0
C0027086|T191|LLT|10061692|MDR|Benign muscle neoplasm|8895/0
C0027086|T191|PT|10061692|MDR|Benign muscle neoplasm|8895/0
C0027086|T191|LLT|10048613|MDR|Benign muscle neoplasm NOS|8895/0
C0027086|T191|LLT|10074632|MDR|Myoma|8895/0
C0027086|T191|MH|D009214|MSH|Myoma|8895/0
C0027086|T191|PM|D009214|MSH|Myomas|8895/0
C0027086|T191|PT|C4882|NCI|Benign Muscle Neoplasm|8895/0
C0027086|T191|SY|C4882|NCI|Benign Muscle Tumor|8895/0
C0027086|T191|SY|C4882|NCI|Benign Neoplasm of Muscle|8895/0
C0027086|T191|SY|C4882|NCI|Benign Neoplasm of the Muscle|8895/0
C0027086|T191|SY|C4882|NCI|Benign Tumor of Muscle|8895/0
C0027086|T191|SY|C4882|NCI|Benign Tumor of the Muscle|8895/0
C0027086|T191|SY|C4882|NCI|Myoma|8895/0
C0027086|T191|PT|X78Vn|RCD|Benign tumour of muscle|8895/0
C0027086|T191|PT|BBK20|RCD|Myoma|8895/0
C0027086|T191|PT|X78Vn|RCDAE|Benign tumor of muscle|8895/0
C0027086|T191|PT|92237006|SNOMEDCT_US|Benign neoplasm of muscle|8895/0
C0027086|T191|IS|92237006|SNOMEDCT_US|Benign neoplasm of muscle, NOS|8895/0
C0027086|T191|SY|92237006|SNOMEDCT_US|Benign tumor of muscle|8895/0
C0027086|T191|SYGB|92237006|SNOMEDCT_US|Benign tumour of muscle|8895/0
C0027086|T191|PT|66357004|SNOMEDCT_US|Myoma|8895/0
C0027086|T191|SY|66357004|SNOMEDCT_US|Myoma, no ICD-O subtype|8895/0
C0027086|T191|SY|66357004|SNOMEDCT_US|Myoma, no International Classification of Diseases for Oncology subtype|8895/0
C0684743|T191|SY|0000044007|CHV|cancer muscle|8895/3
C0684743|T191|SY|0000044007|CHV|cancer muscles|8895/3
C0684743|T191|SY|0000044007|CHV|cancer of muscle|8895/3
C0684743|T191|SY|0000044007|CHV|cancer of the muscle|8895/3
C0684743|T191|PT|0000044007|CHV|muscle cancer|8895/3
C0684743|T191|SY|0000044007|CHV|muscle cancers|8895/3
C0027095|T191|PT|0000008439|CHV|myosarcoma|8895/3
C0684743|T191|ET|C49|ICD10CM|malignant neoplasm of muscle|8895/3
C0684743|T191|PTN|L71015|ICPC2P|malignant neosplasm of the muscles|8895/3
C0684743|T191|PT|sh2010009786|LCH_NW|Muscles--Cancer|8895/3
C0684743|T191|LA|LA10546-2|LNC|Muscle Cancer|8895/3
C0684743|T191|LLT|10062050|MDR|Malignant muscle neoplasm|8895/3
C0684743|T191|PT|10062050|MDR|Malignant muscle neoplasm|8895/3
C0684743|T191|LLT|10050530|MDR|Malignant muscle neoplasm NOS|8895/3
C0684743|T191|PT|352781|MEDCIN|malignant neoplasm of muscle|8895/3
C0027095|T191|PT|271520|MEDCIN|myosarcoma|8895/3
C0684743|T191|PEP|D019042|MSH|Cancer of Muscle|8895/3
C0684743|T191|ET|D019042|MSH|Cancer of the Muscle|8895/3
C0684743|T191|PM|D019042|MSH|Cancer, Muscle|8895/3
C0684743|T191|PM|D019042|MSH|Cancers, Muscle|8895/3
C0684743|T191|ET|D019042|MSH|Muscle Cancer|8895/3
C0684743|T191|PM|D019042|MSH|Muscle Cancers|8895/3
C0027095|T191|MH|D009217|MSH|Myosarcoma|8895/3
C0027095|T191|PM|D009217|MSH|Myosarcomas|8895/3
C0684743|T191|PN|NOCODE|MTH|Malignant neoplasm of muscle|8895/3
C0027095|T191|PN|NOCODE|MTH|Myosarcoma|8895/3
C0684743|T191|PT|C4883|NCI|Malignant Muscle Neoplasm|8895/3
C0684743|T191|SY|C4883|NCI|Malignant Muscle Tumor|8895/3
C0684743|T191|SY|C4883|NCI|Malignant Neoplasm of Muscle|8895/3
C0684743|T191|SY|C4883|NCI|Malignant Neoplasm of the Muscle|8895/3
C0684743|T191|SY|C4883|NCI|Malignant Tumor of Muscle|8895/3
C0684743|T191|SY|C4883|NCI|Malignant Tumor of the Muscle|8895/3
C0684743|T191|SY|C4883|NCI|Myosarcoma|8895/3
C0684743|T191|PT|C4883|NCI_CPTAC|Malignant Muscle Neoplasm|8895/3
C0684743|T191|DN|C4883|NCI_CTRP|Malignant Muscle Neoplasm|8895/3
C0684743|T191|SY|CDR0000039804|PDQ|malignant muscle neoplasm|8895/3
C0684743|T191|SY|CDR0000039804|PDQ|malignant muscle tumor|8895/3
C0684743|T191|SY|CDR0000039804|PDQ|malignant neoplasm of muscle|8895/3
C0684743|T191|SY|CDR0000039804|PDQ|malignant neoplasm of the muscle|8895/3
C0684743|T191|SY|CDR0000039804|PDQ|malignant tumor of muscle|8895/3
C0684743|T191|SY|CDR0000039804|PDQ|malignant tumor of the muscle|8895/3
C0684743|T191|PT|CDR0000039804|PDQ|muscle cancer|8895/3
C0684743|T191|SY|CDR0000039804|PDQ|myosarcoma|8895/3
C0684743|T191|SY|X78Vm|RCD|CA - Cancer of muscle|8895/3
C0684743|T191|SY|X78Vm|RCD|Cancer of muscle|8895/3
C0684743|T191|PT|X78Vm|RCD|Malignant tumour of muscle|8895/3
C0027095|T191|PT|BBK21|RCD|Myosarcoma|8895/3
C0684743|T191|PT|X78Vm|RCDAE|Malignant tumor of muscle|8895/3
C0684743|T191|SY|363495004|SNOMEDCT_US|CA - Cancer of muscle|8895/3
C0684743|T191|SY|363495004|SNOMEDCT_US|Cancer of muscle|8895/3
C0684743|T191|IS|93913006|SNOMEDCT_US|Malignant neoplasm of muscle|8895/3
C0684743|T191|IS|93913006|SNOMEDCT_US|Malignant neoplasm of muscle, NOS|8895/3
C0684743|T191|PT|363495004|SNOMEDCT_US|Malignant tumor of muscle|8895/3
C0684743|T191|PTGB|363495004|SNOMEDCT_US|Malignant tumour of muscle|8895/3
C0027095|T191|PT|20667008|SNOMEDCT_US|Myosarcoma|8895/3
C2347314|T191|PT|C67563|NCI|Myxoid Leiomyoma|8896/0
C2347314|T191|PT|703635008|SNOMEDCT_US|Myxoid leiomyoma|8896/0
C0205816|T191|PT|271523|MEDCIN|myxoid leiomyosarcoma|8896/3
C0205816|T191|PEP|D007890|MSH|Leiomyosarcoma, Myxoid|8896/3
C0205816|T191|PM|D007890|MSH|Leiomyosarcomas, Myxoid|8896/3
C0205816|T191|PM|D007890|MSH|Myxoid Leiomyosarcoma|8896/3
C0205816|T191|PM|D007890|MSH|Myxoid Leiomyosarcomas|8896/3
C0205816|T191|PT|C3701|NCI|Myxoid Leiomyosarcoma|8896/3
C0205816|T191|PT|X77of|RCD|Myxoid leiomyosarcoma|8896/3
C0205816|T191|OAP|189792003|SNOMEDCT_US|Myxoid leiomyosarcoma|8896/3
C0205816|T191|OF|189792003|SNOMEDCT_US|Myxoid leiomyosarcoma|8896/3
C0205816|T191|PT|16090008|SNOMEDCT_US|Myxoid leiomyosarcoma|8896/3
C0206658|T191|SY|0000021001|CHV|muscle smooth tumor|8897/1
C0206658|T191|PT|0000021001|CHV|smooth muscle tumor|8897/1
C0206658|T191|SY|0000021001|CHV|smooth muscle tumors|8897/1
C0206658|T191|PT|sh86005515|LCH_NW|Smooth muscle--Tumors|8897/1
C0206658|T191|PM|D018235|MSH|Muscle Tumor, Smooth|8897/1
C0206658|T191|PM|D018235|MSH|Muscle Tumors, Smooth|8897/1
C0206658|T191|MH|D018235|MSH|Smooth Muscle Tumor|8897/1
C0206658|T191|PM|D018235|MSH|Smooth Muscle Tumors|8897/1
C0206658|T191|PM|D018235|MSH|Tumor, Smooth Muscle|8897/1
C0206658|T191|PM|D018235|MSH|Tumors, Smooth Muscle|8897/1
C1519864|T191|SY|C40177|NCI|Borderline Uterine Corpus Smooth Muscle Neoplasm|8897/1
C0206658|T191|SY|C3751|NCI|Neoplasm of Smooth Muscle|8897/1
C0206658|T191|SY|C3751|NCI|Neoplasm of the Smooth Muscle|8897/1
C0206658|T191|PT|C3751|NCI|Smooth Muscle Neoplasm|8897/1
C0206658|T191|SY|C3751|NCI|Smooth Muscle Tumor|8897/1
C0206658|T191|SY|C3751|NCI|Tumor of Smooth Muscle|8897/1
C0206658|T191|SY|C3751|NCI|Tumor of the Smooth Muscle|8897/1
C1519864|T191|SY|C40177|NCI|Uterine Corpus Smooth Muscle Neoplasm of Uncertain Malignant Potential|8897/1
C1519864|T191|PT|C40177|NCI|Uterine Corpus Smooth Muscle Tumor of Uncertain Malignant Potential|8897/1
C1519864|T191|AB|C40177|NCI|Uterine Corpus STUMP|8897/1
C0206658|T191|PT|X77oi|RCD|Smooth muscle tumour|8897/1
C0206658|T191|PT|X77oi|RCDAE|Smooth muscle tumor|8897/1
C0206658|T191|OP|BBK38|RCDSA|Smooth muscle tumor NOS|8897/1
C0206658|T191|OP|BBK38|RCDSY|Smooth muscle tumour NOS|8897/1
C0206658|T191|PT|75109009|SNOMEDCT_US|Smooth muscle tumor|8897/1
C0206658|T191|SY|75109009|SNOMEDCT_US|Smooth muscle tumor of uncertain malignant potential|8897/1
C0206658|T191|IS|75109009|SNOMEDCT_US|Smooth muscle tumor, NOS|8897/1
C0206658|T191|PTGB|75109009|SNOMEDCT_US|Smooth muscle tumour|8897/1
C0206658|T191|SYGB|75109009|SNOMEDCT_US|Smooth muscle tumour of uncertain malignant potential|8897/1
C1266132|T191|SY|0000056690|CHV|metastasising leiomyoma|8898/1
C1266132|T191|PT|0000056690|CHV|metastasizing leiomyoma|8898/1
C1511090|T191|PT|C40173|NCI|Benign Metastasizing Leiomyoma of the Uterine Corpus|8898/1
C1511090|T191|SY|C40173|NCI|Uterine Corpus Metastasizing Leiomyoma|8898/1
C1266132|T191|PTGB|128747005|SNOMEDCT_US|Metastasising leiomyoma|8898/1
C1266132|T191|PT|128747005|SNOMEDCT_US|Metastasizing leiomyoma|8898/1
C0035411|T191|ET|0000004541|AOD|rhabdomyoma|8900/0
C0035411|T191|PT|0000010836|CHV|rhabdomyoma|8900/0
C0035411|T191|SY|0000010836|CHV|rhabdomyomas|8900/0
C0035411|T191|PT|HP:0009730|HPO|Rhabdomyoma|8900/0
C0035411|T191|LLT|10028633|MDR|Myoma striocellulare|8900/0
C0035411|T191|LLT|10039021|MDR|Rhabdomyoma|8900/0
C0035411|T191|PT|10039021|MDR|Rhabdomyoma|8900/0
C0035411|T191|MH|D012207|MSH|Rhabdomyoma|8900/0
C0035411|T191|PM|D012207|MSH|Rhabdomyomas|8900/0
C0035411|T191|PN|NOCODE|MTH|Rhabdomyoma|8900/0
C0035411|T191|PT|C3358|NCI|Rhabdomyoma|8900/0
C0035411|T191|PT|C3358|NCI_CDISC|RHABDOMYOMA, BENIGN|8900/0
C0035411|T191|PT|C3358|NCI_NICHD|Rhabdomyoma|8900/0
C0035411|T191|SY|C3358|NCI_NICHD|Rhabdomyomatous Neoplasm|8900/0
C0035411|T191|PT|Xa99x|RCD|Rhabdomyoma|8900/0
C0035411|T191|PT|BBK30|RCDSY|Rhabdomyoma NOS|8900/0
C0035411|T191|OA|BBK3z|RCDSY|Rhabdomyomatous neopl.NOS|8900/0
C0035411|T191|OP|BBK3z|RCDSY|Rhabdomyomatous neoplasm NOS|8900/0
C0035411|T191|OP|BBK3.|RCDSY|Rhabdomyomatous neoplasms|8900/0
C0035411|T191|PT|302846007|SNOMEDCT_US|Rhabdomyoma|8900/0
C0035411|T191|PT|43375002|SNOMEDCT_US|Rhabdomyoma|8900/0
C0035411|T191|SY|43375002|SNOMEDCT_US|Rhabdomyoma, no ICD-O subtype|8900/0
C0035411|T191|SY|43375002|SNOMEDCT_US|Rhabdomyoma, no International Classification of Diseases for Oncology subtype|8900/0
C0035411|T191|IS|43375002|SNOMEDCT_US|Rhabdomyoma, NOS|8900/0
C0035411|T191|PT|402877008|SNOMEDCT_US|Rhabdomyomatous neoplasm|8900/0
C0035412|T191|ET|0000004534|AOD|rhabdomyosarcoma|8900/3
C0035412|T191|PT|0041857|CCPSS|RHABDOMYOSARCOMA|8900/3
C0035412|T191|PT|0000010837|CHV|rhabdomyosarcoma|8900/3
C0035412|T191|SY|0000010837|CHV|rhabdomyosarcomas|8900/3
C0035412|T191|SY|0000010837|CHV|rhabdosarcoma|8900/3
C0035412|T191|PT|NOCODE|COSTAR|Rhabdomyosarcoma|8900/3
C0035412|T191|ET|2011-4200|CSP|rhabdomyoblastoma|8900/3
C0035412|T191|PT|2011-4200|CSP|rhabdomyosarcoma|8900/3
C0035412|T191|ET|2011-4200|CSP|rhabdosarcoma|8900/3
C0035412|T191|DI|U001679|DXP|RHABDOMYOSARCOMA|8900/3
C0035412|T191|PT|HP:0002859|HPO|Rhabdomyosarcoma|8900/3
C0035412|T191|PT|U004115|LCH|Rhabdomyosarcoma|8900/3
C0035412|T191|PT|sh85113568|LCH_NW|Rhabdomyosarcoma|8900/3
C0035412|T191|LLT|10039022|MDR|Rhabdomyosarcoma|8900/3
C0035412|T191|PT|10039022|MDR|Rhabdomyosarcoma|8900/3
C0035412|T191|LLT|10039024|MDR|Rhabdomyosarcoma NOS|8900/3
C0035412|T191|HT|10039023|MDR|Rhabdomyosarcomas|8900/3
C0035412|T191|LLT|10039028|MDR|Rhabdosarcoma|8900/3
C0035412|T191|SY|31683|MEDCIN|malignant neoplasm myosarcoma rhabdomyosarcoma|8900/3
C0035412|T191|PT|31683|MEDCIN|rhabdomyosarcoma|8900/3
C0035412|T191|ET|495|MEDLINEPLUS|Rhabdomyosarcoma|8900/3
C0035412|T191|MH|D012208|MSH|Rhabdomyosarcoma|8900/3
C0035412|T191|PM|D012208|MSH|Rhabdomyosarcomas|8900/3
C0035412|T191|PN|NOCODE|MTH|Rhabdomyosarcoma|8900/3
C0035412|T191|PT|C3359|NCI|Rhabdomyosarcoma|8900/3
C0035412|T191|PT|C3359|NCI_CDISC|RHABDOMYOSARCOMA, MALIGNANT|8900/3
C0035412|T191|PT|C3359|NCI_CPTAC|Rhabdomyosarcoma|8900/3
C0035412|T191|PT|10039024|NCI_CTEP-SDC|Rhabdomyosarcoma, NOS|8900/3
C0035412|T191|PT|CDR0000045872|NCI_NCI-GLOSS|rhabdomyosarcoma|8900/3
C0035412|T191|PT|C3359|NCI_NICHD|Rhabdomyosarcoma|8900/3
C0035412|T191|PT|Xa99y|RCD|Rhabdomyosarcoma|8900/3
C0035412|T191|SY|Xa99y|RCD|Rhabdosarcoma|8900/3
C0035412|T191|PT|BBK31|RCDSY|Rhabdomyosarcoma NOS|8900/3
C0035412|T191|PT|302847003|SNOMEDCT_US|Rhabdomyosarcoma|8900/3
C0035412|T191|PT|30924005|SNOMEDCT_US|Rhabdomyosarcoma|8900/3
C0035412|T191|SY|30924005|SNOMEDCT_US|Rhabdomyosarcoma, no subtype|8900/3
C0035412|T191|IS|30924005|SNOMEDCT_US|Rhabdomyosarcoma, NOS|8900/3
C0035412|T191|SY|30924005|SNOMEDCT_US|Rhabdosarcoma|8900/3
C0035412|T191|SY|302847003|SNOMEDCT_US|Rhabdosarcoma|8900/3
C0334480|T191|PT|0000029993|CHV|pleomorphic rhabdomyosarcoma|8901/3
C0334480|T191|SY|0000029993|CHV|rhabdomyosarcoma pleomorphic|8901/3
C0334480|T191|PT|MTHU060031|ICPC2ICD10ENG|pleomorphic; rhabdomyosarcoma|8901/3
C0334480|T191|PT|MTHU064737|ICPC2ICD10ENG|rhabdomyosarcoma; pleomorphic|8901/3
C0334480|T191|PT|271525|MEDCIN|adult type pleomorphic rhabdomyosarcoma|8901/3
C0334480|T191|SY|271525|MEDCIN|malignant myosarcoma rhabdomyosarcoma pleomorphic adult type|8901/3
C0334480|T191|SY|271525|MEDCIN|pleomorphic, adult type rhabdomyosarcoma|8901/3
C0334480|T191|PN|NOCODE|MTH|Pleomorphic Rhabdomyosarcoma|8901/3
C1332211|T191|PT|C27369|NCI|Adult Pleomorphic Rhabdomyosarcoma|8901/3
C0334480|T191|PT|C4258|NCI|Pleomorphic Rhabdomyosarcoma|8901/3
C0334480|T191|PT|BBK32|RCD|Pleomorphic rhabdomyosarcoma|8901/3
C0334480|T191|PT|77455004|SNOMEDCT_US|Pleomorphic rhabdomyosarcoma|8901/3
C0334480|T191|PT|404054005|SNOMEDCT_US|Pleomorphic rhabdomyosarcoma|8901/3
C0334480|T191|SY|77455004|SNOMEDCT_US|Pleomorphic rhabdomyosarcoma, adult type|8901/3
C0334481|T191|PT|MTHU064736|ICPC2ICD10ENG|rhabdomyosarcoma; mixed type|8902/3
C0334481|T191|SY|271526|MEDCIN|malignant neoplasm myosarcoma rhabdomyosarcoma mixed type|8902/3
C0334481|T191|PT|271526|MEDCIN|mixed type rhabdomyosarcoma|8902/3
C1709053|T191|PN|NOCODE|MTH|Rhabdomyosarcoma with Mixed Embryonal and Alveolar Features|8902/3
C1709053|T191|SY|C4259|NCI|Mixed Alveolar Rhabdomyosarcoma|8902/3
C1709053|T191|SY|C4259|NCI|Mixed Type Alveolar Rhabdomyosarcoma|8902/3
C1709053|T191|PT|C4259|NCI|Rhabdomyosarcoma with Mixed Embryonal and Alveolar Features|8902/3
C0334481|T191|PT|BBK33|RCD|Mixed type rhabdomyosarcoma|8902/3
C0334481|T191|SY|62383007|SNOMEDCT_US|Mixed embryonal rhabdomyosarcoma and alveolar rhabdomyosarcoma|8902/3
C0334481|T191|PT|62383007|SNOMEDCT_US|Mixed type rhabdomyosarcoma|8902/3
C0334482|T191|PT|MTHU029075|ICPC2ICD10ENG|fetal; rhabdomyoma|8903/0
C0334482|T191|PT|MTHU064731|ICPC2ICD10ENG|rhabdomyoma; fetal|8903/0
C0334482|T191|PT|C4260|NCI|Fetal Rhabdomyoma|8903/0
C0334482|T191|PT|BBK34|RCD|Fetal rhabdomyoma|8903/0
C0334482|T191|PT|404049001|SNOMEDCT_US|Fetal rhabdomyoma|8903/0
C0334482|T191|PT|40123003|SNOMEDCT_US|Fetal rhabdomyoma|8903/0
C0334482|T191|SY|404049001|SNOMEDCT_US|Foetal rhabdomyoma|8903/0
C0334482|T191|SY|40123003|SNOMEDCT_US|Foetal rhabdomyoma|8903/0
C4055487|T191|PT|C4261|NCI|Adult Extracardiac Rhabdomyoma|8904/0
C4055487|T191|SY|C4261|NCI|Adult Extracardiac Rhabdomyomatous Hamartoma|8904/0
C0334483|T191|PT|BBK35|RCD|Adult rhabdomyoma|8904/0
C0334483|T191|SY|BBK35|RCD|Glycogenic rhabdomyoma|8904/0
C0334483|T191|PT|404048009|SNOMEDCT_US|Adult rhabdomyoma|8904/0
C0334483|T191|PT|16107003|SNOMEDCT_US|Adult rhabdomyoma|8904/0
C0334483|T191|SY|16107003|SNOMEDCT_US|Glycogenic rhabdomyoma|8904/0
C1266133|T191|PT|C6517|NCI|Genital Rhabdomyoma|8905/0
C1266133|T191|PT|128748000|SNOMEDCT_US|Genital rhabdomyoma|8905/0
C1266133|T191|PT|404050001|SNOMEDCT_US|Genital rhabdomyoma|8905/0
C1266133|T191|SY|128748000|SNOMEDCT_US|Genital type rhabdomyoma|8905/0
C0206656|T191|PT|0000021000|CHV|embryonal rhabdomyosarcoma|8910/3
C0206656|T191|PT|HP:0006743|HPO|Embryonal rhabdomyosarcoma|8910/3
C1306573|T191|PT|MTHU012345|ICPC2ICD10ENG|botryoid; sarcoma|8910/3
C0206656|T191|PT|MTHU025480|ICPC2ICD10ENG|embryonal; rhabdomyosarcoma|8910/3
C0206656|T191|PT|MTHU064735|ICPC2ICD10ENG|rhabdomyosarcoma; embryonal|8910/3
C1306573|T191|PT|MTHU065888|ICPC2ICD10ENG|sarcoma; botryoid|8910/3
C0206656|T191|LLT|10065868|MDR|Embryonal rhabdomyosarcoma|8910/3
C0206656|T191|PT|10065868|MDR|Embryonal rhabdomyosarcoma|8910/3
C1306573|T191|LLT|10078566|MDR|Sarcoma botryoides|8910/3
C0206656|T191|PT|271527|MEDCIN|embryonal rhabdomyosarcoma|8910/3
C0206656|T191|SY|271527|MEDCIN|malignant neoplasm myosarcoma rhabdomyosarcoma embryonal|8910/3
C0206656|T191|PM|D018233|MSH|Embryonal Rhabdomyosarcoma|8910/3
C0206656|T191|PM|D018233|MSH|Embryonal Rhabdomyosarcomas|8910/3
C0206656|T191|MH|D018233|MSH|Rhabdomyosarcoma, Embryonal|8910/3
C0206656|T191|PM|D018233|MSH|Rhabdomyosarcomas, Embryonal|8910/3
C1306573|T191|PN|NOCODE|MTH|Botryoid-Type Embryonal Rhabdomyosarcoma|8910/3
C0206656|T191|PN|NOCODE|MTH|Embryonal Rhabdomyosarcoma|8910/3
C1306573|T191|SY|C9150|NCI|Botryoid Sarcoma|8910/3
C1306573|T191|PT|C9150|NCI|Botryoid-Type Embryonal Rhabdomyosarcoma|8910/3
C0206656|T191|PT|C8971|NCI|Embryonal Rhabdomyosarcoma|8910/3
C1306573|T191|SY|C9150|NCI|Sarcoma Botryoides|8910/3
C0206656|T191|PT|10065868|NCI_CTEP-SDC|Embryonal rhabdomyosarcoma|8910/3
C0206656|T191|PT|CDR0000044497|NCI_NCI-GLOSS|embryonal rhabdomyosarcoma|8910/3
C0206656|T191|PT|CDR0000641930|NCI_NCI-GLOSS|ERMS|8910/3
C1306573|T191|SY|BBK36|RCD|Botryoid sarcoma|8910/3
C0206656|T191|PT|BBK36|RCD|Embryonal rhabdomyosarcoma|8910/3
C1306573|T191|SY|BBK36|RCD|Sarcoma botryoides|8910/3
C1306573|T191|SY|14269005|SNOMEDCT_US|Botryoid sarcoma|8910/3
C1306573|T191|PT|405943005|SNOMEDCT_US|Botryoid sarcoma|8910/3
C0206656|T191|PT|404051002|SNOMEDCT_US|Embryonal rhabdomyosarcoma|8910/3
C0206656|T191|PT|14269005|SNOMEDCT_US|Embryonal rhabdomyosarcoma|8910/3
C1306573|T191|SY|404052009|SNOMEDCT_US|Sarcoma botryoides|8910/3
C1306573|T191|SY|405943005|SNOMEDCT_US|Sarcoma botryoides|8910/3
C1306573|T191|SY|14269005|SNOMEDCT_US|Sarcoma botryoides|8910/3
C1266134|T191|SY|271528|MEDCIN|malignant neoplasm myosarcoma rhabdomyosarcoma spindle cell|8912/3
C1266134|T191|PT|271528|MEDCIN|spindle cell rhabdomyosarcoma|8912/3
C1266134|T191|PT|C6519|NCI|Spindle Cell Rhabdomyosarcoma|8912/3
C1266134|T191|PT|C6519|NCI_NICHD|Spindle Cell Rhabdomyosarcoma|8912/3
C1266134|T191|PT|CDR0000776840|PDQ|spindle cell rhabdomyosarcoma|8912/3
C1266134|T191|PT|404055006|SNOMEDCT_US|Spindle cell rhabdomyosarcoma|8912/3
C1266134|T191|PT|128749008|SNOMEDCT_US|Spindle cell rhabdomyosarcoma|8912/3
C0206655|T191|PT|0000020999|CHV|alveolar rhabdomyosarcoma|8920/3
C0206655|T191|SY|0000020999|CHV|alveolar rhabdomyosarcomas|8920/3
C0206655|T191|PT|HP:0006779|HPO|Alveolar rhabdomyosarcoma|8920/3
C0206655|T191|PT|MTHU005107|ICPC2ICD10ENG|alveolar; rhabdomyosarcoma|8920/3
C0206655|T191|PT|MTHU064734|ICPC2ICD10ENG|rhabdomyosarcoma; alveolar|8920/3
C0206655|T191|PT|10065867|MDR|Alveolar rhabdomyosarcoma|8920/3
C0206655|T191|LLT|10065867|MDR|Alveolar rhabdomyosarcoma|8920/3
C0206655|T191|PT|271534|MEDCIN|alveolar rhabdomyosarcoma|8920/3
C0206655|T191|SY|271534|MEDCIN|malignant neoplasm myosarcoma rhabdomyosarcoma alveolar|8920/3
C0206655|T191|PM|D018232|MSH|Alveolar Rhabdomyosarcoma|8920/3
C0206655|T191|PM|D018232|MSH|Alveolar Rhabdomyosarcomas|8920/3
C0206655|T191|ET|D018232|MSH|Rhabdomyosarcoma 2|8920/3
C0206655|T191|MH|D018232|MSH|Rhabdomyosarcoma, Alveolar|8920/3
C0206655|T191|PM|D018232|MSH|Rhabdomyosarcomas, Alveolar|8920/3
C0206655|T191|PN|NOCODE|MTH|Alveolar rhabdomyosarcoma|8920/3
C0206655|T191|PT|C3749|NCI|Alveolar Rhabdomyosarcoma|8920/3
C0206655|T191|AB|C3749|NCI|ARMS|8920/3
C0206655|T191|SY|C3749|NCI|Monomorphous Round Cell Rhabdomyosarcoma|8920/3
C0206655|T191|PT|10065867|NCI_CTEP-SDC|Alveolar rhabdomyosarcoma|8920/3
C0206655|T191|PT|CDR0000641927|NCI_NCI-GLOSS|alveolar rhabdomyosarcoma|8920/3
C0206655|T191|PT|CDR0000641928|NCI_NCI-GLOSS|ARMS|8920/3
C0206655|T191|PT|BBK37|RCD|Alveolar rhabdomyosarcoma|8920/3
C0206655|T191|PT|404053004|SNOMEDCT_US|Alveolar rhabdomyosarcoma|8920/3
C0206655|T191|PT|63449009|SNOMEDCT_US|Alveolar rhabdomyosarcoma|8920/3
C0431111|T191|PT|271535|MEDCIN|rhabdomyosarcoma with ganglionic differentiation|8921/3
C0431111|T191|PT|C4716|NCI|Ectomesenchymoma|8921/3
C0431111|T191|SY|C4716|NCI|Malignant Ectomesenchymoma|8921/3
C0431111|T191|SY|C4716|NCI|Sarcoma with Ganglionic or Neuroectodermal Differentiation|8921/3
C0431111|T191|PT|CDR0000518306|NCI_NCI-GLOSS|ectomesenchymoma|8921/3
C0431111|T191|PT|CDR0000539499|NCI_NCI-GLOSS|malignant ectomesenchymoma|8921/3
C0431111|T191|SY|X77pW|RCD|Ectomesenchymoma|8921/3
C0431111|T191|PT|X77pW|RCD|Gangliorhabdomyosarcoma|8921/3
C0431111|T191|SY|128750008|SNOMEDCT_US|Ectomesenchymoma|8921/3
C0431111|T191|SY|128750008|SNOMEDCT_US|Gangliorhabdomyosarcoma|8921/3
C0431111|T191|PT|128750008|SNOMEDCT_US|Rhabdomyosarcoma with ganglionic differentiation|8921/3
C0334485|T191|PN|NOCODE|MTH|Endometrial stromal nodule|8930/0
C0334485|T191|PT|C4262|NCI|Endometrial Stromal Nodule|8930/0
C0334485|T191|PT|X77oq|RCD|Endometrial stromal nodule|8930/0
C0334485|T191|OF|189810002|SNOMEDCT_US|Endometrial stromal nodule|8930/0
C0334485|T191|PT|70971005|SNOMEDCT_US|Endometrial stromal nodule|8930/0
C0334485|T191|OAP|189810002|SNOMEDCT_US|Endometrial stromal nodule|8930/0
C0206630|T191|SY|0000020980|CHV|endometrial sarcoma|8930/3
C0206630|T191|PT|0000020980|CHV|endometrial stromal sarcoma|8930/3
C0206630|T191|SY|0000020980|CHV|endometrial stromal sarcomas|8930/3
C0206630|T191|SY|0000020980|CHV|sarcoma endometrium|8930/3
C0206630|T191|SY|0000020980|CHV|sarcoma stromal|8930/3
C0206630|T191|SY|0000020980|CHV|stromal sarcoma|8930/3
C0206630|T191|PT|10048397|MDR|Endometrial stromal sarcoma|8930/3
C0206630|T191|LLT|10048397|MDR|Endometrial stromal sarcoma|8930/3
C0206630|T191|ET|D018203|MSH|Endometrial Stromal Sarcoma|8930/3
C0206630|T191|PM|D018203|MSH|Endometrial Stromal Sarcomas|8930/3
C0206630|T191|MH|D018203|MSH|Sarcoma, Endometrial Stromal|8930/3
C0206630|T191|PM|D018203|MSH|Sarcomas, Endometrial Stromal|8930/3
C0206630|T191|PM|D018203|MSH|Stromal Sarcoma, Endometrial|8930/3
C0206630|T191|PM|D018203|MSH|Stromal Sarcomas, Endometrial|8930/3
C0206630|T191|PN|NOCODE|MTH|Endometrial Stromal Sarcoma|8930/3
C2239246|T191|PN|NOCODE|MTH|Endometrial stromal sarcoma, high grade|8930/3
C0206630|T191|SY|C8973|NCI|Endometrial Stromal Sarcoma|8930/3
C0206630|T191|PT|C8973|NCI|Endometrioid Stromal Sarcoma|8930/3
C0206630|T191|AB|C8973|NCI|ESS|8930/3
C2239246|T191|SY|C8972|NCI|Undifferentiated Uterine Sarcoma|8930/3
C2239246|T191|SY|C8972|NCI|Uterine Corpus Undifferentiated Endometrial Sarcoma|8930/3
C2239246|T191|PT|C8972|NCI|Uterine Corpus Undifferentiated Sarcoma|8930/3
C0206630|T191|SY|C8973|NCI_CDISC|ESS|8930/3
C0206630|T191|PT|C8973|NCI_CDISC|STROMAL SARCOMA, ENDOMETRIAL, MALIGNANT|8930/3
C0206630|T191|PT|10048397|NCI_CTEP-SDC|Endometrial stromal sarcoma|8930/3
C0206630|T191|DN|C8973|NCI_CTRP|Endometrioid Stromal Sarcoma|8930/3
C0206630|T191|PT|CDR0000041019|PDQ|endometrial stromal sarcoma|8930/3
C0206630|T191|AB|CDR0000041019|PDQ|ESS|8930/3
C0206630|T191|SY|CDR0000041019|PDQ|stromal sarcoma, endometrial|8930/3
C0206630|T191|SY|BBL0.|RCD|Endometrial sarcoma|8930/3
C0206630|T191|PT|BBL0.|RCD|Endometrial stromal sarcoma|8930/3
C0206630|T191|SY|BBL0.|RCD|Stromal sarcoma|8930/3
C0206630|T191|SY|70555003|SNOMEDCT_US|Endometrial sarcoma|8930/3
C0206630|T191|IS|70555003|SNOMEDCT_US|Endometrial sarcoma, NOS|8930/3
C0206630|T191|PT|699356008|SNOMEDCT_US|Endometrial stromal sarcoma|8930/3
C0206630|T191|SY|70555003|SNOMEDCT_US|Endometrial stromal sarcoma|8930/3
C2959946|T191|PT|446578007|SNOMEDCT_US|Endometrial stromal sarcoma - category|8930/3
C2239246|T191|PT|70555003|SNOMEDCT_US|Endometrial stromal sarcoma, high grade|8930/3
C2239246|T191|SY|70555003|SNOMEDCT_US|Endometrioid stromal sarcoma, high grade|8930/3
C2239246|T191|PT|699358009|SNOMEDCT_US|High grade endometrial stromal sarcoma|8930/3
C0206630|T191|SY|699356008|SNOMEDCT_US|Primary malignant stromal sarcoma of endometrium|8930/3
C0206630|T191|IS|70555003|SNOMEDCT_US|Stromal sarcoma, NOS|8930/3
C0334486|T191|SY|0000029994|CHV|endolymphatic stromal myosis|8931/3
C0334486|T191|PT|0000029994|CHV|stromal myosis|8931/3
C0334486|T191|PT|MTHU026117|ICPC2ICD10ENG|endometriosis; stromal|8931/3
C0334486|T191|PT|MTHU051224|ICPC2ICD10ENG|myosis; stromal|8931/3
C0334486|T191|PT|MTHU070955|ICPC2ICD10ENG|stromal; endometriosis|8931/3
C0334486|T191|PT|MTHU070956|ICPC2ICD10ENG|stromal; myosis|8931/3
C0334486|T191|PT|MTHU070959|ICPC2ICD10ENG|stromatosis; endometrial|8931/3
C0334486|T191|PM|D036821|MSH|Endolymphatic Stromal Myoses|8931/3
C0334486|T191|ET|D036821|MSH|Endolymphatic Stromal Myosis|8931/3
C0334486|T191|PM|D036821|MSH|Myoses, Endolymphatic Stromal|8931/3
C0334486|T191|PM|D036821|MSH|Myosis, Endolymphatic Stromal|8931/3
C0334486|T191|PEP|D036821|MSH|Sarcoma, Endometrial Stromal, Low-Grade|8931/3
C0334486|T191|PM|D036821|MSH|Stromal Myoses, Endolymphatic|8931/3
C0334486|T191|PM|D036821|MSH|Stromal Myosis, Endolymphatic|8931/3
C0334486|T191|PN|NOCODE|MTH|Low Grade Endometrial Stromal Sarcoma|8931/3
C0334486|T191|SY|C4263|NCI|Endolymphatic Stromal Myosis|8931/3
C0334486|T191|PT|C4263|NCI|Low Grade Endometrioid Stromal Sarcoma|8931/3
C0334486|T191|PT|BBL1.|RCD|Endolymphatic stromal myosis|8931/3
C0334486|T191|SY|BBL1.|RCD|Endometrial stromatosis|8931/3
C0334486|T191|SY|BBL1.|RCD|Stromal endometriosis|8931/3
C0334486|T191|SY|BBL1.|RCD|Stromal myosis|8931/3
C0334486|T191|OAP|81158008|SNOMEDCT_US|Endolymphatic stromal myosis|8931/3
C0334486|T191|SY|128726006|SNOMEDCT_US|Endolymphatic stromal myosis|8931/3
C0334486|T191|IS|81158008|SNOMEDCT_US|Endolymphatic stromal myosis -RETIRED-|8931/3
C0334486|T191|OF|81158008|SNOMEDCT_US|Endolymphatic stromal myosis -RETIRED-|8931/3
C0334486|T191|PT|128726006|SNOMEDCT_US|Endometrial stromal sarcoma, low grade|8931/3
C0334486|T191|IS|81158008|SNOMEDCT_US|Endometrial stromatosis|8931/3
C0334486|T191|SY|128726006|SNOMEDCT_US|Endometrial stromatosis|8931/3
C0334486|T191|SY|128726006|SNOMEDCT_US|Endometrioid stromal sarcoma, low grade|8931/3
C0334486|T191|PT|699357004|SNOMEDCT_US|Low grade endometrial stromal sarcoma|8931/3
C0334486|T191|IS|81158008|SNOMEDCT_US|Stromal endometriosis|8931/3
C0334486|T191|SY|128726006|SNOMEDCT_US|Stromal endometriosis|8931/3
C0334486|T191|SY|128726006|SNOMEDCT_US|Stromal myosis|8931/3
C0334486|T191|IS|81158008|SNOMEDCT_US|Stromal myosis, NOS|8931/3
C0206622|T191|PT|0000020974|CHV|adenomyoma|8932/0
C0206622|T191|LLT|10063549|MDR|Adenomyoma|8932/0
C0206622|T191|MH|D018194|MSH|Adenomyoma|8932/0
C0206622|T191|PM|D018194|MSH|Adenomyomas|8932/0
C0206622|T191|PT|C3726|NCI|Adenomyoma|8932/0
C1300347|T191|PT|C6895|NCI|Atypical Polypoid Adenomyoma|8932/0
C0206622|T191|PT|C3726|NCI_CDISC|ADENOMYOMA, BENIGN|8932/0
C0206622|T191|PT|BBL2.|RCD|Adenomyoma|8932/0
C0206622|T191|PT|40293003|SNOMEDCT_US|Adenomyoma|8932/0
C1300347|T191|PT|388987001|SNOMEDCT_US|Atypical polypoid adenomyoma|8932/0
C1300347|T191|SY|40293003|SNOMEDCT_US|Atypical polypoid adenomyoma|8932/0
C0001442|T191|PT|0000000719|CHV|adenosarcoma|8933/3
C0001442|T191|MH|D018195|MSH|Adenosarcoma|8933/3
C0001442|T191|PM|D018195|MSH|Adenosarcomas|8933/3
C0001442|T191|PN|NOCODE|MTH|Adenosarcoma|8933/3
C0001442|T191|PT|C9474|NCI|Adenosarcoma|8933/3
C0001442|T191|SY|C9474|NCI|Mullerian Adenosarcoma|8933/3
C0001442|T191|PT|C9474|NCI_CTRP|Adenosarcoma|8933/3
C0001442|T191|DN|C9474|NCI_CTRP|Adenosarcoma|8933/3
C0001442|T191|PT|CDR0000641990|NCI_NCI-GLOSS|adenosarcoma|8933/3
C0001442|T191|PT|BBLE.|RCD|Adenosarcoma|8933/3
C0001442|T191|OAP|189804002|SNOMEDCT_US|Adenosarcoma|8933/3
C0001442|T191|OF|189804002|SNOMEDCT_US|Adenosarcoma|8933/3
C0001442|T191|PT|31470003|SNOMEDCT_US|Adenosarcoma|8933/3
C1266135|T191|PT|271536|MEDCIN|carcinofibroma|8934/3
C1883485|T191|PT|C40182|NCI|Uterine Corpus Carcinofibroma|8934/3
C1266135|T191|PT|128751007|SNOMEDCT_US|Carcinofibroma|8934/3
C0474833|T191|ET|D21|ICD10CM|benign stromal tumors|8935/0
C0474833|T191|OP|C66772|NCI|Benign Stromal Tumor|8935/0
C0474833|T191|PT|C66772|NCI|Benign Stromal Tumor|8935/0
C0474833|T191|PT|X77op|RCD|Benign stromal tumour|8935/0
C0474833|T191|PT|X77op|RCDAE|Benign stromal tumor|8935/0
C0474833|T191|OAP|253049000|SNOMEDCT_US|Benign stromal tumor|8935/0
C0474833|T191|PT|447644002|SNOMEDCT_US|Benign stromal tumor|8935/0
C0474833|T191|OAP|253049000|SNOMEDCT_US|Benign stromal tumour|8935/0
C0474833|T191|PTGB|447644002|SNOMEDCT_US|Benign stromal tumour|8935/0
C0879615|T191|PT|0000052059|CHV|stromal tumor|8935/1
C0879615|T191|SY|0000052059|CHV|stromal tumors|8935/1
C0879615|T191|SY|0000052059|CHV|stromal tumour|8935/1
C0879615|T191|SY|0000052059|CHV|stromal tumours|8935/1
C0879615|T191|SY|0000052059|CHV|tumor stromal|8935/1
C0879615|T191|SY|0000052059|CHV|tumors stromal|8935/1
C0334695|T191|PM|D036821|MSH|Endometrial Stromal Tumor|8935/1
C0334695|T191|MH|D036821|MSH|Endometrial Stromal Tumors|8935/1
C0334695|T191|PM|D036821|MSH|Stromal Tumor, Endometrial|8935/1
C0334695|T191|PM|D036821|MSH|Stromal Tumors, Endometrial|8935/1
C0334695|T191|PM|D036821|MSH|Tumor, Endometrial Stromal|8935/1
C0334695|T191|PM|D036821|MSH|Tumors, Endometrial Stromal|8935/1
C0879615|T191|PN|NOCODE|MTH|Stromal Neoplasm|8935/1
C1285519|T191|PT|C157749|NCI|Metanephric Stromal Tumor|8935/1
C0879615|T191|SY|C6781|NCI|Stromal Cell Tumor|8935/1
C0879615|T191|PT|C6781|NCI|Stromal Neoplasm|8935/1
C0879615|T191|SY|C6781|NCI|Stromal Tumor|8935/1
C0879615|T191|PT|CDR0000044929|NCI_NCI-GLOSS|stromal tumor|8935/1
C0334695|T191|PT|446887007|SNOMEDCT_US|Endometrial stromal tumor|8935/1
C0334695|T191|PT|68738004|SNOMEDCT_US|Endometrial stromal tumor|8935/1
C0334695|T191|IS|68738004|SNOMEDCT_US|Endometrial stromal tumor, NOS|8935/1
C0334695|T191|PTGB|446887007|SNOMEDCT_US|Endometrial stromal tumour|8935/1
C0334695|T191|PTGB|68738004|SNOMEDCT_US|Endometrial stromal tumour|8935/1
C1285519|T191|PT|363658005|SNOMEDCT_US|Metanephric stromal tumor|8935/1
C1285519|T191|PTGB|363658005|SNOMEDCT_US|Metanephric stromal tumour|8935/1
C0879615|T191|PT|128752000|SNOMEDCT_US|Stromal tumor|8935/1
C0879615|T191|PTGB|128752000|SNOMEDCT_US|Stromal tumour|8935/1
C1370723|T191|PT|MTHU065934|ICPC2ICD10ENG|sarcoma; stromal|8935/3
C1370723|T191|PT|MTHU070957|ICPC2ICD10ENG|stromal; sarcoma|8935/3
C1370723|T191|PT|271499|MEDCIN|stromal sarcoma|8935/3
C1370723|T191|PN|NOCODE|MTH|Stromal sarcoma|8935/3
C1370723|T191|PT|C6926|NCI|Stromal Sarcoma|8935/3
C1370723|T191|PT|C6926|NCI_CDISC|STROMAL SARCOMA, MALIGNANT|8935/3
C1370723|T191|SY|C6926|NCI_CDISC|Stromal Tumor, Malignant|8935/3
C1370723|T191|PT|X77oj|RCD|Malignant stromal tumour|8935/3
C1370723|T191|PT|X77oj|RCDAE|Malignant stromal tumor|8935/3
C1370723|T191|PT|253048008|SNOMEDCT_US|Malignant stromal tumor|8935/3
C1370723|T191|PTGB|253048008|SNOMEDCT_US|Malignant stromal tumour|8935/3
C1370723|T191|PT|128753005|SNOMEDCT_US|Stromal sarcoma|8935/3
C1266136|T191|PT|C53998|NCI|Benign Gastrointestinal Stromal Tumor|8936/0
C1266136|T191|PT|C53998|NCI_CDISC|GASTROINTESTINAL STROMAL TUMOR, BENIGN|8936/0
C1266136|T191|SY|C53998|NCI_CDISC|GIST, Benign|8936/0
C1266136|T191|PT|128754004|SNOMEDCT_US|Gastrointestinal stromal tumor, benign|8936/0
C1266136|T191|PTGB|128754004|SNOMEDCT_US|Gastrointestinal stromal tumour, benign|8936/0
C1266136|T191|SY|128754004|SNOMEDCT_US|GIST, benign|8936/0
C0238198|T191|PT|0030321|CCPSS|GASTROINTESTINAL TUMOR STROMAL|8936/1
C0238198|T191|SY|0000023965|CHV|gant|8936/1
C0238198|T191|SY|0000023965|CHV|gants|8936/1
C0238198|T191|SY|0000023965|CHV|gastrointestinal stromal tumor|8936/1
C0238198|T191|SY|0000023965|CHV|gastrointestinal stromal tumors|8936/1
C0238198|T191|SY|0000023965|CHV|gastrointestinal stromal tumour|8936/1
C0238198|T191|SY|0000023965|CHV|gastrointestinal stromal tumours|8936/1
C0238198|T191|PT|0000023965|CHV|gist|8936/1
C0238198|T191|SY|0000023965|CHV|gists|8936/1
C0238198|T191|PT|HP:0100723|HPO|Gastrointestinal stroma tumor|8936/1
C0238198|T191|SY|HP:0100723|HPO|Gastrointestinal stromal tumor|8936/1
C0238198|T191|ET|HP:0100723|HPO|Gastrointestinal stromal tumors|8936/1
C0238198|T191|SY|HP:0100723|HPO|GI stroma tumor|8936/1
C0238198|T191|SY|HP:0100723|HPO|GIST|8936/1
C0238198|T191|AB|C49.A|ICD10CM|Gastrointestinal stromal tumor|8936/1
C0238198|T191|HT|C49.A|ICD10CM|Gastrointestinal stromal tumor|8936/1
C0238198|T191|PT|sh2006007119|LCH_NW|Gastrointestinal stromal tumors|8936/1
C0238198|T191|MTH_PT|10051066|MDR|Gastrointestinal stromal tumor|8936/1
C0238198|T191|LLT|10062427|MDR|Gastrointestinal stromal tumor|8936/1
C0238198|T191|LLT|10051066|MDR|Gastrointestinal stromal tumour|8936/1
C0238198|T191|PT|10051066|MDR|Gastrointestinal stromal tumour|8936/1
C0238198|T191|PT|355286|MEDCIN|gastrointestinal stromal neoplasm|8936/1
C0238198|T191|SY|355286|MEDCIN|neoplasm gastrointestinal tract stromal|8936/1
C0238198|T191|ET|3652|MEDLINEPLUS|Gastrointestinal Stromal Tumors|8936/1
C0238198|T191|ET|D046152|MSH|Gastrointestinal Stromal Neoplasm|8936/1
C0238198|T191|ET|D046152|MSH|Gastrointestinal Stromal Neoplasms|8936/1
C0238198|T191|ET|D046152|MSH|Gastrointestinal Stromal Tumor|8936/1
C0238198|T191|MH|D046152|MSH|Gastrointestinal Stromal Tumors|8936/1
C0238198|T191|PM|D046152|MSH|Neoplasm, Gastrointestinal Stromal|8936/1
C0238198|T191|PM|D046152|MSH|Neoplasms, Gastrointestinal Stromal|8936/1
C0238198|T191|PM|D046152|MSH|Stromal Neoplasm, Gastrointestinal|8936/1
C0238198|T191|PM|D046152|MSH|Stromal Neoplasms, Gastrointestinal|8936/1
C0238198|T191|PM|D046152|MSH|Stromal Tumor, Gastrointestinal|8936/1
C0238198|T191|PM|D046152|MSH|Stromal Tumors, Gastrointestinal|8936/1
C0238198|T191|PM|D046152|MSH|Tumor, Gastrointestinal Stromal|8936/1
C0238198|T191|PM|D046152|MSH|Tumors, Gastrointestinal Stromal|8936/1
C0238198|T191|PN|NOCODE|MTH|Gastrointestinal Stromal Tumors|8936/1
C0238198|T191|SY|C3868|NCI|Gastrointestinal Stromal Neoplasm|8936/1
C0238198|T191|PT|C3868|NCI|Gastrointestinal Stromal Tumor|8936/1
C1704399|T191|HD|C54000|NCI|Gastrointestinal Stromal Tumor of Uncertain Malignant Potential|8936/1
C1704399|T191|PT|C54000|NCI|Gastrointestinal Stromal Tumor of Uncertain Malignant Potential|8936/1
C0238198|T191|AB|C3868|NCI|GIST|8936/1
C0238198|T191|PT|C3868|NCI_CPTAC|Gastrointestinal Stromal Tumor|8936/1
C0238198|T191|PT|10051066|NCI_CTEP-SDC|Gastrointestinal stromal tumor|8936/1
C0238198|T191|PT|CDR0000044998|NCI_NCI-GLOSS|gastrointestinal stromal tumor|8936/1
C0238198|T191|PT|CDR0000044406|NCI_NCI-GLOSS|GIST|8936/1
C0238198|T191|PSC|CDR0000038161|PDQ|gastrointestinal stromal tumor|8936/1
C0238198|T191|AB|CDR0000038161|PDQ|GIST|8936/1
C0238198|T191|SY|CDR0000038161|PDQ|stromal tumor, gastrointestinal|8936/1
C0238198|T191|SY|128755003|SNOMEDCT_US|Gastrointestinal pacemaker cell tumor|8936/1
C0238198|T191|SYGB|128755003|SNOMEDCT_US|Gastrointestinal pacemaker cell tumour|8936/1
C0238198|T191|SY|128755003|SNOMEDCT_US|Gastrointestinal stromal tumor|8936/1
C0238198|T191|PT|420120006|SNOMEDCT_US|Gastrointestinal stromal tumor|8936/1
C1704399|T191|PT|128755003|SNOMEDCT_US|Gastrointestinal stromal tumor, uncertain malignant potential|8936/1
C0238198|T191|SYGB|128755003|SNOMEDCT_US|Gastrointestinal stromal tumour|8936/1
C0238198|T191|PTGB|420120006|SNOMEDCT_US|Gastrointestinal stromal tumour|8936/1
C1704399|T191|PTGB|128755003|SNOMEDCT_US|Gastrointestinal stromal tumour, uncertain malignant potential|8936/1
C0238198|T191|SY|128755003|SNOMEDCT_US|GIST|8936/1
C0238198|T191|SY|420120006|SNOMEDCT_US|GIST - Gastrointestinal stromal tumor|8936/1
C0238198|T191|SYGB|420120006|SNOMEDCT_US|GIST - Gastrointestinal stromal tumour|8936/1
C3179349|T191|LA|LA26516-7|LNC|Gastrointestinal stromal tumor, malignant|8936/3
C3179349|T191|PEP|D046152|MSH|Gastrointestinal Stromal Sarcoma|8936/3
C3179349|T191|PT|C53999|NCI|Malignant Gastrointestinal Stromal Tumor|8936/3
C3179349|T191|PT|C53999|NCI_CDISC|GASTROINTESTINAL STROMA TUMOR, MALIGNANT|8936/3
C3179349|T191|SY|C53999|NCI_CDISC|GIST, Malignant|8936/3
C3179349|T191|SY|420120006|SNOMEDCT_US|Gastrointestinal stromal sarcoma|8936/3
C3179349|T191|PT|128756002|SNOMEDCT_US|Gastrointestinal stromal sarcoma|8936/3
C3179349|T191|SY|128756002|SNOMEDCT_US|Gastrointestinal stromal tumor, malignant|8936/3
C3179349|T191|SYGB|128756002|SNOMEDCT_US|Gastrointestinal stromal tumour, malignant|8936/3
C3179349|T191|SY|128756002|SNOMEDCT_US|GIST, malignant|8936/3
C0026277|T191|SY|0000008198|CHV|adenoma pleomorphic|8940/0
C0026277|T191|SY|0000008198|CHV|chondroid syringoma|8940/0
C0026277|T191|SY|0000008198|CHV|mixed tumor|8940/0
C0026277|T191|SY|0000008198|CHV|mixed tumors|8940/0
C0026277|T191|PT|0000008198|CHV|pleomorphic adenoma|8940/0
C0026277|T191|SY|0000008198|CHV|pleomorphic adenomas|8940/0
C0026277|T191|SY|0000008198|CHV|tumor mix|8940/0
C0026277|T191|SY|0000008198|CHV|tumour mix|8940/0
C0026277|T191|PT|MTHU016347|ICPC2ICD10ENG|chondroid; syringoma|8940/0
C0026277|T191|PT|MTHU073180|ICPC2ICD10ENG|syringoma; chondroid|8940/0
C0026277|T191|PT|10073372|MDR|Pleomorphic adenoma|8940/0
C0026277|T191|LLT|10073372|MDR|Pleomorphic adenoma|8940/0
C0026277|T191|MH|D008949|MSH|Adenoma, Pleomorphic|8940/0
C0026277|T191|PM|D008949|MSH|Adenomas, Pleomorphic|8940/0
C0026277|T191|PM|D008949|MSH|Chondroid Syringoma|8940/0
C0026277|T191|PM|D008949|MSH|Chondroid Syringomas|8940/0
C0026277|T191|ET|D008949|MSH|Mixed Salivary Gland Tumor|8940/0
C0026277|T191|PM|D008949|MSH|Pleomorphic Adenoma|8940/0
C0026277|T191|PM|D008949|MSH|Pleomorphic Adenomas|8940/0
C0026277|T191|ET|D008949|MSH|Salivary Gland Tumor, Mixed|8940/0
C0026277|T191|ET|D008949|MSH|Syringoma, Chondroid|8940/0
C0026277|T191|PM|D008949|MSH|Syringomas, Chondroid|8940/0
C0346026|T191|PN|NOCODE|MTH|Eccrine mixed tumor of skin|8940/0
C0026277|T191|PN|NOCODE|MTH|Mixed Salivary Gland Tumor|8940/0
C0346026|T191|SY|C4474|NCI|Benign Mixed Tumor of Skin|8940/0
C0346026|T191|SY|C4474|NCI|Benign Mixed Tumor of the Skin|8940/0
C0346026|T191|SY|C4474|NCI|Chondroid Syringoma|8940/0
C0026277|T191|SY|C35691|NCI|Mixed Tumor of Salivary Gland|8940/0
C0026277|T191|PT|C35691|NCI|Mixed Tumor of the Salivary Gland|8940/0
C0026277|T191|PT|C8602|NCI|Pleomorphic Adenoma|8940/0
C0026277|T191|PT|C8602|NCI_CDISC|TUMOR, MIXED, BENIGN|8940/0
C0026277|T191|SY|BBL3.|RCD|Chondroid syringoma|8940/0
C0346026|T191|PT|X78Sv|RCD|Eccrine mixed tumour|8940/0
C0026277|T191|SY|BBL3.|RCD|Mixed salivary gland tumour|8940/0
C0026277|T191|SY|BBL3.|RCD|Mixed tumour|8940/0
C0346026|T191|SY|X78Sv|RCD|Mixed tumour of skin|8940/0
C0026277|T191|PT|BBL3.|RCD|Pleomorphic adenoma|8940/0
C0346026|T191|PT|X78Sv|RCDAE|Eccrine mixed tumor|8940/0
C0026277|T191|SY|BBL3.|RCDAE|Mixed salivary gland tumor|8940/0
C0026277|T191|SY|BBL3.|RCDAE|Mixed tumor|8940/0
C0346026|T191|SY|X78Sv|RCDAE|Mixed tumor of skin|8940/0
C0026277|T191|SY|8360001|SNOMEDCT_US|Chondroid syringoma|8940/0
C0346026|T191|PT|400144002|SNOMEDCT_US|Eccrine mixed tumor|8940/0
C0346026|T191|PT|254720009|SNOMEDCT_US|Eccrine mixed tumor|8940/0
C0346026|T191|SY|254720009|SNOMEDCT_US|Eccrine mixed tumor of skin|8940/0
C0346026|T191|PTGB|400144002|SNOMEDCT_US|Eccrine mixed tumour|8940/0
C0346026|T191|PTGB|254720009|SNOMEDCT_US|Eccrine mixed tumour|8940/0
C0346026|T191|SYGB|254720009|SNOMEDCT_US|Eccrine mixed tumour of skin|8940/0
C0026277|T191|SY|8360001|SNOMEDCT_US|Mixed salivary gland tumor|8940/0
C0026277|T191|SYGB|8360001|SNOMEDCT_US|Mixed salivary gland tumour|8940/0
C0026277|T191|SY|8360001|SNOMEDCT_US|Mixed tumor|8940/0
C0346026|T191|SY|254720009|SNOMEDCT_US|Mixed tumor of skin|8940/0
C0026277|T191|IS|8360001|SNOMEDCT_US|Mixed tumor, NOS|8940/0
C0026277|T191|SY|8360001|SNOMEDCT_US|Mixed tumor, salivary gland type|8940/0
C0026277|T191|IS|8360001|SNOMEDCT_US|Mixed tumor, salivary gland type, NOS|8940/0
C0026277|T191|SYGB|8360001|SNOMEDCT_US|Mixed tumour|8940/0
C0346026|T191|SYGB|254720009|SNOMEDCT_US|Mixed tumour of skin|8940/0
C0026277|T191|SYGB|8360001|SNOMEDCT_US|Mixed tumour, salivary gland type|8940/0
C0026277|T191|PT|8360001|SNOMEDCT_US|Pleomorphic adenoma|8940/0
C1368354|T191|PN|NOCODE|MTH|Mixed Neoplasm|8940/1
C1368354|T191|PT|C6930|NCI|Mixed Neoplasm|8940/1
C1368354|T191|SY|C6930|NCI|Mixed Tumor|8940/1
C0206625|T191|PT|MTHU031232|ICPC2ICD10ENG|mixed; tumor, malignant|8940/3
C0206625|T191|PT|MTHU077092|ICPC2ICD10ENG|tumor; malignant, mixed|8940/3
C0206625|T191|PT|MTHU077062|ICPC2ICD10ENG|tumor; mixed, malignant|8940/3
C0206625|T191|PT|271537|MEDCIN|malignant mixed tumor|8940/3
C1321781|T191|PT|231704|MEDCIN|malignant mixed tumor of skin|8940/3
C0206625|T191|PM|D018198|MSH|Malignant Mixed Tumor|8940/3
C0206625|T191|PM|D018198|MSH|Malignant Mixed Tumors|8940/3
C0206625|T191|MH|D018198|MSH|Mixed Tumor, Malignant|8940/3
C0206625|T191|PM|D018198|MSH|Mixed Tumors, Malignant|8940/3
C0206625|T191|PM|D018198|MSH|Tumor, Malignant Mixed|8940/3
C0206625|T191|PM|D018198|MSH|Tumors, Malignant Mixed|8940/3
C1321781|T191|PN|NOCODE|MTH|Malignant chondroid syringoma|8940/3
C0206625|T191|PN|U002408|MTH|Malignant Mixed Tumor|8940/3
C0206625|T191|PT|C3729|NCI|Malignant Mixed Neoplasm|8940/3
C0206625|T191|SY|C3729|NCI|Malignant Mixed Tumor|8940/3
C0206625|T191|SY|C3729|NCI_CDISC|Malignant Mixed Tumor|8940/3
C0206625|T191|PT|C3729|NCI_CDISC|TUMOR, MIXED, MALIGNANT|8940/3
C0206625|T191|PT|C3729|NCI_CPTAC|Malignant Mixed Neoplasm|8940/3
C0206625|T191|PT|XM1FO|RCD|Malignant mixed tumour|8940/3
C0206625|T191|PT|XM1FO|RCDAE|Malignant mixed tumor|8940/3
C0206625|T191|OA|BBL4.|RCDSA|Mixed tumor, malignant NOS|8940/3
C0206625|T191|OP|BBL4.|RCDSA|Mixed tumor, malignant, NOS|8940/3
C0206625|T191|OA|BBL4.|RCDSY|Mixed tumour, malignant NOS|8940/3
C0206625|T191|OP|BBL4.|RCDSY|Mixed tumour, malignant, NOS|8940/3
C1321781|T191|SY|403943008|SNOMEDCT_US|Eccrine mixed tumor, malignant|8940/3
C1321781|T191|SYGB|403943008|SNOMEDCT_US|Eccrine mixed tumour, malignant|8940/3
C1321781|T191|PT|400124008|SNOMEDCT_US|Malignant chondroid syringoma|8940/3
C1321781|T191|PT|403943008|SNOMEDCT_US|Malignant chondroid syringoma|8940/3
C1321781|T191|SY|8145008|SNOMEDCT_US|Malignant chondroid syringoma|8940/3
C1321781|T191|SY|403943008|SNOMEDCT_US|Malignant chondroid syringoma of skin|8940/3
C0206625|T191|SY|8145008|SNOMEDCT_US|Malignant mixed tumor|8940/3
C1321781|T191|SY|403943008|SNOMEDCT_US|Malignant mixed tumor of the skin|8940/3
C0334696|T191|PT|40459000|SNOMEDCT_US|Malignant mixed tumor, carcinomatous type|8940/3
C0334697|T191|PT|82993000|SNOMEDCT_US|Malignant mixed tumor, chondrosarcomatous type|8940/3
C0334698|T191|PT|4392007|SNOMEDCT_US|Malignant mixed tumor, osteosarcomatous type|8940/3
C0206625|T191|SYGB|8145008|SNOMEDCT_US|Malignant mixed tumour|8940/3
C1321781|T191|SYGB|403943008|SNOMEDCT_US|Malignant mixed tumour of the skin|8940/3
C0334696|T191|PTGB|40459000|SNOMEDCT_US|Malignant mixed tumour, carcinomatous type|8940/3
C0334697|T191|PTGB|82993000|SNOMEDCT_US|Malignant mixed tumour, chondrosarcomatous type|8940/3
C0334698|T191|PTGB|4392007|SNOMEDCT_US|Malignant mixed tumour, osteosarcomatous type|8940/3
C0206625|T191|PT|8145008|SNOMEDCT_US|Mixed tumor, malignant|8940/3
C0206625|T191|PTGB|8145008|SNOMEDCT_US|Mixed tumour, malignant|8940/3
C0344460|T191|LLT|10077435|MDR|Carcinoma ex-pleomorphic adenoma|8941/3
C0344460|T191|PT|10077435|MDR|Carcinoma ex-pleomorphic adenoma|8941/3
C0344460|T191|PT|271451|MEDCIN|carcinoma ex pleomorphic adenoma|8941/3
C0344460|T191|SY|271451|MEDCIN|malignant neoplasm carcinoma ex pleomorphic adenoma|8941/3
C0344460|T191|PT|C4397|NCI|Carcinoma ex Pleomorphic Adenoma|8941/3
C0344460|T191|SY|C4397|NCI|Carcinoma in Pleomorphic Adenoma|8941/3
C0344460|T191|AB|X77ok|RCD|Ca in pleomorphic adenoma|8941/3
C0344460|T191|PT|X77ok|RCD|Carcinoma in pleomorphic adenoma|8941/3
C0344460|T191|AB|X77ok|RCDSY|Carcin in pleomorph adenoma|8941/3
C0344460|T191|PT|17264009|SNOMEDCT_US|Carcinoma ex pleomorphic adenoma|8941/3
C0344460|T191|OAP|189811003|SNOMEDCT_US|Carcinoma in pleomorphic adenoma|8941/3
C0344460|T191|OF|189811003|SNOMEDCT_US|Carcinoma in pleomorphic adenoma|8941/3
C0344460|T191|SY|17264009|SNOMEDCT_US|Carcinoma in pleomorphic adenoma|8941/3
C3698226|T191|SY|698255000|SNOMEDCT_US|Intracapsular carcinoma ex pleomorphic adenoma|8941/3
C3698226|T191|PT|698255000|SNOMEDCT_US|Noninvasive carcinoma ex pleomorphic adenoma|8941/3
C0206627|T191|PT|0046136|CCPSS|MULLERIAN MIXED TUMOR|8950/3
C0206627|T191|PT|0000020977|CHV|mixed mullerian tumor|8950/3
C0206627|T191|SY|0000020977|CHV|mixed mullerian tumors|8950/3
C0206627|T191|SY|0000020977|CHV|mixed mullerian tumour|8950/3
C0206627|T191|SY|0000020977|CHV|mullerian mixed tumor|8950/3
C0206627|T191|SY|0000020977|CHV|mullerian mixed tumour|8950/3
C0206627|T191|PT|271538|MEDCIN|Mullerian mixed tumor|8950/3
C0206627|T191|MH|D018200|MSH|Mixed Tumor, Mullerian|8950/3
C0206627|T191|PM|D018200|MSH|Mullerian Mixed Tumor|8950/3
C0206627|T191|PM|D018200|MSH|Tumor, Mullerian Mixed|8950/3
C0206627|T191|PN|NOCODE|MTH|Mixed Tumor, Mullerian|8950/3
C0206627|T191|SY|C3730|NCI|Mixed Müllerian Tumor|8950/3
C0206627|T191|PT|CDR0000335077|NCI_NCI-GLOSS|Mullerian tumor|8950/3
C0206627|T191|PT|BBL5.|RCD|Mullerian mixed tumour|8950/3
C0206627|T191|PT|BBL5.|RCDAE|Mullerian mixed tumor|8950/3
C0206627|T191|SY|84427001|SNOMEDCT_US|Malignant mixed mesodermal tumor|8950/3
C0206627|T191|SYGB|84427001|SNOMEDCT_US|Malignant mixed mesodermal tumour|8950/3
C0206627|T191|SY|84427001|SNOMEDCT_US|Malignant mixed Mullerian tumor|8950/3
C0206627|T191|SYGB|84427001|SNOMEDCT_US|Malignant mixed Mullerian tumour|8950/3
C0206627|T191|PT|84427001|SNOMEDCT_US|Mullerian mixed tumor|8950/3
C0206627|T191|PTGB|84427001|SNOMEDCT_US|Mullerian mixed tumour|8950/3
C0206627|T191|PT|0046136|CCPSS|MULLERIAN MIXED TUMOR|8951/3
C1334603|T191|PT|0000020976|CHV|mesodermal mixed tumor|8951/3
C1334603|T191|SY|0000020976|CHV|mixed mesodermal tumor|8951/3
C1334603|T191|SY|0000020976|CHV|mixed mesodermal tumors|8951/3
C0206627|T191|PT|0000020977|CHV|mixed mullerian tumor|8951/3
C0206627|T191|SY|0000020977|CHV|mixed mullerian tumors|8951/3
C0206627|T191|SY|0000020977|CHV|mixed mullerian tumour|8951/3
C0206627|T191|SY|0000020977|CHV|mullerian mixed tumor|8951/3
C0206627|T191|SY|0000020977|CHV|mullerian mixed tumour|8951/3
C1334603|T191|PT|271539|MEDCIN|mesodermal mixed tumor|8951/3
C0206627|T191|PT|271538|MEDCIN|Mullerian mixed tumor|8951/3
C1334603|T191|PM|D018199|MSH|Mesodermal Mixed Tumor|8951/3
C1334603|T191|PM|D018199|MSH|Mesodermal Mixed Tumors|8951/3
C1334603|T191|MH|D018199|MSH|Mixed Tumor, Mesodermal|8951/3
C0206627|T191|MH|D018200|MSH|Mixed Tumor, Mullerian|8951/3
C1334603|T191|PM|D018199|MSH|Mixed Tumors, Mesodermal|8951/3
C0206627|T191|PM|D018200|MSH|Mullerian Mixed Tumor|8951/3
C1334603|T191|PM|D018199|MSH|Tumor, Mesodermal Mixed|8951/3
C0206627|T191|PM|D018200|MSH|Tumor, Mullerian Mixed|8951/3
C1334603|T191|PM|D018199|MSH|Tumors, Mesodermal Mixed|8951/3
C0206627|T191|PN|NOCODE|MTH|Mixed Tumor, Mullerian|8951/3
C1334603|T191|SY|C8975|NCI|Malignant Mixed Mesodermal Tumor|8951/3
C1334603|T191|SY|C8975|NCI|Malignant Mixed Mullerian Tumor|8951/3
C0206627|T191|SY|C3730|NCI|Mixed Müllerian Tumor|8951/3
C1334603|T191|AB|C8975|NCI|MMMT|8951/3
C1334603|T191|SY|C8975|NCI_CDISC|Malignant Mixed Mesodermal Tumor|8951/3
C1334603|T191|SY|C8975|NCI_CDISC|MMMT|8951/3
C1334603|T191|PT|C8975|NCI_CDISC|MULLERIAN TUMOR, MIXED, MALIGNANT|8951/3
C1334603|T191|PT|CDR0000335078|NCI_NCI-GLOSS|malignant mixed Mullerian tumor|8951/3
C1334603|T191|SY|CDR0000533838|NCI_NCI-GLOSS|MMMT|8951/3
C0206627|T191|PT|CDR0000335077|NCI_NCI-GLOSS|Mullerian tumor|8951/3
C1334603|T191|PT|BBL6.|RCD|Mesodermal mixed tumour|8951/3
C0206627|T191|PT|BBL5.|RCD|Mullerian mixed tumour|8951/3
C1334603|T191|PT|BBL6.|RCDAE|Mesodermal mixed tumor|8951/3
C0206627|T191|PT|BBL5.|RCDAE|Mullerian mixed tumor|8951/3
C0206627|T191|SY|84427001|SNOMEDCT_US|Malignant mixed mesodermal tumor|8951/3
C1334603|T191|OAS|112684005|SNOMEDCT_US|Malignant mixed mesodermal tumor|8951/3
C1334603|T191|OAS|112684005|SNOMEDCT_US|Malignant mixed mesodermal tumour|8951/3
C0206627|T191|SYGB|84427001|SNOMEDCT_US|Malignant mixed mesodermal tumour|8951/3
C0206627|T191|SY|84427001|SNOMEDCT_US|Malignant mixed Mullerian tumor|8951/3
C0206627|T191|SYGB|84427001|SNOMEDCT_US|Malignant mixed Mullerian tumour|8951/3
C1334603|T191|OAP|112684005|SNOMEDCT_US|Mesodermal mixed tumor|8951/3
C1334603|T191|OAP|112684005|SNOMEDCT_US|Mesodermal mixed tumour|8951/3
C0206627|T191|PT|84427001|SNOMEDCT_US|Mullerian mixed tumor|8951/3
C0206627|T191|PTGB|84427001|SNOMEDCT_US|Mullerian mixed tumour|8951/3
C1266138|T191|PT|C7504|NCI|Adult Cystic Nephroma|8959/0
C1266138|T191|DN|C7504|NCI_CTRP|Cystic Nephroma|8959/0
C1266138|T191|SY|CDR0000582682|PDQ|Benign Cystic Nephroma|8959/0
C1266138|T191|PT|CDR0000582682|PDQ|cystic nephroma|8959/0
C1266138|T191|PT|128757006|SNOMEDCT_US|Benign cystic nephroma|8959/0
C1266139|T191|SY|234226|MEDCIN|malignant cystic nephroma|8959/1
C1266139|T191|PT|234226|MEDCIN|malignant cystic nephroma of kidney|8959/1
C1266139|T191|PN|NOCODE|MTH|Cystic Partially Differentiated Nephroblastoma|8959/1
C1266139|T191|PT|C6897|NCI|Cystic Partially Differentiated Kidney Nephroblastoma|8959/1
C1266139|T191|SY|C6897|NCI|Malignant Cystic Nephroma|8959/1
C1266139|T191|SY|C6897|NCI|Malignant Multilocular Cystic Nephroma|8959/1
C1266139|T191|PT|C6897|NCI_NICHD|Cystic Partially Differentiated Nephroblastoma|8959/1
C1266139|T191|PT|128758001|SNOMEDCT_US|Cystic partially differentiated nephroblastoma|8959/1
C1266139|T191|PT|128759009|SNOMEDCT_US|Malignant cystic nephroma|8959/1
C1266139|T191|SY|128759009|SNOMEDCT_US|Malignant multilocular cystic nephroma|8959/1
C1266139|T191|SY|234226|MEDCIN|malignant cystic nephroma|8959/3
C1266139|T191|PT|234226|MEDCIN|malignant cystic nephroma of kidney|8959/3
C1266139|T191|PN|NOCODE|MTH|Cystic Partially Differentiated Nephroblastoma|8959/3
C1266139|T191|PT|C6897|NCI|Cystic Partially Differentiated Kidney Nephroblastoma|8959/3
C1266139|T191|SY|C6897|NCI|Malignant Cystic Nephroma|8959/3
C1266139|T191|SY|C6897|NCI|Malignant Multilocular Cystic Nephroma|8959/3
C1266139|T191|PT|C6897|NCI_NICHD|Cystic Partially Differentiated Nephroblastoma|8959/3
C1266139|T191|PT|128758001|SNOMEDCT_US|Cystic partially differentiated nephroblastoma|8959/3
C1266139|T191|PT|128759009|SNOMEDCT_US|Malignant cystic nephroma|8959/3
C1266139|T191|SY|128759009|SNOMEDCT_US|Malignant multilocular cystic nephroma|8959/3
C0206628|T191|PT|0000020978|CHV|mesoblastic nephroma|8960/1
C1332965|T191|PT|HP:0100881|HPO|Congenital mesoblastic nephroma|8960/1
C0206628|T191|PT|MTHU048909|ICPC2ICD10ENG|mesoblastic; nephroma|8960/1
C0206628|T191|PT|MTHU052070|ICPC2ICD10ENG|nephroma; mesoblastic|8960/1
C0206628|T191|PT|10070665|MDR|Mesoblastic nephroma|8960/1
C0206628|T191|LLT|10070665|MDR|Mesoblastic nephroma|8960/1
C0206628|T191|PT|351906|MEDCIN|Mesoblastic nephroma|8960/1
C1332965|T191|DEV|D018201|MSH|CONGEN MESOBLASTIC NEPHROMA|8960/1
C1332965|T191|PEP|D018201|MSH|Congenital Mesoblastic Nephroma|8960/1
C1332965|T191|PM|D018201|MSH|Congenital Mesoblastic Nephromas|8960/1
C0206628|T191|ET|D018201|MSH|Mesoblastic Nephroma|8960/1
C1332965|T191|PM|D018201|MSH|Mesoblastic Nephroma, Congenital|8960/1
C1332965|T191|PM|D018201|MSH|Mesoblastic Nephromas, Congenital|8960/1
C1332965|T191|PM|D018201|MSH|Nephroma, Congenital Mesoblastic|8960/1
C0206628|T191|MH|D018201|MSH|Nephroma, Mesoblastic|8960/1
C1332965|T191|PM|D018201|MSH|Nephromas, Congenital Mesoblastic|8960/1
C0206628|T191|PM|D018201|MSH|Nephromas, Mesoblastic|8960/1
C1332965|T191|PN|NOCODE|MTH|Congenital Mesoblastic Nephroma|8960/1
C0206628|T191|PN|NOCODE|MTH|Mesoblastic Nephroma|8960/1
C1332965|T191|AB|C6569|NCI|CMN|8960/1
C1332965|T191|PT|C6569|NCI|Congenital Mesoblastic Nephroma|8960/1
C1332965|T191|SY|C6569|NCI|Mesoblastic Nephroma|8960/1
C1332965|T191|SY|C6569|NCI_CDISC|CMN|8960/1
C1332965|T191|PT|C6569|NCI_CDISC|STROMAL NEPHROMA, MALIGNANT|8960/1
C1332965|T191|DN|C6569|NCI_CTRP|Congenital Mesoblastic Nephroma|8960/1
C1332965|T191|PT|CDR0000534218|NCI_NCI-GLOSS|congenital mesoblastic nephroma|8960/1
C1332965|T191|PT|C6569|NCI_NICHD|Congenital Mesoblastic Nephroma|8960/1
C1332965|T191|AB|CDR0000566112|PDQ|CMN|8960/1
C1332965|T191|PT|CDR0000566112|PDQ|congenital mesoblastic nephroma|8960/1
C1332965|T191|SY|CDR0000566112|PDQ|Mesoblastic Nephroma|8960/1
C0206628|T191|PT|XaBAx|RCD|Mesoblastic nephroma|8960/1
C0206628|T191|PT|BBL70|RCDSY|Mesoblastic nephroma|8960/1
C0206628|T191|PT|307604008|SNOMEDCT_US|Mesoblastic nephroma|8960/1
C0206628|T191|PT|11793003|SNOMEDCT_US|Mesoblastic nephroma|8960/1
C1320471|T191|PT|405941007|SNOMEDCT_US|Mesoblastic nephroma, cellular|8960/1
C1320470|T191|PT|405940008|SNOMEDCT_US|Mesoblastic nephroma, classical|8960/1
C1320472|T191|PT|405942000|SNOMEDCT_US|Mesoblastic nephroma, mixed|8960/1
C0027708|T191|ET|0000004550|AOD|nephroblastoma|8960/3
C0027708|T191|NP|0000023021|AOD|Wilms tumor|8960/3
C0027708|T191|PT|0048278|CCPSS|WILMS TUMOR|8960/3
C0027708|T191|SY|0000008581|CHV|nephroblastoma|8960/3
C0027708|T191|SY|0000008581|CHV|nephroma|8960/3
C0027708|T191|SY|0000008581|CHV|nephromas|8960/3
C0027708|T191|SY|0000008581|CHV|tumor wilm's|8960/3
C0027708|T191|SY|0000008581|CHV|tumor wilms|8960/3
C0027708|T191|SY|0000008581|CHV|tumor wilms'|8960/3
C0027708|T191|SY|0000008581|CHV|tumor wilms's|8960/3
C0027708|T191|SY|0000008581|CHV|tumors wilm's|8960/3
C0027708|T191|SY|0000008581|CHV|tumors wilms|8960/3
C0027708|T191|SY|0000008581|CHV|wilm tumor|8960/3
C0027708|T191|SY|0000008581|CHV|wilm's tumor|8960/3
C0027708|T191|PT|0000008581|CHV|wilms tumor|8960/3
C0027708|T191|SY|0000008581|CHV|wilms tumour|8960/3
C0027708|T191|SY|0000008581|CHV|wilms' tumor|8960/3
C0027708|T191|SY|0000008581|CHV|wilms' tumour|8960/3
C0027708|T191|PT|NOCODE|COSTAR|Wilm's Tumor|8960/3
C0027708|T191|PT|2021-2990|CSP|nephroblastoma|8960/3
C0027708|T191|PT|4001-0143|CSP|Wilms' tumor|8960/3
C0027708|T191|GT|CARCINOMA|CST|WILMS TUMOR|8960/3
C0027708|T191|SY|NOCODE|DXP|KIDNEY, ADENOMYOSARCOMA, EMBRYONAL|8960/3
C0027708|T191|SY|NOCODE|DXP|KIDNEY, CARCINOSARCOMA, EMBRYONAL|8960/3
C0027708|T191|SY|NOCODE|DXP|KIDNEY, EMBRYOMA|8960/3
C0027708|T191|SY|NOCODE|DXP|KIDNEY, EMBRYONAL MIXED TUMOR|8960/3
C0027708|T191|SY|NOCODE|DXP|NEPHROBLASTOMA|8960/3
C0027708|T191|SY|NOCODE|DXP|RENAL CANCER, WILMS|8960/3
C0027708|T191|DI|U002025|DXP|WILMS TUMOR|8960/3
C0027708|T191|PT|HP:0002667|HPO|Nephroblastoma|8960/3
C0027708|T191|SY|HP:0002667|HPO|Wilm's tumor|8960/3
C0027708|T191|SY|HP:0002667|HPO|Wilms tumor|8960/3
C0027708|T191|PT|MTHU025491|ICPC2ICD10ENG|embryoma; kidney|8960/3
C0027708|T191|PT|MTHU052990|ICPC2ICD10ENG|kidney; embryoma|8960/3
C0027708|T191|PT|MTHU052063|ICPC2ICD10ENG|nephroblastoma|8960/3
C0027708|T191|PT|MTHU052069|ICPC2ICD10ENG|nephroma|8960/3
C0027708|T191|PT|MTHU077184|ICPC2ICD10ENG|tumor; Wilms|8960/3
C0027708|T191|PT|MTHU082457|ICPC2ICD10ENG|Wilms|8960/3
C0027708|T191|PT|MTHU082458|ICPC2ICD10ENG|Wilms; tumor|8960/3
C0027708|T191|PT|sh85090858|LCH_NW|Nephroblastoma|8960/3
C0027708|T191|PT|10029145|MDR|Nephroblastoma|8960/3
C0027708|T191|LLT|10029145|MDR|Nephroblastoma|8960/3
C0027708|T191|LLT|10047985|MDR|Wilms tumor|8960/3
C0027708|T191|LLT|10047986|MDR|Wilms tumour|8960/3
C0027708|T191|LLT|10047987|MDR|Wilms' tumor|8960/3
C0027708|T191|SY|31531|MEDCIN|nephroblastoma|8960/3
C0027708|T191|PT|31531|MEDCIN|nephroblastoma of kidney|8960/3
C0027708|T191|SY|3075|MEDLINEPLUS|Nephroblastoma|8960/3
C0027708|T191|ET|3075|MEDLINEPLUS|Nephroblastoma|8960/3
C0027708|T191|PT|3075|MEDLINEPLUS|Wilms Tumor|8960/3
C0027708|T191|ET|D009396|MSH|Nephroblastoma|8960/3
C0027708|T191|PM|D009396|MSH|Nephroblastomas|8960/3
C0027708|T191|PM|D009396|MSH|Tumor, Wilms|8960/3
C0027708|T191|PM|D009396|MSH|Tumor, Wilms'|8960/3
C0027708|T191|PM|D009396|MSH|Wilm Tumor|8960/3
C0027708|T191|PM|D009396|MSH|Wilm's Tumor|8960/3
C0027708|T191|MH|D009396|MSH|Wilms Tumor|8960/3
C0027708|T191|ET|D009396|MSH|Wilms Tumor 1|8960/3
C0027708|T191|ET|D009396|MSH|Wilms' Tumor|8960/3
C0027708|T191|PN|NOCODE|MTH|Nephroblastoma|8960/3
C0027708|T191|SY|C40407|NCI|Kidney Nephroblastoma|8960/3
C0027708|T191|PT|C40407|NCI|Kidney Wilms Tumor|8960/3
C0027708|T191|SY|C3267|NCI|Nephroblastoma|8960/3
C0027708|T191|SY|C40407|NCI|Renal Wilms Tumor|8960/3
C0027708|T191|SY|C40407|NCI|Renal Wilms' Tumor|8960/3
C0027708|T191|PT|C3267|NCI|Wilms Tumor|8960/3
C0027708|T191|SY|C40407|NCI|Wilms Tumor of the Kidney|8960/3
C0027708|T191|SY|C3267|NCI|Wilms' Tumor|8960/3
C0027708|T191|SY|C40407|NCI|Wilms' Tumor of the Kidney|8960/3
C0027708|T191|SY|C40407|NCI_CDISC|Embryonal Nephroma|8960/3
C0027708|T191|SY|C40407|NCI_CDISC|Nephroblastoma|8960/3
C0027708|T191|PT|C40407|NCI_CDISC|NEPHROBLASTOMA, MALIGNANT|8960/3
C0027708|T191|SY|C40407|NCI_CDISC|Renal Wilms' Tumor|8960/3
C0027708|T191|SY|C40407|NCI_CDISC|Wilms Tumor of the Kidney|8960/3
C0027708|T191|SY|C40407|NCI_CDISC|Wilms' Tumor of the Kidney|8960/3
C0027708|T191|PT|C3267|NCI_CPTAC|Wilms Tumor|8960/3
C0027708|T191|DN|C3267|NCI_CTRP|Wilms Tumor|8960/3
C0027708|T191|PT|C3267|NCI_CTRP|Wilms Tumor|8960/3
C0027708|T191|PT|CDR0000045946|NCI_NCI-GLOSS|Wilms' tumor|8960/3
C0027708|T191|PT|C40407|NCI_NICHD|Nephroblastoma|8960/3
C0027708|T191|PT|C3267|NCI_NICHD|Wilms Tumor|8960/3
C0027708|T191|SY|CDR0000042957|PDQ|nephroblastoma|8960/3
C0027708|T191|SY|CDR0000042957|PDQ|tumor, Wilms'|8960/3
C0027708|T191|SY|CDR0000042957|PDQ|Wilm's tumor|8960/3
C0027708|T191|SY|CDR0000042957|PDQ|Wilms tumor|8960/3
C0027708|T191|ET|CDR0000042957|PDQ|Wilms tumor|8960/3
C0027708|T191|PSC|CDR0000042957|PDQ|Wilms tumor and other childhood kidney tumors|8960/3
C0027708|T191|SY|CDR0000042957|PDQ|Wilms' tumor and other childhood kidney tumors|8960/3
C0027708|T191|PT|Xa9A0|RCD|Nephroblastoma|8960/3
C0027708|T191|SY|Xa9A0|RCD|Nephroma|8960/3
C0027708|T191|SY|Xa9A0|RCD|Wilms' tumour|8960/3
C0027708|T191|SY|Xa9A0|RCDAE|Wilms' tumor|8960/3
C0027708|T191|SY|BBLE.|RCDSY|Nephroblastoma NOS|8960/3
C0027708|T191|SY|25081006|SNOMEDCT_US|Embryonal adenosarcoma|8960/3
C0027708|T191|SY|25081006|SNOMEDCT_US|Embryonal nephroma|8960/3
C0027708|T191|PT|25081006|SNOMEDCT_US|Nephroblastoma|8960/3
C0027708|T191|PT|302849000|SNOMEDCT_US|Nephroblastoma|8960/3
C1319302|T191|PT|405939006|SNOMEDCT_US|Nephroblastoma, diffuse anaplasia|8960/3
C1319300|T191|PT|405937008|SNOMEDCT_US|Nephroblastoma, favorable histology|8960/3
C1319300|T191|PTGB|405937008|SNOMEDCT_US|Nephroblastoma, favourable histology|8960/3
C1319301|T191|PT|405938003|SNOMEDCT_US|Nephroblastoma, focal anaplasia|8960/3
C0027708|T191|IS|25081006|SNOMEDCT_US|Nephroblastoma, NOS|8960/3
C0027708|T191|SY|302849000|SNOMEDCT_US|Nephroma|8960/3
C0027708|T191|SY|25081006|SNOMEDCT_US|Nephroma|8960/3
C0027708|T191|IS|25081006|SNOMEDCT_US|Nephroma, NOS|8960/3
C0027708|T191|IS|302849000|SNOMEDCT_US|Perlman syndrome|8960/3
C0027708|T191|SY|25081006|SNOMEDCT_US|Renal adenosarcoma|8960/3
C0027708|T191|SY|302849000|SNOMEDCT_US|Wilm's tumor|8960/3
C0027708|T191|SY|302849000|SNOMEDCT_US|Wilms tumor|8960/3
C0027708|T191|SYGB|302849000|SNOMEDCT_US|Wilms tumour|8960/3
C0027708|T191|SY|25081006|SNOMEDCT_US|Wilms' tumor|8960/3
C0027708|T191|IS|302849000|SNOMEDCT_US|Wilms' tumor|8960/3
C1319302|T191|SY|405939006|SNOMEDCT_US|Wilms' tumor, diffuse anaplasia|8960/3
C1319300|T191|SY|405937008|SNOMEDCT_US|Wilms' tumor, favorable histology|8960/3
C1319301|T191|SY|405938003|SNOMEDCT_US|Wilms' tumor, focal anaplasia|8960/3
C0027708|T191|IS|302849000|SNOMEDCT_US|Wilms' tumour|8960/3
C0027708|T191|SYGB|25081006|SNOMEDCT_US|Wilms' tumour|8960/3
C1319302|T191|SYGB|405939006|SNOMEDCT_US|Wilms' tumour, diffuse anaplasia|8960/3
C1319300|T191|SYGB|405937008|SNOMEDCT_US|Wilms' tumour, favourable histology|8960/3
C1319301|T191|SYGB|405938003|SNOMEDCT_US|Wilms' tumour, focal anaplasia|8960/3
C0206743|T191|SY|0000021063|CHV|malignant rhabdoid tumor|8963/3
C0206743|T191|SY|0000021063|CHV|rhabdoid sarcoma|8963/3
C0206743|T191|PT|0000021063|CHV|rhabdoid tumor|8963/3
C0206743|T191|SY|0000021063|CHV|rhabdoid tumors|8963/3
C0206743|T191|SY|0000021063|CHV|sarcoma rhabdoid|8963/3
C0206743|T191|MTH_PT|10073334|MDR|Rhabdoid tumor|8963/3
C0206743|T191|LLT|10073335|MDR|Rhabdoid tumor|8963/3
C0206743|T191|LLT|10073334|MDR|Rhabdoid tumour|8963/3
C0206743|T191|PT|10073334|MDR|Rhabdoid tumour|8963/3
C0206743|T191|MH|D018335|MSH|Rhabdoid Tumor|8963/3
C0206743|T191|PM|D018335|MSH|Rhabdoid Tumors|8963/3
C0206743|T191|PM|D018335|MSH|Tumor, Rhabdoid|8963/3
C0206743|T191|PM|D018335|MSH|Tumors, Rhabdoid|8963/3
C0206743|T191|PN|NOCODE|MTH|Rhabdoid Tumor|8963/3
C0206743|T191|OP|C3808|NCI|Rhabdoid Sarcoma|8963/3
C0206743|T191|PT|C3808|NCI|Rhabdoid Tumor|8963/3
C0206743|T191|PT|CDR0000046139|NCI_NCI-GLOSS|rhabdoid tumor|8963/3
C0206743|T191|PT|C3808|NCI_NICHD|Rhabdoid Tumor|8963/3
C0206743|T191|PT|X77ol|RCD|Rhabdoid sarcoma|8963/3
C0206743|T191|PT|83118000|SNOMEDCT_US|Malignant rhabdoid tumor|8963/3
C0206743|T191|PTGB|83118000|SNOMEDCT_US|Malignant rhabdoid tumour|8963/3
C0206743|T191|OAP|189812005|SNOMEDCT_US|Rhabdoid sarcoma|8963/3
C0206743|T191|OF|189812005|SNOMEDCT_US|Rhabdoid sarcoma|8963/3
C0206743|T191|SY|83118000|SNOMEDCT_US|Rhabdoid sarcoma|8963/3
C0206743|T191|SY|83118000|SNOMEDCT_US|Rhabdoid tumor|8963/3
C0206743|T191|SYGB|83118000|SNOMEDCT_US|Rhabdoid tumour|8963/3
C0334488|T191|SY|0000029995|CHV|clear cell sarcoma kidney|8964/3
C0334488|T191|PT|0000029995|CHV|clear cell sarcoma of the kidney|8964/3
C0334488|T191|PT|MTHU016917|ICPC2ICD10ENG|clear cell; sarcoma, kidney|8964/3
C0334488|T191|PT|MTHU052961|ICPC2ICD10ENG|kidney; clear cell sarcoma|8964/3
C0334488|T191|PT|MTHU053092|ICPC2ICD10ENG|kidney; sarcoma, clear cell|8964/3
C0334488|T191|PT|MTHU065893|ICPC2ICD10ENG|sarcoma; clear cell, kidney|8964/3
C0334488|T191|LLT|10009253|MDR|Clear cell sarcoma of the kidney|8964/3
C0334488|T191|PT|10009253|MDR|Clear cell sarcoma of the kidney|8964/3
C0334488|T191|PT|234210|MEDCIN|clear cell sarcoma of kidney|8964/3
C0334488|T191|PN|NOCODE|MTH|Clear cell sarcoma of kidney|8964/3
C0334488|T191|AB|C4264|NCI|CCSK|8964/3
C0334488|T191|SY|C4264|NCI|Childhood Clear Cell Sarcoma of the Kidney|8964/3
C0334488|T191|SY|C4264|NCI|Childhood Kidney Clear Cell Sarcoma|8964/3
C0334488|T191|SY|C4264|NCI|Childhood Renal Clear Cell Sarcoma|8964/3
C0334488|T191|SY|C4264|NCI|Clear Cell Sarcoma of Kidney|8964/3
C0334488|T191|PT|C4264|NCI|Clear Cell Sarcoma of the Kidney|8964/3
C0334488|T191|SY|C4264|NCI|Kidney Clear Cell Sarcoma|8964/3
C0334488|T191|SY|C4264|NCI|Pediatric Kidney Clear Cell Sarcoma|8964/3
C0334488|T191|SY|C4264|NCI|Pediatric Renal Clear Cell Sarcoma|8964/3
C0334488|T191|SY|C4264|NCI|Renal Clear Cell Sarcoma|8964/3
C0334488|T191|SY|10009253|NCI_CTEP-SDC|Clear cell sarcoma - kidney|8964/3
C0334488|T191|PT|10009253|NCI_CTEP-SDC|Clear cell sarcoma of the kidney|8964/3
C0334488|T191|DN|C4264|NCI_CTRP|Clear Cell Sarcoma of the Kidney|8964/3
C0334488|T191|PT|CDR0000044997|NCI_NCI-GLOSS|clear cell sarcoma of the kidney|8964/3
C0334488|T191|PT|C4264|NCI_NICHD|Clear Cell Sarcoma of the Kidney|8964/3
C0334488|T191|AB|CDR0000038146|PDQ|CCSK|8964/3
C0334488|T191|SY|CDR0000038146|PDQ|Childhood Clear Cell Sarcoma of the Kidney|8964/3
C0334488|T191|SY|CDR0000038146|PDQ|Childhood Kidney Clear Cell Sarcoma|8964/3
C0334488|T191|SY|CDR0000038146|PDQ|Childhood Renal Clear Cell Sarcoma|8964/3
C0334488|T191|SY|CDR0000038146|PDQ|Clear Cell Sarcoma of Kidney|8964/3
C0334488|T191|PT|CDR0000038146|PDQ|clear cell sarcoma of the kidney|8964/3
C0334488|T191|SY|CDR0000038146|PDQ|kidney clear cell sarcoma|8964/3
C0334488|T191|SY|CDR0000038146|PDQ|Pediatric Kidney Clear Cell Sarcoma|8964/3
C0334488|T191|SY|CDR0000038146|PDQ|Pediatric Renal Clear Cell Sarcoma|8964/3
C0334488|T191|SY|CDR0000038146|PDQ|Renal Clear Cell Sarcoma|8964/3
C0334488|T191|PT|X77om|RCD|Clear cell sarcoma of kidney|8964/3
C0334488|T191|OP|BBLJ.|RCDSY|Clear cell sarcoma of kidney|8964/3
C0334488|T191|OA|BBLJ.|RCDSY|Clear cell sarcoma,kidney|8964/3
C0334488|T191|PT|24007003|SNOMEDCT_US|Clear cell sarcoma of kidney|8964/3
C1266141|T191|PT|C39812|NCI|Metanephric Adenofibroma|8965/0
C1266141|T191|SY|C39812|NCI|Nephrogenic Adenofibroma|8965/0
C1266141|T191|SY|128760004|SNOMEDCT_US|Metanephric adenofibroma|8965/0
C1266141|T191|PT|128760004|SNOMEDCT_US|Nephrogenic adenofibroma|8965/0
C1266142|T191|PT|HP:0008696|HPO|Renal hamartoma|8966/0
C1266142|T191|SY|C5100|NCI|Fibroma of Renal Medulla|8966/0
C1266142|T191|SY|C5100|NCI|Kidney Fibroma|8966/0
C1266142|T191|SY|C5100|NCI|Medullary Fibroma|8966/0
C1266142|T191|SY|C5100|NCI|Renal Hamartoma|8966/0
C1266142|T191|PT|C5100|NCI|Renomedullary Interstitial Cell Tumor|8966/0
C1266142|T191|SY|128761000|SNOMEDCT_US|Renomedullary fibroma|8966/0
C1266142|T191|PT|128761000|SNOMEDCT_US|Renomedullary interstitial cell tumor|8966/0
C1266142|T191|PTGB|128761000|SNOMEDCT_US|Renomedullary interstitial cell tumour|8966/0
C1882198|T191|AB|C66774|NCI|ORTI|8967/0
C1882198|T191|PT|C66774|NCI|Ossifying Renal Tumor of Infancy|8967/0
C1266143|T191|PT|128762007|SNOMEDCT_US|Ossifying renal tumor|8967/0
C1266143|T191|PTGB|128762007|SNOMEDCT_US|Ossifying renal tumour|8967/0
C0206624|T191|PT|0000020975|CHV|hepatoblastoma|8970/3
C0206624|T191|PT|4003-0022|CSP|hepatoblastoma|8970/3
C0206624|T191|DI|U000819|DXP|HEPATOBLASTOMA|8970/3
C0206624|T191|PT|HP:0002884|HPO|Hepatoblastoma|8970/3
C0206624|T191|PT|C22.2|ICD10|Hepatoblastoma|8970/3
C0206624|T191|AB|C22.2|ICD10CM|Hepatoblastoma|8970/3
C0206624|T191|PT|C22.2|ICD10CM|Hepatoblastoma|8970/3
C0206624|T191|PT|MTHU025478|ICPC2ICD10ENG|embryonal; hepatoma|8970/3
C0206624|T191|PT|MTHU034359|ICPC2ICD10ENG|hepatoblastoma|8970/3
C0206624|T191|PT|MTHU034386|ICPC2ICD10ENG|hepatoma; embryonal|8970/3
C0206624|T191|PT|10062001|MDR|Hepatoblastoma|8970/3
C0206624|T191|LLT|10062001|MDR|Hepatoblastoma|8970/3
C0206624|T191|LLT|10019822|MDR|Hepatoblastoma NOS|8970/3
C0206624|T191|HT|10019825|MDR|Hepatoblastomas|8970/3
C0206624|T191|SY|36086|MEDCIN|hepatoblastoma|8970/3
C0206624|T191|PT|36086|MEDCIN|hepatoblastoma of liver|8970/3
C0206624|T191|ET|309|MEDLINEPLUS|Hepatoblastoma|8970/3
C0206624|T191|MH|D018197|MSH|Hepatoblastoma|8970/3
C0206624|T191|PM|D018197|MSH|Hepatoblastomas|8970/3
C0206624|T191|PN|NOCODE|MTH|Hepatoblastoma|8970/3
C0206624|T191|ET|155.0|MTHICD9|Hepatoblastoma|8970/3
C0206624|T191|AB|C3728|NCI|HBL|8970/3
C0206624|T191|PT|C3728|NCI|Hepatoblastoma|8970/3
C1333982|T191|PT|C7093|NCI|Hepatoblastoma with Pure Fetal Epithelial Differentiation|8970/3
C1334784|T191|PT|C7097|NCI|Mixed Epithelial and Mesenchymal Hepatoblastoma|8970/3
C0206624|T191|SY|C3728|NCI|Pediatric Embryonal Hepatoma|8970/3
C0206624|T191|SY|C3728|NCI|Pediatric Hepatoblastoma|8970/3
C0206624|T191|SY|C3728|NCI_CDISC|HBL|8970/3
C0206624|T191|PT|C3728|NCI_CDISC|HEPATOBLASTOMA, MALIGNANT|8970/3
C0206624|T191|SY|C3728|NCI_CDISC|Pediatric Embryonal Hepatoma|8970/3
C0206624|T191|SY|C3728|NCI_CDISC|Pediatric Hepatoblastoma|8970/3
C0206624|T191|PT|C3728|NCI_CPTAC|Hepatoblastoma|8970/3
C0206624|T191|PT|10019822|NCI_CTEP-SDC|Hepatoblastoma|8970/3
C0206624|T191|PT|C3728|NCI_CTRP|Hepatoblastoma|8970/3
C0206624|T191|DN|C3728|NCI_CTRP|Hepatoblastoma|8970/3
C0206624|T191|PT|CDR0000046160|NCI_NCI-GLOSS|hepatoblastoma|8970/3
C0206624|T191|PT|C3728|NCI_NICHD|Hepatoblastoma|8970/3
C1333982|T191|PT|C7093|NCI_NICHD|Hepatoblastoma with Pure Fetal Epithelial Differentiation|8970/3
C1334784|T191|PT|C7097|NCI_NICHD|Mixed Epithelial and Mesenchymal Hepatoblastoma|8970/3
C0206624|T191|PT|CDR0000043722|PDQ|childhood hepatoblastoma|8970/3
C0206624|T191|AB|CDR0000043722|PDQ|HBL|8970/3
C0206624|T191|SY|CDR0000043722|PDQ|Hepatoblastoma|8970/3
C0206624|T191|SY|CDR0000043722|PDQ|hepatoblastoma, childhood|8970/3
C0206624|T191|SY|CDR0000043722|PDQ|Pediatric Embryonal Hepatoma|8970/3
C0206624|T191|SY|CDR0000043722|PDQ|pediatric hepatoblastoma|8970/3
C0206624|T191|SY|BBL8.|RCD|Embryonal hepatoma|8970/3
C0206624|T191|SY|BBL8.|RCD|HBL - Hepatoblastoma|8970/3
C0206624|T191|PT|BBL8.|RCD|Hepatoblastoma|8970/3
C0206624|T191|PT|B1501|RCD|Hepatoblastoma of liver|8970/3
C0206624|T191|SY|45024009|SNOMEDCT_US|Embryonal hepatoma|8970/3
C4518346|T191|PT|734035004|SNOMEDCT_US|Epithelial variant hepatoblastoma|8970/3
C0206624|T191|SY|45024009|SNOMEDCT_US|HBL - Hepatoblastoma|8970/3
C0206624|T191|PT|109843000|SNOMEDCT_US|Hepatoblastoma|8970/3
C0206624|T191|PT|45024009|SNOMEDCT_US|Hepatoblastoma|8970/3
C0206624|T191|SY|109843000|SNOMEDCT_US|Hepatoblastoma of liver|8970/3
C4518346|T191|SY|734035004|SNOMEDCT_US|Hepatoblastoma, epithelial variant|8970/3
C1334784|T191|SY|734033006|SNOMEDCT_US|Hepatoblastoma, mixed epithelial-mesenchymal|8970/3
C1334784|T191|PT|734033006|SNOMEDCT_US|Mixed epithelial-mesenchymal hepatoblastoma|8970/3
C0334489|T191|PT|0000029996|CHV|pancreatoblastoma|8971/3
C0334489|T191|PT|HP:0100757|HPO|Pancreatoblastoma|8971/3
C0334489|T191|LLT|10073367|MDR|Pancreatoblastoma|8971/3
C0334489|T191|PT|10073367|MDR|Pancreatoblastoma|8971/3
C0334489|T191|PT|38726|MEDCIN|pancreatoblastoma|8971/3
C0334489|T191|NM|C537162|MSH|Pancreatoblastoma|8971/3
C0334489|T191|PT|C4265|NCI|Pancreatoblastoma|8971/3
C0334489|T191|PT|X77on|RCD|Pancreatoblastoma|8971/3
C0334489|T191|PT|53618008|SNOMEDCT_US|Pancreatoblastoma|8971/3
C0334489|T191|OAP|189814006|SNOMEDCT_US|Pancreatoblastoma|8971/3
C0334489|T191|OF|189814006|SNOMEDCT_US|Pancreatoblastoma|8971/3
C0206629|T191|PT|0004173|CCPSS|PULMONARY BLASTOMA|8972/3
C0206629|T191|SY|0000020979|CHV|pneumoblastoma|8972/3
C0206629|T191|PT|0000020979|CHV|pulmonary blastoma|8972/3
C0206629|T191|DEV|D018202|MSH|BLASTOMA PULM|8972/3
C0206629|T191|ET|D018202|MSH|Blastoma, Pulmonary|8972/3
C0206629|T191|DEV|D018202|MSH|BLASTOMAS PULM|8972/3
C0206629|T191|ET|D018202|MSH|Blastomas, Pulmonary|8972/3
C0206629|T191|DEV|D018202|MSH|PULM BLASTOMA|8972/3
C0206629|T191|DEV|D018202|MSH|PULM BLASTOMAS|8972/3
C0206629|T191|MH|D018202|MSH|Pulmonary Blastoma|8972/3
C0206629|T191|ET|D018202|MSH|Pulmonary Blastomas|8972/3
C0206629|T191|SY|C3732|NCI|Blastoma of Lung|8972/3
C0206629|T191|SY|C3732|NCI|Blastoma of the Lung|8972/3
C0206629|T191|SY|C3732|NCI|Lung Blastoma|8972/3
C0206629|T191|SY|C3732|NCI|Pneumoblastoma|8972/3
C0206629|T191|PT|C3732|NCI|Pulmonary Blastoma|8972/3
C0206629|T191|SY|X77oo|RCD|Pneumoblastoma|8972/3
C0206629|T191|PT|X77oo|RCD|Pulmonary blastoma|8972/3
C0206629|T191|SY|43149009|SNOMEDCT_US|Pneumoblastoma|8972/3
C0206629|T191|PT|189815007|SNOMEDCT_US|Pulmonary blastoma|8972/3
C0206629|T191|PT|43149009|SNOMEDCT_US|Pulmonary blastoma|8972/3
C0206629|T191|OF|189815007|SNOMEDCT_US|Pulmonary blastoma|8972/3
C1266144|T191|PT|HP:0100528|HPO|Pleuropulmonary blastoma|8973/3
C1266144|T191|PT|10080682|MDR|Pleuropulmonary blastoma|8973/3
C1266144|T191|LLT|10080682|MDR|Pleuropulmonary blastoma|8973/3
C1266144|T191|NM|C537516|MSH|Pleuropulmonary blastoma|8973/3
C1266144|T191|PN|NOCODE|MTH|Pleuropulmonary blastoma|8973/3
C1266144|T191|PT|C5669|NCI|Pleuropulmonary Blastoma|8973/3
C1266144|T191|SY|C5669|NCI|Pulmonary Blastoma of Childhood|8973/3
C1266144|T191|PT|C5669|NCI_CPTAC|Pleuropulmonary Blastoma|8973/3
C1266144|T191|PT|C5669|NCI_CTRP|Pleuropulmonary Blastoma|8973/3
C1266144|T191|DN|C5669|NCI_CTRP|Pleuropulmonary Blastoma|8973/3
C1266144|T191|PT|CDR0000446557|NCI_NCI-GLOSS|pleuropulmonary blastoma|8973/3
C1266144|T191|PT|C5669|NCI_NICHD|Pleuropulmonary Blastoma|8973/3
C1266144|T191|PT|CDR0000582828|PDQ|pleuropulmonary blastoma|8973/3
C1266144|T191|SY|CDR0000582828|PDQ|Pulmonary Blastoma of Childhood|8973/3
C1266144|T191|SY|707670009|SNOMEDCT_US|Pleuro-pulmonary blastoma|8973/3
C1266144|T191|PT|707670009|SNOMEDCT_US|Pleuropulmonary blastoma|8973/3
C1266144|T191|PT|128763002|SNOMEDCT_US|Pleuropulmonary blastoma|8973/3
C1335911|T191|PT|C35837|NCI|Salivary Gland Sialoblastoma|8974/1
C1266145|T191|PT|128764008|SNOMEDCT_US|Sialoblastoma|8974/1
C3273067|T191|PT|C96830|NCI|Calcifying Nested Epithelial Stromal Tumor of the Liver|8975/1
C3472610|T191|PT|450898007|SNOMEDCT_US|Calcifying nested epithelial stromal tumor|8975/1
C3472610|T191|PTGB|450898007|SNOMEDCT_US|Calcifying nested epithelial stromal tumour|8975/1
C0007140|T191|PT|0000002439|CHV|carcinosarcoma|8980/3
C0007140|T191|SY|0000002439|CHV|carcinosarcomas|8980/3
C0007140|T191|PT|2000-3358|CSP|carcinosarcoma|8980/3
C0007140|T191|PT|271530|MEDCIN|carcinosarcoma|8980/3
C0007140|T191|MH|D002296|MSH|Carcinosarcoma|8980/3
C0007140|T191|PM|D002296|MSH|Carcinosarcomas|8980/3
C0007140|T191|PN|NOCODE|MTH|Carcinosarcoma|8980/3
C0007140|T191|PT|C34448|NCI|Carcinosarcoma|8980/3
C0007140|T191|PT|C34448|NCI_CDISC|CARCINOSARCOMA, MALIGNANT|8980/3
C0007140|T191|PT|C34448|NCI_CTRP|Carcinosarcoma|8980/3
C0007140|T191|DN|C34448|NCI_CTRP|Carcinosarcoma|8980/3
C0007140|T191|PT|CDR0000044003|NCI_NCI-GLOSS|carcinosarcoma|8980/3
C0007140|T191|PT|Xa9A1|RCD|Carcinosarcoma|8980/3
C0007140|T191|OP|BBL9.|RCDSY|Carcinosarcoma NOS|8980/3
C0007140|T191|PT|63264007|SNOMEDCT_US|Carcinosarcoma|8980/3
C0007140|T191|IS|63264007|SNOMEDCT_US|Carcinosarcoma, NOS|8980/3
C0334490|T191|PT|271531|MEDCIN|embryonal carcinosarcoma|8981/3
C0936282|T191|PT|C8997|NCI|Blastoma|8981/3
C0936282|T191|SY|C8997|NCI|Embryoma|8981/3
C0936282|T191|PT|CDR0000367443|NCI_NCI-GLOSS|embryoma|8981/3
C0936282|T191|SY|BB02.|RCD|Blastoma|8981/3
C0334490|T191|PT|BBLA.|RCD|Embryonal carcinosarcoma,|8981/3
C0936282|T191|SY|86049000|SNOMEDCT_US|Blastoma|8981/3
C0936282|T191|IS|86049000|SNOMEDCT_US|Blastoma, NOS|8981/3
C0334490|T191|PT|112685006|SNOMEDCT_US|Carcinosarcoma, embryonal|8981/3
C0334490|T191|SY|112685006|SNOMEDCT_US|Embryonal carcinosarcoma|8981/3
C0334490|T191|IS|112685006|SNOMEDCT_US|Embryonal carcinosarcoma,|8981/3
C0027070|T191|SY|0000008429|CHV|myoepithelial tumor|8982/0
C0027070|T191|PT|0000008429|CHV|myoepithelioma|8982/0
C0027070|T191|ET|D009208|MSH|Myoepithelial Tumor|8982/0
C0027070|T191|PM|D009208|MSH|Myoepithelial Tumors|8982/0
C0027070|T191|MH|D009208|MSH|Myoepithelioma|8982/0
C0027070|T191|PM|D009208|MSH|Myoepitheliomas|8982/0
C0027070|T191|PM|D009208|MSH|Tumor, Myoepithelial|8982/0
C0027070|T191|PM|D009208|MSH|Tumors, Myoepithelial|8982/0
C0027070|T191|PN|NOCODE|MTH|Myoepithelioma|8982/0
C0027070|T191|SY|C40392|NCI|Myoepithelial Neoplasm|8982/0
C0027070|T191|PT|C40392|NCI|Myoepithelial Tumor|8982/0
C0027070|T191|SY|C40392|NCI|Myoepithelioma|8982/0
C0027070|T191|SY|BBLB.|RCD|Myoepithelial tumour|8982/0
C0027070|T191|PT|BBLB.|RCD|Myoepithelioma|8982/0
C0027070|T191|SY|BBLB.|RCDAE|Myoepithelial tumor|8982/0
C0027070|T191|SY|69291002|SNOMEDCT_US|Myoepithelial adenoma|8982/0
C0027070|T191|SY|69291002|SNOMEDCT_US|Myoepithelial tumor|8982/0
C0027070|T191|SYGB|69291002|SNOMEDCT_US|Myoepithelial tumour|8982/0
C0027070|T191|PT|69291002|SNOMEDCT_US|Myoepithelioma|8982/0
C0027070|T191|SY|0000008429|CHV|myoepithelial tumor|8982/1
C0027070|T191|PT|0000008429|CHV|myoepithelioma|8982/1
C0027070|T191|ET|D009208|MSH|Myoepithelial Tumor|8982/1
C0027070|T191|PM|D009208|MSH|Myoepithelial Tumors|8982/1
C0027070|T191|MH|D009208|MSH|Myoepithelioma|8982/1
C0027070|T191|PM|D009208|MSH|Myoepitheliomas|8982/1
C0027070|T191|PM|D009208|MSH|Tumor, Myoepithelial|8982/1
C0027070|T191|PM|D009208|MSH|Tumors, Myoepithelial|8982/1
C0027070|T191|PN|NOCODE|MTH|Myoepithelioma|8982/1
C0027070|T191|SY|C40392|NCI|Myoepithelial Neoplasm|8982/1
C0027070|T191|PT|C40392|NCI|Myoepithelial Tumor|8982/1
C0027070|T191|SY|C40392|NCI|Myoepithelioma|8982/1
C0027070|T191|SY|BBLB.|RCD|Myoepithelial tumour|8982/1
C0027070|T191|PT|BBLB.|RCD|Myoepithelioma|8982/1
C0027070|T191|SY|BBLB.|RCDAE|Myoepithelial tumor|8982/1
C0027070|T191|SY|69291002|SNOMEDCT_US|Myoepithelial adenoma|8982/1
C0027070|T191|SY|69291002|SNOMEDCT_US|Myoepithelial tumor|8982/1
C0027070|T191|SYGB|69291002|SNOMEDCT_US|Myoepithelial tumour|8982/1
C0027070|T191|PT|69291002|SNOMEDCT_US|Myoepithelioma|8982/1
C0334699|T191|PT|0000030023|CHV|myoepithelial carcinoma|8982/3
C0334699|T191|PT|271532|MEDCIN|malignant myoepithelioma|8982/3
C0334699|T191|PN|NOCODE|MTH|Malignant myoepithelioma|8982/3
C0334699|T191|PT|C7596|NCI|Malignant Myoepithelioma|8982/3
C0334699|T191|SY|C7596|NCI|Myoepithelial Carcinoma|8982/3
C0334699|T191|SY|C7596|NCI_CDISC|Malignant Myoepithelioma|8982/3
C0334699|T191|SY|C7596|NCI_CDISC|Myoepithelial Carcinoma|8982/3
C0334699|T191|PT|C7596|NCI_CDISC|MYOEPITHELIOMA, MALIGNANT|8982/3
C0334699|T191|PT|C7596|NCI_CPTAC|Malignant Myoepithelioma|8982/3
C0334699|T191|PT|CDR0000778443|PDQ|malignant myoepithelioma|8982/3
C0334699|T191|SY|CDR0000778443|PDQ|myoepithelial carcinoma|8982/3
C0334699|T191|SY|128884000|SNOMEDCT_US|Infiltrating myoepithelioma|8982/3
C0334699|T191|OAP|24292006|SNOMEDCT_US|Malignant myoepithelioma|8982/3
C0334699|T191|PT|128884000|SNOMEDCT_US|Malignant myoepithelioma|8982/3
C0334699|T191|IS|24292006|SNOMEDCT_US|Malignant myoepithelioma -RETIRED-|8982/3
C0334699|T191|OF|24292006|SNOMEDCT_US|Malignant myoepithelioma -RETIRED-|8982/3
C0334699|T191|SY|128884000|SNOMEDCT_US|Myoepithelial carcinoma|8982/3
C1266146|T191|MH|D055331|MSH|Adenomyoepithelioma|8983/0
C1266146|T191|PM|D055331|MSH|Adenomyoepitheliomas|8983/0
C1266146|T191|PN|NOCODE|MTH|Adenomyoepithelioma|8983/0
C1510795|T191|SY|C6899|NCI|Adenomyoepithelioma of the Breast|8983/0
C1510795|T191|PT|C6899|NCI|Breast Adenomyoepithelioma|8983/0
C1266146|T191|PT|C124607|NCI|Experimental Organism Benign Adenomyoepithelioma|8983/0
C1266146|T191|PT|C124607|NCI_CDISC|ADENOMYOEPITHELIOMA, BENIGN|8983/0
C1266146|T191|PT|128765009|SNOMEDCT_US|Adenomyoepithelioma|8983/0
C1266146|T191|SY|128765009|SNOMEDCT_US|Adenomyoepithelioma, benign|8983/0
C3839546|T191|PT|703644009|SNOMEDCT_US|Adenomyoepithelioma with carcinoma|8983/3
C3839546|T191|SY|703644009|SNOMEDCT_US|Malignant adenomyoepithelioma|8983/3
C3814879|T191|MTH_PT|10079470|MDR|Phosphaturic mesenchymal tumor|8990/0
C3814879|T191|LLT|10079478|MDR|Phosphaturic mesenchymal tumor|8990/0
C3814879|T191|LLT|10079470|MDR|Phosphaturic mesenchymal tumour|8990/0
C3814879|T191|PT|10079470|MDR|Phosphaturic mesenchymal tumour|8990/0
C0334491|T191|PN|NOCODE|MTH|Benign Mesenchymoma|8990/0
C3814879|T191|PN|NOCODE|MTH|Phosphaturic mesenchymal tumor, benign|8990/0
C0334491|T191|OP|C4267|NCI|Benign Mesenchymoma|8990/0
C0334491|T191|PT|C4267|NCI|Benign Mesenchymoma|8990/0
C3814879|T191|PT|C121788|NCI|Benign Phosphaturic Mesenchymal Tumor|8990/0
C0334491|T191|PT|C4267|NCI_CDISC|MESENCHYMAL TUMOR, BENIGN|8990/0
C0334491|T191|PT|BBLC0|RCD|Benign mesenchymoma|8990/0
C0334491|T191|SY|38406003|SNOMEDCT_US|Benign mesenchymoma|8990/0
C0334491|T191|PT|38406003|SNOMEDCT_US|Mesenchymoma, benign|8990/0
C3814879|T191|SY|703649004|SNOMEDCT_US|Phosphaturic mesenchymal tumor|8990/0
C3814879|T191|PT|703649004|SNOMEDCT_US|Phosphaturic mesenchymal tumor, benign|8990/0
C3814879|T191|SYGB|703649004|SNOMEDCT_US|Phosphaturic mesenchymal tumour|8990/0
C3814879|T191|PTGB|703649004|SNOMEDCT_US|Phosphaturic mesenchymal tumour, benign|8990/0
C0025464|T191|ET|0000004537|AOD|mesenchymoma|8990/1
C0025464|T191|PT|0000007982|CHV|mesenchymoma|8990/1
C1300127|T191|PT|0000057615|CHV|pecoma|8990/1
C1300127|T191|SY|0000057615|CHV|pecomas|8990/1
C0025464|T191|PT|2000-4749|CSP|mesenchymoma|8990/1
C0025464|T191|MH|D008637|MSH|Mesenchymoma|8990/1
C0025464|T191|PM|D008637|MSH|Mesenchymomas|8990/1
C1300127|T191|ET|D054973|MSH|Neoplasms, Perivascular Epithelioid Cell|8990/1
C1300127|T191|PM|D054973|MSH|PEComa|8990/1
C1300127|T191|ET|D054973|MSH|PEComas|8990/1
C1300127|T191|MH|D054973|MSH|Perivascular Epithelioid Cell Neoplasms|8990/1
C1300127|T191|ET|D054973|MSH|Perivascular Epithelioid Cell Tumors|8990/1
C0025464|T191|OP|C3233|NCI|Mesenchymoma|8990/1
C0025464|T191|PT|C3233|NCI|Mesenchymoma|8990/1
C1300127|T191|SY|C38150|NCI|Neoplasm with Perivascular Epithelioid Cell Differentiation|8990/1
C1300127|T191|PT|C38150|NCI|PEComa|8990/1
C1300127|T191|SY|C38150|NCI|Tumor with Perivascular Epithelioid Cell Differentiation|8990/1
C1300127|T191|SY|CDR0000778387|PDQ|neoplasm with perivascular epithelioid cell differentiation|8990/1
C1300127|T191|PT|CDR0000778387|PDQ|PEComa|8990/1
C1300127|T191|SY|CDR0000778387|PDQ|tumor with perivascular epithelioid cell differentiation|8990/1
C0025464|T191|SY|BBLC.|RCD|Mesenchymoma|8990/1
C0025464|T191|SY|BBLC.|RCD|Mixed mesenchymal tumour|8990/1
C0025464|T191|SY|BBLC.|RCDAE|Mixed mesenchymal tumor|8990/1
C0025464|T191|OP|BBLCz|RCDSY|Mesenchymoma NOS|8990/1
C0025464|T191|PT|BBLC.|RCDSY|Mesenchymomas|8990/1
C0025464|T191|PT|44524009|SNOMEDCT_US|Mesenchymoma|8990/1
C0025464|T191|IS|44524009|SNOMEDCT_US|Mesenchymoma, NOS|8990/1
C0025464|T191|SY|44524009|SNOMEDCT_US|Mesenchymomas|8990/1
C0025464|T191|SY|44524009|SNOMEDCT_US|Mixed mesenchymal tumor|8990/1
C0025464|T191|SYGB|44524009|SNOMEDCT_US|Mixed mesenchymal tumour|8990/1
C1300127|T191|SY|388601000|SNOMEDCT_US|PEComa|8990/1
C1300127|T191|SY|388601000|SNOMEDCT_US|Perivascular epithelial cell tumor|8990/1
C1300127|T191|SYGB|388601000|SNOMEDCT_US|Perivascular epithelial cell tumour|8990/1
C1300127|T191|PT|388601000|SNOMEDCT_US|Perivascular epithelioid cell tumor|8990/1
C1300127|T191|PTGB|388601000|SNOMEDCT_US|Perivascular epithelioid cell tumour|8990/1
C5230988|T191|PT|817951007|SNOMEDCT_US|Primitive non-neural granular cell tumor|8990/1
C5230988|T191|PTGB|817951007|SNOMEDCT_US|Primitive non-neural granular cell tumour|8990/1
C0334492|T191|PT|0000029997|CHV|malignant mesenchymoma|8990/3
C0334492|T191|SY|0000029997|CHV|malignant mesenchymomas|8990/3
C0334492|T191|LLT|10061526|MDR|Malignant mesenchymoma|8990/3
C0334492|T191|PT|10061526|MDR|Malignant mesenchymoma|8990/3
C0334492|T191|LLT|10025676|MDR|Malignant mesenchymoma NOS|8990/3
C0334492|T191|LLT|10025678|MDR|Malignant mesenchymoma stage unspecified|8990/3
C0334492|T191|HT|10025673|MDR|Mesenchymomas malignant|8990/3
C0334492|T191|PT|271540|MEDCIN|malignant mesenchymoma|8990/3
C0334492|T191|NM|C535700|MSH|Malignant mesenchymal tumor|8990/3
C0334492|T191|CE|C535700|MSH|Malignant mesenchymoma|8990/3
C0334492|T191|PN|NOCODE|MTH|Malignant mesenchymal tumor|8990/3
C0334492|T191|OP|C4268|NCI|Malignant Mesenchymoma|8990/3
C0334492|T191|PT|C4268|NCI|Malignant Mesenchymoma|8990/3
C3839061|T191|PT|C121789|NCI|Malignant Phosphaturic Mesenchymal Tumor|8990/3
C0334492|T191|PT|C4268|NCI_CDISC|MESENCHYMOMA, MALIGNANT|8990/3
C0334492|T191|PT|BBLC1|RCD|Malignant mesenchymoma|8990/3
C0334492|T191|SY|BBLC1|RCD|Mixed mesenchymal sarcoma|8990/3
C0334492|T191|SY|89623007|SNOMEDCT_US|Malignant mesenchymoma|8990/3
C0334492|T191|PT|89623007|SNOMEDCT_US|Mesenchymoma, malignant|8990/3
C0334492|T191|SY|89623007|SNOMEDCT_US|Mixed mesenchymal sarcoma|8990/3
C3839061|T191|PT|703650004|SNOMEDCT_US|Phosphaturic mesenchymal tumor, malignant|8990/3
C3839061|T191|PTGB|703650004|SNOMEDCT_US|Phosphaturic mesenchymal tumour, malignant|8990/3
C0855073|T191|PT|0000050298|CHV|undifferentiated sarcoma|8991/3
C0855073|T191|PT|MTHU025481|ICPC2ICD10ENG|embryonal; sarcoma|8991/3
C0855073|T191|PT|MTHU065894|ICPC2ICD10ENG|sarcoma; embryonal|8991/3
C0855073|T191|LLT|10045515|MDR|Undifferentiated sarcoma|8991/3
C0855073|T191|PT|10045515|MDR|Undifferentiated sarcoma|8991/3
C0855073|T191|PT|271500|MEDCIN|embryonal sarcoma|8991/3
C0855073|T191|PT|271497|MEDCIN|undifferentiated sarcoma|8991/3
C0855073|T191|SY|C27096|NCI|Embryonal Sarcoma|8991/3
C0855073|T191|AB|C27096|NCI|UES|8991/3
C0855073|T191|SY|C27096|NCI|Undifferentiated Sarcoma|8991/3
C0855073|T191|SY|C27096|NCI_CDISC|Embryonal Sarcoma, Undifferentiated|8991/3
C0855073|T191|PT|C27096|NCI_CDISC|SARCOMA, UNDIFFERENTIATED, MALIGNANT|8991/3
C0855073|T191|PT|BBLD.|RCD|Embryonal sarcoma|8991/3
C0855073|T191|PT|59583009|SNOMEDCT_US|Embryonal sarcoma|8991/3
C0855073|T191|PT|128734000|SNOMEDCT_US|Undifferentiated sarcoma|8991/3
C0006160|T191|PT|0021673|CCPSS|BRENNER TUMOR|9000/0
C0006160|T191|PT|0000002163|CHV|brenner tumor|9000/0
C0006160|T191|SY|0000002163|CHV|brenner tumors|9000/0
C0006160|T191|SY|0000002163|CHV|brenner tumour|9000/0
C0006160|T191|SY|NOCODE|DXP|OVARIAN CANCER, BRENNER|9000/0
C0006160|T191|DI|U001366|DXP|OVARY, BRENNER TUMOR|9000/0
C0006160|T191|SY|NOCODE|DXP|OVARY, FIBROEPITHELIOMA|9000/0
C0006160|T191|PT|MTHU012689|ICPC2ICD10ENG|Brenner; tumor|9000/0
C0006160|T191|PT|MTHU077029|ICPC2ICD10ENG|tumor; Brenner|9000/0
C0006160|T191|LLT|10073271|MDR|Brenner tumor|9000/0
C0006160|T191|MTH_PT|10073258|MDR|Brenner tumor|9000/0
C0006160|T191|LLT|10073258|MDR|Brenner tumour|9000/0
C0006160|T191|PT|10073258|MDR|Brenner tumour|9000/0
C0474834|T191|PT|34922|MEDCIN|benign Brenner tumor of ovary|9000/0
C0474834|T191|PEP|D001948|MSH|Benign Brenner Tumor|9000/0
C0006160|T191|MH|D001948|MSH|Brenner Tumor|9000/0
C0006160|T191|ET|D001948|MSH|Brenner Tumor of Ovary|9000/0
C0474834|T191|PM|D001948|MSH|Brenner Tumor, Benign|9000/0
C0006160|T191|ET|D001948|MSH|Ovarian Brenner Tumor|9000/0
C0006160|T191|PM|D001948|MSH|Ovary Brenner Tumor|9000/0
C0006160|T191|PN|NOCODE|MTH|Brenner Tumor|9000/0
C4551593|T191|PN|NOCODE|MTH|Surface epithelial-stromal tumor|9000/0
C0474834|T191|SY|C4746|NCI|Benign Brenner Neoplasm of Ovary|9000/0
C0474834|T191|SY|C4746|NCI|Benign Brenner Neoplasm of the Ovary|9000/0
C0474834|T191|SY|C4746|NCI|Benign Brenner Tumor of Ovary|9000/0
C0474834|T191|SY|C4746|NCI|Benign Brenner Tumor of the Ovary|9000/0
C0474834|T191|SY|C4746|NCI|Benign Ovarian Brenner Neoplasm|9000/0
C0474834|T191|PT|C4746|NCI|Benign Ovarian Brenner Tumor|9000/0
C0006160|T191|SY|C3872|NCI|Brenner Neoplasm of Ovary|9000/0
C0006160|T191|SY|C3872|NCI|Brenner Neoplasm of the Ovary|9000/0
C0006160|T191|SY|C3872|NCI|Brenner Tumor|9000/0
C0006160|T191|PT|C39954|NCI|Brenner Tumor|9000/0
C0006160|T191|SY|C3872|NCI|Brenner Tumor of Ovary|9000/0
C0006160|T191|SY|C3872|NCI|Brenner Tumor of the Ovary|9000/0
C0006160|T191|SY|C3872|NCI|Ovarian Brenner Neoplasm|9000/0
C0006160|T191|PT|C3872|NCI|Ovarian Brenner Tumor|9000/0
C0006160|T191|DN|C3872|NCI_CTRP|Ovarian Brenner Tumor|9000/0
C0006160|T191|SY|CDR0000043342|PDQ|Brenner neoplasm of ovary|9000/0
C0006160|T191|SY|CDR0000043342|PDQ|Brenner neoplasm of the ovary|9000/0
C0006160|T191|PT|CDR0000043342|PDQ|Brenner tumor|9000/0
C0006160|T191|SY|CDR0000043342|PDQ|Brenner tumor of ovary|9000/0
C0006160|T191|SY|CDR0000043342|PDQ|Brenner tumor of the ovary|9000/0
C0006160|T191|SY|CDR0000043342|PDQ|ovarian Brenner neoplasm|9000/0
C0006160|T191|SY|CDR0000043342|PDQ|ovarian Brenner tumor|9000/0
C0474834|T191|PT|X77os|RCD|Benign Brenner tumour|9000/0
C4551593|T191|PT|XM1FP|RCD|Brenner tumour|9000/0
C0006160|T191|PT|X78Ww|RCD|Brenner tumour of ovary|9000/0
C0474834|T191|PT|X77os|RCDAE|Benign Brenner tumor|9000/0
C4551593|T191|PT|XM1FP|RCDAE|Brenner tumor|9000/0
C0006160|T191|PT|X78Ww|RCDAE|Brenner tumor of ovary|9000/0
C0006160|T191|OP|BBM0z|RCDSA|Brenner tumor NOS|9000/0
C0006160|T191|OP|BBM0.|RCDSA|Brenner tumors|9000/0
C0006160|T191|OP|BBM0z|RCDSY|Brenner tumour NOS|9000/0
C0006160|T191|OP|BBM0.|RCDSY|Brenner tumours|9000/0
C0474834|T191|PT|253051001|SNOMEDCT_US|Benign Brenner tumor|9000/0
C0474834|T191|PTGB|253051001|SNOMEDCT_US|Benign Brenner tumour|9000/0
C4551593|T191|PT|768795009|SNOMEDCT_US|Brenner tumor|9000/0
C0006160|T191|OAP|74739000|SNOMEDCT_US|Brenner tumor|9000/0
C0006160|T191|PT|254859006|SNOMEDCT_US|Brenner tumor of ovary|9000/0
C0006160|T191|IS|74739000|SNOMEDCT_US|Brenner tumor, NOS|9000/0
C0006160|T191|OAP|74739000|SNOMEDCT_US|Brenner tumour|9000/0
C4551593|T191|PTGB|768795009|SNOMEDCT_US|Brenner tumour|9000/0
C0006160|T191|PTGB|254859006|SNOMEDCT_US|Brenner tumour of ovary|9000/0
C4551593|T191|SY|768795009|SNOMEDCT_US|Surface epithelial-stromal tumor|9000/0
C4551593|T191|SYGB|768795009|SNOMEDCT_US|Surface epithelial-stromal tumour|9000/0
C0334494|T191|PT|MTHU012111|ICPC2ICD10ENG|borderline malignancy; Brenner tumor|9000/1
C0334494|T191|PT|MTHU012690|ICPC2ICD10ENG|Brenner; tumor, borderline malignancy|9000/1
C0334494|T191|PT|MTHU012692|ICPC2ICD10ENG|Brenner; tumor, proliferating|9000/1
C0334494|T191|PT|MTHU062032|ICPC2ICD10ENG|proliferating; Brenner tumor|9000/1
C0334494|T191|PT|MTHU077030|ICPC2ICD10ENG|tumor; Brenner, borderline malignancy|9000/1
C0334494|T191|PT|MTHU077032|ICPC2ICD10ENG|tumor; Brenner, proliferating|9000/1
C0334494|T191|PN|NOCODE|MTH|Proliferating Brenner Tumor|9000/1
C0334494|T191|SY|C9459|NCI|Borderline Brenner Neoplasm of Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Borderline Brenner Neoplasm of the Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Borderline Brenner Tumor of Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Borderline Brenner Tumor of the Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Borderline Ovarian Brenner Neoplasm|9000/1
C0334494|T191|SY|C9459|NCI|Borderline Ovarian Brenner Tumor|9000/1
C0334494|T191|PT|C9459|NCI|Borderline Ovarian Brenner Tumor/Atypical Proliferative Ovarian Brenner Tumor|9000/1
C0334494|T191|SY|C9459|NCI|Low Malignancy Potential Brenner Neoplasm of Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Low Malignancy Potential Brenner Neoplasm of the Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Low Malignancy Potential Brenner Tumor of Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Low Malignancy Potential Brenner Tumor of the Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Low Malignancy Potential Ovarian Brenner Neoplasm|9000/1
C0334494|T191|SY|C9459|NCI|Low Malignancy Potential Ovarian Brenner Tumor|9000/1
C0334494|T191|SY|C9459|NCI|Proliferating Brenner Neoplasm of Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Proliferating Brenner Neoplasm of the Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Proliferating Brenner Tumor of Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Proliferating Brenner Tumor of the Ovary|9000/1
C0334494|T191|SY|C9459|NCI|Proliferating Ovarian Brenner Neoplasm|9000/1
C0334494|T191|SY|C9459|NCI|Proliferating Ovarian Brenner Tumor|9000/1
C0334494|T191|AB|BBM00|RCD|Brenner tumour - border malign|9000/1
C0334494|T191|PT|BBM00|RCD|Brenner tumour - borderline malignancy|9000/1
C0334494|T191|SY|BBM00|RCD|Proliferating Brenner tumour|9000/1
C0334494|T191|AB|BBM00|RCDAE|Brenner tumor - border malign|9000/1
C0334494|T191|PT|BBM00|RCDAE|Brenner tumor - borderline malignancy|9000/1
C0334494|T191|SY|BBM00|RCDAE|Proliferating Brenner tumor|9000/1
C0334494|T191|SY|89996007|SNOMEDCT_US|Borderline Brenner tumor|9000/1
C0334494|T191|SYGB|89996007|SNOMEDCT_US|Borderline Brenner tumour|9000/1
C0334494|T191|SY|89996007|SNOMEDCT_US|Brenner tumor - borderline malignancy|9000/1
C0334494|T191|SY|89996007|SNOMEDCT_US|Brenner tumor, atypical proliferative|9000/1
C0334494|T191|PT|89996007|SNOMEDCT_US|Brenner tumor, borderline malignancy|9000/1
C0334494|T191|SY|89996007|SNOMEDCT_US|Brenner tumor, proliferating|9000/1
C0334494|T191|SYGB|89996007|SNOMEDCT_US|Brenner tumour - borderline malignancy|9000/1
C0334494|T191|SYGB|89996007|SNOMEDCT_US|Brenner tumour, atypical proliferative|9000/1
C0334494|T191|PTGB|89996007|SNOMEDCT_US|Brenner tumour, borderline malignancy|9000/1
C0334494|T191|SYGB|89996007|SNOMEDCT_US|Brenner tumour, proliferating|9000/1
C0334494|T191|SY|89996007|SNOMEDCT_US|Proliferating Brenner tumor|9000/1
C0334494|T191|SYGB|89996007|SNOMEDCT_US|Proliferating Brenner tumour|9000/1
C0334495|T191|PT|MTHU012691|ICPC2ICD10ENG|Brenner; tumor, malignant|9000/3
C0334495|T191|PT|MTHU077031|ICPC2ICD10ENG|tumor; Brenner, malignant|9000/3
C0334495|T191|PT|34899|MEDCIN|malignant Brenner tumor of ovary|9000/3
C0334495|T191|PM|D001948|MSH|Brenner Tumor, Malignant|9000/3
C0334495|T191|PEP|D001948|MSH|Malignant Brenner Tumor|9000/3
C0334495|T191|SY|C4270|NCI|Malignant Brenner Tumor of Ovary|9000/3
C0334495|T191|SY|C4270|NCI|Malignant Brenner Tumor of the Ovary|9000/3
C0334495|T191|PT|C4270|NCI|Malignant Ovarian Brenner Tumor|9000/3
C0334495|T191|DN|C4270|NCI_CTRP|Malignant Ovarian Brenner Tumor|9000/3
C0334495|T191|PT|BBM01|RCD|Malignant Brenner tumour|9000/3
C0334495|T191|PT|BBM01|RCDAE|Malignant Brenner tumor|9000/3
C0334495|T191|PT|42194009|SNOMEDCT_US|Brenner tumor, malignant|9000/3
C0334495|T191|PTGB|42194009|SNOMEDCT_US|Brenner tumour, malignant|9000/3
C0334495|T191|SY|42194009|SNOMEDCT_US|Malignant Brenner tumor|9000/3
C0334495|T191|SYGB|42194009|SNOMEDCT_US|Malignant Brenner tumour|9000/3
C0178421|T191|SY|0000018289|CHV|adenofibroma breast|9010/0
C0178421|T191|PT|0000018289|CHV|breast fibroadenoma|9010/0
C0178421|T191|SY|0000018289|CHV|breast fibroadenomas|9010/0
C0178421|T191|SY|0000018289|CHV|breast mouse|9010/0
C0206650|T191|PT|0000020995|CHV|fibroadenoma|9010/0
C0178421|T191|SY|0000018289|CHV|fibroadenoma breast|9010/0
C0178421|T191|SY|0000018289|CHV|fibroadenoma of breast|9010/0
C0206650|T191|SY|0000020995|CHV|fibroadenomas|9010/0
C0178421|T191|PT|U000289|COSTAR|FIBROADENOMA OF BREAST|9010/0
C0178421|T191|SY|NOCODE|DXP|BREAST, ADENOFIBROMA|9010/0
C0178421|T191|DI|U000247|DXP|BREAST, FIBROADENOMA|9010/0
C0178421|T191|SY|HP:0010619|HPO|Breast fibroadenoma|9010/0
C0178421|T191|SY|HP:0010619|HPO|Breast fibroadenomas|9010/0
C0178421|T191|PT|HP:0010619|HPO|Fibroadenoma of the breast|9010/0
C0178421|T191|ET|D24|ICD10CM|fibroadenoma of breast|9010/0
C0206650|T191|PT|MTHU028164|ICPC2ICD10ENG|fibroadenoma; unspecified site|9010/0
C0178421|T191|LLT|10006276|MDR|Breast mouse|9010/0
C0206650|T191|LLT|10063384|MDR|Fibroadenoma|9010/0
C0178421|T191|LLT|10016613|MDR|Fibroadenoma of breast|9010/0
C0178421|T191|PT|10016613|MDR|Fibroadenoma of breast|9010/0
C0178421|T191|PT|31650|MEDCIN|fibroadenoma of breast|9010/0
C0206650|T191|MH|D018226|MSH|Fibroadenoma|9010/0
C0206650|T191|PM|D018226|MSH|Fibroadenomas|9010/0
C0206650|T191|PN|NOCODE|MTH|Fibroadenoma|9010/0
C0178421|T191|PN|NOCODE|MTH|Fibroadenoma of breast|9010/0
C0178421|T191|PT|C3744|NCI|Breast Fibroadenoma|9010/0
C0178421|T191|SY|C3744|NCI|Fibroadenoma|9010/0
C0178421|T191|SY|C3744|NCI|Fibroadenoma of Breast|9010/0
C0178421|T191|SY|C3744|NCI|Fibroadenoma of the Breast|9010/0
C0178421|T191|SY|C3744|NCI_CDISC|Breast Fibroadenoma|9010/0
C0178421|T191|SY|C3744|NCI_CDISC|Fibroadenoma of Breast|9010/0
C0178421|T191|SY|C3744|NCI_CDISC|Fibroadenoma of the Breast|9010/0
C0178421|T191|PT|C3744|NCI_CDISC|FIBROADENOMA, BENIGN|9010/0
C0178421|T191|PT|CDR0000523438|NCI_NCI-GLOSS|fibroadenoma|9010/0
C0178421|T191|SY|X78WY|RCD|Breast mouse|9010/0
C0206650|T191|PT|Xa9A3|RCD|Fibroadenoma|9010/0
C0178421|T191|PT|X78WY|RCD|Fibroadenoma of breast|9010/0
C0206650|T191|OP|BBM1.|RCDSY|Fibroadenoma NOS|9010/0
C0178421|T191|OAS|269640007|SNOMEDCT_US|Breast fibroadenoma|9010/0
C0178421|T191|SY|254845004|SNOMEDCT_US|Breast mouse|9010/0
C0206650|T191|PT|65877006|SNOMEDCT_US|Fibroadenoma|9010/0
C0178421|T191|OAS|269640007|SNOMEDCT_US|Fibroadenoma of breast|9010/0
C0178421|T191|OAS|189102001|SNOMEDCT_US|Fibroadenoma of breast|9010/0
C0178421|T191|PT|254845004|SNOMEDCT_US|Fibroadenoma of breast|9010/0
C0206650|T191|SY|65877006|SNOMEDCT_US|Fibroadenoma, no ICD-O subtype|9010/0
C0206650|T191|SY|65877006|SNOMEDCT_US|Fibroadenoma, no International Classification of Diseases for Oncology subtype|9010/0
C0206650|T191|IS|65877006|SNOMEDCT_US|Fibroadenoma, NOS|9010/0
C0334496|T191|SY|NOCODE|DXP|BREAST, FIBROADENOMA, INTRACANALICULAR|9011/0
C0334496|T191|PT|C4271|NCI|Breast Intracanalicular Fibroadenoma|9011/0
C0334496|T191|SY|C4271|NCI|Intracanalicular Breast Fibroadenoma|9011/0
C0334496|T191|SY|C4271|NCI|Intracanalicular Fibroadenoma|9011/0
C0334496|T191|SY|C4271|NCI|Intracanalicular Fibroadenoma of Breast|9011/0
C0334496|T191|SY|C4271|NCI|Intracanalicular Fibroadenoma of the Breast|9011/0
C0334496|T191|PT|Xa9A4|RCD|Intracanalicular fibroadenoma|9011/0
C0334496|T191|OA|BBM2.|RCDSY|Intracanal.fibroadenoma NOS|9011/0
C0334496|T191|OP|BBM2.|RCDSY|Intracanalicular fibroadenoma NOS|9011/0
C0334496|T191|PT|72905006|SNOMEDCT_US|Intracanalicular fibroadenoma|9011/0
C0334496|T191|IS|72905006|SNOMEDCT_US|Intracanalicular fibroadenoma, NOS|9011/0
C0334497|T191|PT|MTHU028165|ICPC2ICD10ENG|fibroadenoma; pericanalicular, unspecified site|9012/0
C0334497|T191|PT|MTHU058604|ICPC2ICD10ENG|pericanalicular; fibroadenoma, unspecified site|9012/0
C0334497|T191|PT|C4272|NCI|Breast Pericanalicular Fibroadenoma|9012/0
C0334497|T191|SY|C4272|NCI|Pericanalicular Breast Fibroadenoma|9012/0
C0334497|T191|SY|C4272|NCI|Pericanalicular Fibroadenoma|9012/0
C0334497|T191|SY|C4272|NCI|Pericanalicular Fibroadenoma of Breast|9012/0
C0334497|T191|SY|C4272|NCI|Pericanalicular Fibroadenoma of the Breast|9012/0
C0334497|T191|PT|BBM3.|RCD|Pericanalicular fibroadenoma|9012/0
C0334497|T191|PT|41382006|SNOMEDCT_US|Pericanalicular fibroadenoma|9012/0
C0001422|T191|PT|0000000711|CHV|adenofibroma|9013/0
C0001422|T191|SY|0000000711|CHV|adenofibromas|9013/0
C0001422|T191|LLT|10072991|MDR|Adenofibroma|9013/0
C0001422|T191|MH|D000232|MSH|Adenofibroma|9013/0
C0001422|T191|PM|D000232|MSH|Adenofibromas|9013/0
C0001422|T191|PN|NOCODE|MTH|Adenofibroma|9013/0
C4520837|T191|PT|C8984|NCI|Female Reproductive System Adenofibroma|9013/0
C4520837|T191|PT|C8984|NCI_CDISC|ADENOFIBROMA, BENIGN|9013/0
C4520837|T191|SY|C8984|NCI_CDISC|Benign Mixed Muellerian Tumor|9013/0
C0001422|T191|PT|Xa9A5|RCD|Adenofibroma|9013/0
C0001422|T191|SY|Xa9A5|RCDSY|Adenofibroma NOS|9013/0
C0001422|T191|PT|2962009|SNOMEDCT_US|Adenofibroma|9013/0
C0001422|T191|OAP|189823009|SNOMEDCT_US|Adenofibroma|9013/0
C0001422|T191|OF|189823009|SNOMEDCT_US|Adenofibroma|9013/0
C0001422|T191|SY|2962009|SNOMEDCT_US|Adenofibroma, no ICD-O subtype|9013/0
C0001422|T191|SY|2962009|SNOMEDCT_US|Adenofibroma, no International Classification of Diseases for Oncology subtype|9013/0
C0001422|T191|IS|2962009|SNOMEDCT_US|Adenofibroma, NOS|9013/0
C0334498|T191|PT|MTHU003432|ICPC2ICD10ENG|adenofibroma; serous, unspecified site|9014/0
C0334498|T191|PT|MTHU067547|ICPC2ICD10ENG|serous; adenofibroma, unspecified site|9014/0
C0334498|T191|PT|C67090|NCI|Serous Adenofibroma|9014/0
C0334498|T191|PT|BBM5.|RCD|Serous adenofibroma|9014/0
C0334498|T191|SY|BBM5.|RCD|Serous cystadenofibroma|9014/0
C3839174|T191|PT|703652007|SNOMEDCT_US|Seromucinous adenofibroma|9014/0
C0334498|T191|PT|2026006|SNOMEDCT_US|Serous adenofibroma|9014/0
C0334498|T191|SY|2026006|SNOMEDCT_US|Serous cystadenofibroma|9014/0
C1511266|T191|PT|C40028|NCI|Borderline Ovarian Serous Adenofibroma|9014/1
C1266152|T191|PT|128885004|SNOMEDCT_US|Serous adenofibroma of borderline malignancy|9014/1
C1266152|T191|SY|128885004|SNOMEDCT_US|Serous cystadenofibroma of borderline malignancy|9014/1
C2212013|T191|PT|233166|MEDCIN|serous adenocarcinofibroma of ovary|9014/3
C2212013|T191|PT|C67092|NCI|Ovarian Serous Adenocarcinofibroma|9014/3
C1266153|T191|SY|128886003|SNOMEDCT_US|Malignant serous adenofibroma|9014/3
C1266153|T191|SY|128886003|SNOMEDCT_US|Malignant serous cystadenofibroma|9014/3
C1266153|T191|PT|128886003|SNOMEDCT_US|Serous adenocarcinofibroma|9014/3
C1266153|T191|SY|128886003|SNOMEDCT_US|Serous cystadenocarcinofibroma|9014/3
C0334499|T191|PT|C8978|NCI|Mucinous Adenofibroma|9015/0
C0334499|T191|PT|BBM6.|RCD|Mucinous adenofibroma|9015/0
C0334499|T191|PT|10705005|SNOMEDCT_US|Mucinous adenofibroma|9015/0
C1881912|T191|PT|C66775|NCI|Borderline Ovarian Mucinous Adenofibroma|9015/1
C1881912|T191|SY|C66775|NCI|Ovarian Mucinous Adenofibroma of Borderline Malignancy|9015/1
C1266154|T191|PT|128887007|SNOMEDCT_US|Mucinous adenofibroma of borderline malignancy|9015/1
C1266154|T191|SY|128887007|SNOMEDCT_US|Mucinous cystadenofibroma of borderline malignancy|9015/1
C2212014|T191|PT|233167|MEDCIN|mucinous adenocarcinofibroma of ovary|9015/3
C2212014|T191|PT|C40034|NCI|Ovarian Mucinous Adenocarcinofibroma|9015/3
C2212014|T191|SY|C40034|NCI|Ovarian Mucinous Malignant Adenofibroma|9015/3
C1266155|T191|SY|128888002|SNOMEDCT_US|Malignant mucinous adenofibroma|9015/3
C1266155|T191|SY|128888002|SNOMEDCT_US|Malignant mucinous cystadenofibroma|9015/3
C1266155|T191|PT|128888002|SNOMEDCT_US|Mucinous adenocarcinofibroma|9015/3
C1266155|T191|SY|128888002|SNOMEDCT_US|Mucinous cystadenocarcinofibroma|9015/3
C0334500|T191|PN|NOCODE|MTH|Giant fibroadenoma|9016/0
C0346157|T191|PN|NOCODE|MTH|Giant fibroadenoma of breast|9016/0
C0346157|T191|PT|C4273|NCI|Breast Giant Fibroadenoma|9016/0
C0346157|T191|SY|C4273|NCI|Giant Breast Fibroadenoma|9016/0
C0346157|T191|SY|C4273|NCI|Giant Fibroadenoma|9016/0
C0346157|T191|SY|C4273|NCI|Giant Fibroadenoma of Breast|9016/0
C0346157|T191|SY|C4273|NCI|Giant Fibroadenoma of the Breast|9016/0
C0334500|T191|PT|X77ot|RCD|Giant fibroadenoma|9016/0
C0346157|T191|PT|X78WZ|RCD|Giant fibroadenoma of breast|9016/0
C0346157|T191|SY|X78WZ|RCD|Serocystic disease of Brodie|9016/0
C0334500|T191|OAP|189827005|SNOMEDCT_US|Giant fibroadenoma|9016/0
C0334500|T191|OF|189827005|SNOMEDCT_US|Giant fibroadenoma|9016/0
C0334500|T191|PT|34882000|SNOMEDCT_US|Giant fibroadenoma|9016/0
C0346157|T191|PT|254846003|SNOMEDCT_US|Giant fibroadenoma of breast|9016/0
C0346157|T191|SY|254846003|SNOMEDCT_US|Serocystic disease of Brodie|9016/0
C0334501|T191|PT|MTHU010311|ICPC2ICD10ENG|benign; Cystosarcoma phyllodes|9020/0
C0334501|T191|PT|MTHU020867|ICPC2ICD10ENG|Cystosarcoma phyllodes; benign|9020/0
C0334501|T191|PT|MTHU028166|ICPC2ICD10ENG|fibroadenoma; phyllodes|9020/0
C0334501|T191|PT|MTHU059414|ICPC2ICD10ENG|phyllodes; fibroadenoma|9020/0
C0334501|T191|PT|MTHU059416|ICPC2ICD10ENG|phyllodes; tumor, benign|9020/0
C0334501|T191|PT|MTHU077136|ICPC2ICD10ENG|tumor; phyllodes, benign|9020/0
C0334501|T191|SY|C4274|NCI|Benign Cystosarcoma Phyllodes|9020/0
C0334501|T191|SY|C4274|NCI|Benign Phyllodes Neoplasm|9020/0
C0334501|T191|PT|C4274|NCI|Benign Phyllodes Tumor|9020/0
C0334501|T191|SY|Xa9A6|RCD|Benign cystosarcoma phyllodes|9020/0
C0334501|T191|PT|Xa9A6|RCD|Benign phyllodes tumour|9020/0
C0334501|T191|PT|Xa9A6|RCDAE|Benign phyllodes tumor|9020/0
C0334501|T191|SY|16566002|SNOMEDCT_US|Benign cystosarcoma phyllodes|9020/0
C0334501|T191|PT|16566002|SNOMEDCT_US|Benign phyllodes tumor|9020/0
C0334501|T191|PTGB|16566002|SNOMEDCT_US|Benign phyllodes tumour|9020/0
C0334501|T191|SY|16566002|SNOMEDCT_US|Cystosarcoma phyllodes, benign|9020/0
C0334501|T191|SY|16566002|SNOMEDCT_US|Phyllodes tumor, benign|9020/0
C0334501|T191|SYGB|16566002|SNOMEDCT_US|Phyllodes tumour, benign|9020/0
C1370913|T191|SY|C7503|NCI|Borderline Phyllodes Neoplasm|9020/1
C1370913|T191|PT|C7503|NCI|Borderline Phyllodes Tumor|9020/1
C1370913|T191|SY|71232009|SNOMEDCT_US|Borderline cystosarcoma phyllodes|9020/1
C1370913|T191|PT|71232009|SNOMEDCT_US|Borderline phyllodes tumor|9020/1
C1370913|T191|PTGB|71232009|SNOMEDCT_US|Borderline phyllodes tumour|9020/1
C1370913|T191|SY|71232009|SNOMEDCT_US|Phyllodes tumor, borderline|9020/1
C1370913|T191|SYGB|71232009|SNOMEDCT_US|Phyllodes tumour, borderline|9020/1
C0600066|T191|PT|0000029998|CHV|malignant phyllodes tumor|9020/3
C0600066|T191|SY|0000029998|CHV|phyllodes malignant tumor|9020/3
C0600066|T191|PM|D003557|MSH|Cystosarcoma Phyllodes, Malignant|9020/3
C0600066|T191|PEP|D003557|MSH|Malignant Cystosarcoma Phyllodes|9020/3
C0600066|T191|PN|NOCODE|MTH|Malignant Cystosarcoma Phyllodes|9020/3
C0600066|T191|SY|C4275|NCI|Malignant Cystosarcoma Phyllodes|9020/3
C0600066|T191|SY|C4275|NCI|Malignant Phyllodes Neoplasm|9020/3
C0600066|T191|PT|C4275|NCI|Malignant Phyllodes Tumor|9020/3
C0600066|T191|OA|BBM9.|RCD|Malig cystosarcoma phyllodes|9020/3
C0600066|T191|OP|BBM9.|RCD|Malignant cystosarcoma phyllodes|9020/3
C0600066|T191|PT|Xa9A8|RCD|Malignant phyllodes tumour|9020/3
C0600066|T191|PT|Xa9A8|RCDAE|Malignant phyllodes tumor|9020/3
C0600066|T191|SY|87913009|SNOMEDCT_US|Cystosarcoma phyllodes, malignant|9020/3
C0600066|T191|SY|87913009|SNOMEDCT_US|Malignant cystosarcoma phyllodes|9020/3
C0600066|T191|OAP|189826001|SNOMEDCT_US|Malignant cystosarcoma phyllodes|9020/3
C0600066|T191|PT|87913009|SNOMEDCT_US|Malignant phyllodes tumor|9020/3
C0600066|T191|OAP|134331008|SNOMEDCT_US|Malignant phyllodes tumor|9020/3
C0600066|T191|PTGB|87913009|SNOMEDCT_US|Malignant phyllodes tumour|9020/3
C0600066|T191|OAP|134331008|SNOMEDCT_US|Malignant phyllodes tumour|9020/3
C3839630|T191|PT|703653002|SNOMEDCT_US|Periductal stromal tumor, low grade|9020/3
C3839630|T191|PTGB|703653002|SNOMEDCT_US|Periductal stromal tumour, low grade|9020/3
C0600066|T191|SY|87913009|SNOMEDCT_US|Phyllodes tumor, malignant|9020/3
C0600066|T191|SYGB|87913009|SNOMEDCT_US|Phyllodes tumour, malignant|9020/3
C0346158|T191|PT|MTHU028163|ICPC2ICD10ENG|fibroadenoma; juvenile|9030/0
C0346158|T191|PT|MTHU040682|ICPC2ICD10ENG|juvenile; fibroadenoma|9030/0
C0346158|T191|PT|C4276|NCI|Breast Juvenile Fibroadenoma|9030/0
C0346158|T191|SY|C4276|NCI|Cellular Fibroadenoma|9030/0
C0346158|T191|SY|C4276|NCI|Juvenile Breast Fibroadenoma|9030/0
C0346158|T191|SY|C4276|NCI|Juvenile Fibroadenoma|9030/0
C0346158|T191|SY|C4276|NCI|Juvenile Fibroadenoma of Breast|9030/0
C0346158|T191|SY|C4276|NCI|Juvenile Fibroadenoma of the Breast|9030/0
C0346158|T191|PT|BBMA.|RCD|Juvenile fibroadenoma|9030/0
C0346158|T191|AB|X78Wa|RCD|Juvenile fibroadenoma breast|9030/0
C0346158|T191|PT|X78Wa|RCD|Juvenile fibroadenoma of breast|9030/0
C0346158|T191|SY|46212000|SNOMEDCT_US|Cellular fibroadenoma|9030/0
C0346158|T191|PT|46212000|SNOMEDCT_US|Juvenile fibroadenoma|9030/0
C0346158|T191|PT|254847007|SNOMEDCT_US|Juvenile fibroadenoma of breast|9030/0
C0221289|T047|SY|NOCODE|DXP|SYNOVIOMA, BENIGN|9040/0
C0221289|T047|SY|C3829|NCI|Benign Neoplasm of Synovium|9040/0
C0221289|T047|SY|C3829|NCI|Benign Neoplasm of the Synovium|9040/0
C0221289|T047|PT|C3829|NCI|Benign Synovial Neoplasm|9040/0
C0221289|T047|SY|C3829|NCI|Benign Synovial Tumor|9040/0
C0221289|T047|SY|C3829|NCI|Benign Synovioma|9040/0
C0221289|T047|SY|C3829|NCI|Benign Tumor of Synovium|9040/0
C0221289|T047|SY|C3829|NCI|Benign Tumor of the Synovium|9040/0
C0221289|T047|SY|C3829|NCI_CDISC|Benign Neoplasm of Synovium|9040/0
C0221289|T047|SY|C3829|NCI_CDISC|Benign Neoplasm of the Synovium|9040/0
C0221289|T047|SY|C3829|NCI_CDISC|Benign Synovial Tumor|9040/0
C0221289|T047|SY|C3829|NCI_CDISC|Benign Synovioma|9040/0
C0221289|T047|SY|C3829|NCI_CDISC|Benign Tumor of Synovium|9040/0
C0221289|T047|SY|C3829|NCI_CDISC|Benign Tumor of the Synovium|9040/0
C0221289|T047|PT|C3829|NCI_CDISC|SYNOVIOMA, BENIGN|9040/0
C0221289|T047|PT|BBN0.|RCD|Benign synovioma|9040/0
C0221289|T047|SY|5178002|SNOMEDCT_US|Benign synovioma|9040/0
C0221289|T047|PT|5178002|SNOMEDCT_US|Synovioma, benign|9040/0
C0039101|T191|SY|0000011982|CHV|sarcoma synovial|9040/3
C0039101|T191|PT|0000011982|CHV|synovial sarcoma|9040/3
C0039101|T191|SY|0000011982|CHV|synovioma|9040/3
C0039101|T191|SY|HP:0012570|HPO|Malignant synovioma|9040/3
C0039101|T191|PT|HP:0012570|HPO|Synovial sarcoma|9040/3
C0039101|T191|PT|U004562|LCH|Synovioma|9040/3
C0039101|T191|PT|sh85131651|LCH_NW|Synovioma|9040/3
C0039101|T191|LLT|10042863|MDR|Synovial sarcoma|9040/3
C0039101|T191|PT|10042863|MDR|Synovial sarcoma|9040/3
C0039101|T191|LLT|10042866|MDR|Synovial sarcoma NOS|9040/3
C0039101|T191|LLT|10069062|MDR|Synovioma|9040/3
C0039101|T191|PT|271501|MEDCIN|synovial sarcoma|9040/3
C0039101|T191|PT|231888|MEDCIN|synovial sarcoma of soft tissue|9040/3
C0039101|T191|SY|31580|MEDCIN|synovioma|9040/3
C0039101|T191|PT|31580|MEDCIN|synovioma of joint|9040/3
C0039101|T191|MH|D013584|MSH|Sarcoma, Synovial|9040/3
C0039101|T191|PM|D013584|MSH|Sarcomas, Synovial|9040/3
C0039101|T191|PM|D013584|MSH|Synovial Sarcoma|9040/3
C0039101|T191|PM|D013584|MSH|Synovial Sarcomas|9040/3
C0039101|T191|ET|D013584|MSH|Synovioma|9040/3
C0039101|T191|PM|D013584|MSH|Synoviomas|9040/3
C0039101|T191|PN|NOCODE|MTH|synovial sarcoma|9040/3
C0039101|T191|AB|C3400|NCI|SS|9040/3
C0039101|T191|PT|C3400|NCI|Synovial Sarcoma|9040/3
C0039101|T191|SY|C3400|NCI|Synovial Sarcoma, NOS|9040/3
C0039101|T191|SY|C3400|NCI|Synovial Sarcoma, Not Otherwise Specified|9040/3
C0039101|T191|PT|C3400|NCI_CDISC|SARCOMA, SYNOVIAL, MALIGNANT|9040/3
C0039101|T191|SY|C3400|NCI_CDISC|SS|9040/3
C0039101|T191|PT|10042866|NCI_CTEP-SDC|Synovial sarcoma|9040/3
C0039101|T191|DN|C3400|NCI_CTRP|Synovial Sarcoma|9040/3
C0039101|T191|PT|CDR0000044626|NCI_NCI-GLOSS|synovial sarcoma|9040/3
C0039101|T191|SY|Xa9A9|RCD|Malignant synovioma|9040/3
C0039101|T191|PT|Xa9A9|RCD|Synovial sarcoma|9040/3
C0039101|T191|SY|BBN1.|RCDSY|Synovial sarcoma NOS|9040/3
C0039101|T191|PT|BBN1.|RCDSY|Synovioma NOS|9040/3
C0039101|T191|SY|302851001|SNOMEDCT_US|Malignant synovioma|9040/3
C0039101|T191|PT|302851001|SNOMEDCT_US|Synovial sarcoma|9040/3
C0039101|T191|PT|63211008|SNOMEDCT_US|Synovial sarcoma|9040/3
C1959647|T191|PT|425535000|SNOMEDCT_US|Synovial sarcoma - category|9040/3
C0039101|T191|IS|63211008|SNOMEDCT_US|Synovial sarcoma, NOS|9040/3
C0039101|T191|SY|63211008|SNOMEDCT_US|Synovioma|9040/3
C0039101|T191|SY|63211008|SNOMEDCT_US|Synovioma, malignant|9040/3
C0039101|T191|IS|63211008|SNOMEDCT_US|Synovioma, NOS|9040/3
C0334505|T191|PT|271503|MEDCIN|spindle cell synovial sarcoma|9041/3
C0334505|T191|SY|271503|MEDCIN|synovial spindle cell sarcoma|9041/3
C0334505|T191|PT|C4277|NCI|Spindle Cell Synovial Sarcoma|9041/3
C0334505|T191|SY|C4277|NCI|Synovial Sarcoma with Spindle Cell Components|9041/3
C0334505|T191|PT|BBN2.|RCD|Synovial sarcoma - spindle cell|9041/3
C0334505|T191|AB|BBN2.|RCD|Synovial sarcoma-spindle cell|9041/3
C0334505|T191|SY|37206003|SNOMEDCT_US|Synovial sarcoma - spindle cell|9041/3
C0334505|T191|SY|37206003|SNOMEDCT_US|Synovial sarcoma, monophasic fibrous|9041/3
C0334505|T191|PT|37206003|SNOMEDCT_US|Synovial sarcoma, spindle cell|9041/3
C0334506|T191|PT|271504|MEDCIN|epithelioid cell synovial sarcoma|9042/3
C0334506|T191|SY|271504|MEDCIN|synovial epithelioid cell sarcoma|9042/3
C0334506|T191|SY|C4278|NCI|Epithelial Sarcoma of Synovium|9042/3
C0334506|T191|SY|C4278|NCI|Epithelial Sarcoma of the Synovium|9042/3
C0334506|T191|PT|C4278|NCI|Epithelial Synovial Sarcoma|9042/3
C0334506|T191|SY|C4278|NCI|Epithelioid Cell Sarcoma of Synovium|9042/3
C0334506|T191|SY|C4278|NCI|Epithelioid Cell Sarcoma of the Synovium|9042/3
C0334506|T191|SY|C4278|NCI|Epithelioid Cell Synovial Sarcoma|9042/3
C0334506|T191|SY|C4278|NCI|Epithelioid Synovial Sarcoma|9042/3
C0334506|T191|AB|BBN3.|RCD|Synov sarcoma-epithelioid cell|9042/3
C0334506|T191|PT|BBN3.|RCD|Synovial sarcoma - epithelioid cell|9042/3
C0334506|T191|SY|56422000|SNOMEDCT_US|Synovial sarcoma - epithelioid cell|9042/3
C0334506|T191|PT|56422000|SNOMEDCT_US|Synovial sarcoma, epithelioid cell|9042/3
C0334507|T191|PT|271505|MEDCIN|biphasic synovial sarcoma|9043/3
C0334507|T191|SY|C4279|NCI|Biphasic Sarcoma of Synovium|9043/3
C0334507|T191|SY|C4279|NCI|Biphasic Sarcoma of the Synovium|9043/3
C0334507|T191|PT|C4279|NCI|Biphasic Synovial Sarcoma|9043/3
C0334507|T191|PT|BBN4.|RCD|Synovial sarcoma - biphasic|9043/3
C0334507|T191|SY|18588008|SNOMEDCT_US|Synovial sarcoma - biphasic|9043/3
C0334507|T191|PT|18588008|SNOMEDCT_US|Synovial sarcoma, biphasic|9043/3
C0206651|T191|LLT|10065865|MDR|Clear cell sarcoma|9044/3
C0206651|T191|PT|10073140|MDR|Clear cell sarcoma of soft tissue|9044/3
C0206651|T191|LLT|10073140|MDR|Clear cell sarcoma of soft tissue|9044/3
C0206651|T191|PT|271506|MEDCIN|clear cell sarcoma|9044/3
C0206651|T191|PT|231892|MEDCIN|clear cell sarcoma of soft tissue|9044/3
C0206651|T191|PT|352929|MEDCIN|malignant melanoma of soft tissue|9044/3
C0206651|T191|SY|352929|MEDCIN|soft tissue neoplasm malignant melanoma|9044/3
C0206651|T191|PM|D018227|MSH|Clear Cell Sarcoma|9044/3
C0206651|T191|ET|D018227|MSH|Clear Cell Sarcoma of Soft Tissue|9044/3
C0206651|T191|PM|D018227|MSH|Clear Cell Sarcomas|9044/3
C0206651|T191|ET|D018227|MSH|Malignant Melanoma of Soft Parts|9044/3
C0206651|T191|ET|D018227|MSH|Melanoma of Soft Parts|9044/3
C0206651|T191|ET|D018227|MSH|Melanoma, Malignant, of Soft Parts|9044/3
C0206651|T191|MH|D018227|MSH|Sarcoma, Clear Cell|9044/3
C0206651|T191|PM|D018227|MSH|Sarcomas, Clear Cell|9044/3
C0206651|T191|PN|NOCODE|MTH|Clear Cell Sarcoma of Soft Tissue|9044/3
C0206651|T191|SY|C3745|NCI|Chordoid Sarcoma|9044/3
C0206651|T191|SY|C3745|NCI|Clear Cell Sarcoma of Soft Parts|9044/3
C0206651|T191|PT|C3745|NCI|Clear Cell Sarcoma of Soft Tissue|9044/3
C0206651|T191|SY|C3745|NCI|Malignant Melanoma of Soft Parts|9044/3
C0206651|T191|SY|C3745|NCI|Malignant Melanoma of the Soft Parts|9044/3
C0206651|T191|SY|10065865|NCI_CTEP-SDC|Clear cell sarcoma - not kidney|9044/3
C0206651|T191|PT|CDR0000641939|NCI_NCI-GLOSS|clear cell sarcoma of soft tissue|9044/3
C0206651|T191|PT|CDR0000656145|NCI_NCI-GLOSS|malignant melanoma of soft parts|9044/3
C0206651|T191|PT|XM0Af|RCD|Clear cell sarcoma|9044/3
C0206651|T191|AB|XM0Af|RCD|Malig melanoma of soft tissue|9044/3
C0206651|T191|SY|XM0Af|RCD|Malignant melanoma of soft tissue|9044/3
C0206651|T191|PT|271944004|SNOMEDCT_US|Clear cell sarcoma|9044/3
C0206651|T191|SY|402561003|SNOMEDCT_US|Clear cell sarcoma|9044/3
C0206651|T191|SY|271944004|SNOMEDCT_US|Malignant melanoma of soft tissue|9044/3
C0206651|T191|PT|402561003|SNOMEDCT_US|Malignant melanoma of soft tissues|9044/3
C0206651|T191|SY|12622007|SNOMEDCT_US|Melanoma, malignant, of soft parts|9044/3
C0206675|T191|NP|0000023024|AOD|adenomatoid tumor|9050/0
C0206675|T191|PT|0000021013|CHV|adenomatoid tumor|9050/0
C0206675|T191|SY|0000021013|CHV|adenomatoid tumors|9050/0
C0206675|T191|ET|D19.9|ICD10CM|Benign mesothelioma NOS|9050/0
C0206675|T191|PT|10061691|MDR|Benign mesothelioma|9050/0
C0206675|T191|LLT|10061691|MDR|Benign mesothelioma|9050/0
C0206675|T191|LLT|10004291|MDR|Benign mesothelioma NOS|9050/0
C0206675|T191|HT|10027413|MDR|Mesotheliomas benign|9050/0
C0206675|T191|MH|D018254|MSH|Adenomatoid Tumor|9050/0
C0206675|T191|PM|D018254|MSH|Adenomatoid Tumors|9050/0
C0206675|T191|PM|D018254|MSH|Tumor, Adenomatoid|9050/0
C0206675|T191|PM|D018254|MSH|Tumors, Adenomatoid|9050/0
C0206675|T191|PT|C3762|NCI|Adenomatoid Tumor|9050/0
C0206675|T191|SY|C3762|NCI|Benign Localized Epithelial Mesothelioma|9050/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelial Neoplasm|9050/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelial Tumor|9050/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelioma|9050/0
C0206675|T191|SY|C3762|NCI|Benign Neoplasm of Mesothelium|9050/0
C0206675|T191|SY|C3762|NCI|Benign Neoplasm of the Mesothelium|9050/0
C0206675|T191|SY|C3762|NCI|Benign Tumor of Mesothelium|9050/0
C0206675|T191|SY|C3762|NCI|Benign Tumor of the Mesothelium|9050/0
C0206675|T191|SY|C3762|NCI|Mesothelioma, Benign|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Adenomatoid Tumor, Benign|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Localized Epithelial Mesothelioma|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelial Neoplasm|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelial Tumor|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelioma|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Neoplasm of Mesothelium|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Neoplasm of the Mesothelium|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Tumor of Mesothelium|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Tumor of the Mesothelium|9050/0
C0206675|T191|PT|C3762|NCI_CDISC|MESOTHELIOMA, BENIGN|9050/0
C0206675|T191|SY|C3762|NCI_CDISC|Mesothelioma, Benign|9050/0
C0206675|T191|PT|Xa9AD|RCD|Adenomatoid tumour|9050/0
C0334514|T191|PT|BBP6.|RCD|Benign biphasic mesothelioma|9050/0
C0206675|T191|PT|BBP0.|RCD|Benign mesothelioma|9050/0
C0206675|T191|PT|Xa9AD|RCDAE|Adenomatoid tumor|9050/0
C0206675|T191|OP|BBP8.|RCDSA|Adenomatoid tumor NOS|9050/0
C0206675|T191|OP|BBP8.|RCDSY|Adenomatoid tumour NOS|9050/0
C0206675|T191|PT|2348006|SNOMEDCT_US|Adenomatoid tumor|9050/0
C0206675|T191|IS|2348006|SNOMEDCT_US|Adenomatoid tumor, NOS|9050/0
C0206675|T191|PTGB|2348006|SNOMEDCT_US|Adenomatoid tumour|9050/0
C0334514|T191|PT|189833001|SNOMEDCT_US|Benign biphasic mesothelioma|9050/0
C0206675|T191|SY|41183007|SNOMEDCT_US|Benign mesothelioma|9050/0
C0206675|T191|PT|41183007|SNOMEDCT_US|Mesothelioma, benign|9050/0
C0334514|T191|OAP|34762006|SNOMEDCT_US|Mesothelioma, biphasic, benign|9050/0
C0334514|T191|IS|34762006|SNOMEDCT_US|Mesothelioma, biphasic, benign -RETIRED-|9050/0
C0334514|T191|OF|34762006|SNOMEDCT_US|Mesothelioma, biphasic, benign -RETIRED-|9050/0
C0345967|T191|PT|0000031033|CHV|malignant mesothelioma|9050/3
C0345967|T191|PT|HP:0100001|HPO|Malignant mesothelioma|9050/3
C0345967|T191|LLT|10027407|MDR|Mesothelioma malignant|9050/3
C0345967|T191|PT|10027407|MDR|Mesothelioma malignant|9050/3
C0345967|T191|LLT|10027410|MDR|Mesothelioma malignant NOS|9050/3
C0345967|T191|SY|335197|MEDCIN|malignant neoplasm mesothelioma|9050/3
C0345967|T191|PT|335197|MEDCIN|mesothelioma|9050/3
C0345967|T191|SY|4014|MEDLINEPLUS|Malignant mesothelioma|9050/3
C0345967|T191|NM|C562839|MSH|Mesothelioma, Malignant|9050/3
C0345967|T191|PN|NOCODE|MTH|Malignant mesothelioma|9050/3
C0345967|T191|SY|C4456|NCI|Malignant Mesothelial Neoplasm|9050/3
C0345967|T191|SY|C4456|NCI|Malignant Mesothelial Tumor|9050/3
C0345967|T191|PT|C4456|NCI|Malignant Mesothelioma|9050/3
C0345967|T191|SY|C4456|NCI|Malignant Neoplasm of Mesothelium|9050/3
C0345967|T191|SY|C4456|NCI|Malignant Neoplasm of the Mesothelium|9050/3
C0345967|T191|SY|C4456|NCI|Malignant Tumor of Mesothelium|9050/3
C0345967|T191|SY|C4456|NCI|Malignant Tumor of the Mesothelium|9050/3
C0345967|T191|SY|C4456|NCI_CDISC|Malignant Mesothelial Neoplasm|9050/3
C0345967|T191|SY|C4456|NCI_CDISC|Malignant Mesothelial Tumor|9050/3
C0345967|T191|SY|C4456|NCI_CDISC|Malignant Neoplasm of Mesothelium|9050/3
C0345967|T191|SY|C4456|NCI_CDISC|Malignant Neoplasm of the Mesothelium|9050/3
C0345967|T191|SY|C4456|NCI_CDISC|Malignant Tumor of Mesothelium|9050/3
C0345967|T191|SY|C4456|NCI_CDISC|Malignant Tumor of the Mesothelium|9050/3
C0345967|T191|PT|C4456|NCI_CDISC|MESOTHELIOMA, MALIGNANT|9050/3
C0345967|T191|PT|C4456|NCI_CPTAC|Malignant Mesothelioma|9050/3
C0345967|T191|DN|C4456|NCI_CTRP|Malignant Mesothelioma|9050/3
C0345967|T191|PT|CDR0000044992|NCI_NCI-GLOSS|malignant mesothelioma|9050/3
C0345967|T191|PSC|CDR0000038142|PDQ|malignant mesothelioma|9050/3
C0345967|T191|SY|CDR0000038142|PDQ|mesothelioma, malignant|9050/3
C0345967|T191|PT|BBP1.|RCD|Malignant mesothelioma|9050/3
C0345967|T191|SY|109378008|SNOMEDCT_US|Cancer, mesothelioma|9050/3
C0345967|T191|SY|109378008|SNOMEDCT_US|Malignant mesothelioma|9050/3
C0345967|T191|SY|62064005|SNOMEDCT_US|Malignant mesothelioma|9050/3
C0345967|T191|PT|62064005|SNOMEDCT_US|Mesothelioma, malignant|9050/3
C1266119|T191|PT|0000056686|CHV|solitary fibrous tumor|9051/0
C1266119|T191|SY|0000056686|CHV|solitary fibrous tumour|9051/0
C1266119|T191|LLT|10024773|MDR|Localised fibrous mesothelioma|9051/0
C1266119|T191|LLT|10062468|MDR|Localized fibrous mesothelioma|9051/0
C1266119|T191|LLT|10082807|MDR|Solitary fibrous tumor|9051/0
C1266119|T191|MTH_PT|10082804|MDR|Solitary fibrous tumor|9051/0
C1266119|T191|LLT|10082804|MDR|Solitary fibrous tumour|9051/0
C1266119|T191|PT|10082804|MDR|Solitary fibrous tumour|9051/0
C0334511|T191|ET|D054363|MSH|Benign Fibrous Mesothelioma|9051/0
C0334511|T191|PM|D054363|MSH|Benign Fibrous Mesotheliomas|9051/0
C0334511|T191|PM|D054363|MSH|Fibroma, Submesothelial|9051/0
C0334511|T191|PM|D054363|MSH|Fibromas, Submesothelial|9051/0
C0334511|T191|ET|D054363|MSH|Fibrous Mesothelioma|9051/0
C0334511|T191|PM|D054363|MSH|Fibrous Mesothelioma, Benign|9051/0
C0334511|T191|PM|D054363|MSH|Fibrous Mesothelioma, Localized|9051/0
C0334511|T191|PM|D054363|MSH|Fibrous Mesothelioma, Solitary|9051/0
C0334511|T191|PM|D054363|MSH|Fibrous Mesotheliomas|9051/0
C0334511|T191|PM|D054363|MSH|Fibrous Mesotheliomas, Benign|9051/0
C0334511|T191|PM|D054363|MSH|Fibrous Mesotheliomas, Localized|9051/0
C0334511|T191|PM|D054363|MSH|Fibrous Mesotheliomas, Solitary|9051/0
C1266119|T191|PM|D054364|MSH|Fibrous Tumor, Solitary|9051/0
C1266119|T191|PM|D054364|MSH|Fibrous Tumors, Solitary|9051/0
C0334511|T191|ET|D054363|MSH|Localized Fibrous Mesothelioma|9051/0
C0334511|T191|PM|D054363|MSH|Localized Fibrous Mesotheliomas|9051/0
C0334511|T191|ET|D054363|MSH|Localized Mesothelioma|9051/0
C0334511|T191|PM|D054363|MSH|Localized Mesotheliomas|9051/0
C0334511|T191|PM|D054363|MSH|Mesothelioma, Benign Fibrous|9051/0
C0334511|T191|PM|D054363|MSH|Mesothelioma, Fibrous|9051/0
C0334511|T191|PM|D054363|MSH|Mesothelioma, Localized|9051/0
C0334511|T191|PM|D054363|MSH|Mesothelioma, Localized Fibrous|9051/0
C0334511|T191|PM|D054363|MSH|Mesothelioma, Solitary Fibrous|9051/0
C0334511|T191|PM|D054363|MSH|Mesotheliomas, Benign Fibrous|9051/0
C0334511|T191|PM|D054363|MSH|Mesotheliomas, Fibrous|9051/0
C0334511|T191|PM|D054363|MSH|Mesotheliomas, Localized|9051/0
C0334511|T191|PM|D054363|MSH|Mesotheliomas, Localized Fibrous|9051/0
C0334511|T191|PM|D054363|MSH|Mesotheliomas, Solitary Fibrous|9051/0
C0334511|T191|ET|D054363|MSH|Solitary Fibrous Mesothelioma|9051/0
C0334511|T191|PM|D054363|MSH|Solitary Fibrous Mesotheliomas|9051/0
C1266119|T191|PM|D054364|MSH|Solitary Fibrous Tumor|9051/0
C0334511|T191|ET|D054363|MSH|Solitary Fibrous Tumor of the Pleura|9051/0
C0334511|T191|MH|D054363|MSH|Solitary Fibrous Tumor, Pleural|9051/0
C1266119|T191|MH|D054364|MSH|Solitary Fibrous Tumors|9051/0
C0334511|T191|ET|D054363|MSH|Submesothelial Fibroma|9051/0
C0334511|T191|PM|D054363|MSH|Submesothelial Fibromas|9051/0
C1266119|T191|PM|D054364|MSH|Tumor, Solitary Fibrous|9051/0
C1266119|T191|PM|D054364|MSH|Tumors, Solitary Fibrous|9051/0
C0334511|T191|PN|NOCODE|MTH|Pleural Solitary Fibrous Tumor|9051/0
C1266119|T191|PN|NOCODE|MTH|Solitary fibrous tumor|9051/0
C0334511|T191|SY|C4457|NCI|Fibroma of Pleura|9051/0
C0334511|T191|SY|C4457|NCI|Fibroma of the Pleura|9051/0
C1266119|T191|OP|C7634|NCI|Hemangiopericytoma|9051/0
C1266119|T191|OP|C7634|NCI|Localized Fibrous Mesothelioma|9051/0
C0334511|T191|OP|C4457|NCI|Localized Fibrous Mesothelioma of Pleura|9051/0
C0334511|T191|OP|C4457|NCI|Localized Fibrous Mesothelioma of the Pleura|9051/0
C1266119|T191|SY|C7634|NCI|Localized Fibrous Tumor|9051/0
C0334511|T191|SY|C4457|NCI|Pleural Fibroma|9051/0
C0334511|T191|PT|C4457|NCI|Pleural Solitary Fibrous Tumor|9051/0
C0334511|T191|OP|C4457|NCI|Pleural Submesothelial Fibroma|9051/0
C1266119|T191|AB|C7634|NCI|SFT|9051/0
C1266119|T191|PT|C7634|NCI|Solitary Fibrous Tumor|9051/0
C0334511|T191|SY|C4457|NCI|Solitary Fibrous Tumor of Pleura|9051/0
C0334511|T191|SY|C4457|NCI|Solitary Fibrous Tumor of the Pleura|9051/0
C1266119|T191|OP|C7634|NCI|Submesothelial Fibroma|9051/0
C0334511|T191|PT|BBP2.|RCD|Benign fibrous mesothelioma|9051/0
C0334511|T191|PT|X78Qe|RCD|Pleural fibroma|9051/0
C0334511|T191|SY|15702005|SNOMEDCT_US|Benign fibrous mesothelioma|9051/0
C0334511|T191|PT|15702005|SNOMEDCT_US|Fibrous mesothelioma, benign|9051/0
C1266119|T191|SYGB|128736003|SNOMEDCT_US|Localised fibrous tumour|9051/0
C0334511|T191|SYGB|254646001|SNOMEDCT_US|Localised fibrous tumour of pleura|9051/0
C1266119|T191|SY|128736003|SNOMEDCT_US|Localized fibrous tumor|9051/0
C0334511|T191|SY|254646001|SNOMEDCT_US|Localized fibrous tumor of pleura|9051/0
C0334511|T191|PT|254646001|SNOMEDCT_US|Pleural fibroma|9051/0
C1266119|T191|PT|128736003|SNOMEDCT_US|Solitary fibrous tumor|9051/0
C0334511|T191|SY|254646001|SNOMEDCT_US|Solitary fibrous tumor of pleura|9051/0
C1266119|T191|PTGB|128736003|SNOMEDCT_US|Solitary fibrous tumour|9051/0
C0334511|T191|SYGB|254646001|SNOMEDCT_US|Solitary fibrous tumour of pleura|9051/0
C0334513|T191|PT|0000029999|CHV|sarcomatoid mesothelioma|9051/3
C0334513|T191|SY|0000029999|CHV|sarcomatous mesothelioma|9051/3
C0334513|T191|PT|MTHU028115|ICPC2ICD10ENG|fibrous; mesothelioma|9051/3
C0334513|T191|PT|MTHU048955|ICPC2ICD10ENG|mesothelioma; fibrous|9051/3
C1270206|T191|LLT|10073063|MDR|Desmoplastic mesothelioma|9051/3
C1270206|T191|PT|10073063|MDR|Desmoplastic mesothelioma|9051/3
C0334513|T191|LLT|10073065|MDR|Sarcomatoid mesothelioma|9051/3
C0334513|T191|PT|10073065|MDR|Sarcomatoid mesothelioma|9051/3
C0334513|T191|PN|NOCODE|MTH|Sarcomatoid Mesothelioma|9051/3
C1270206|T191|PT|C6747|NCI|Desmoplastic Mesothelioma|9051/3
C0334513|T191|PT|C45655|NCI|Sarcomatoid Mesothelioma|9051/3
C1270206|T191|DN|C6747|NCI_CTRP|Desmoplastic Mesothelioma|9051/3
C0334513|T191|DN|C45655|NCI_CTRP|Sarcomatoid Mesothelioma|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|fibrous mesothelial sarcoma|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|fibrous mesothelioma|9051/3
C0334513|T191|SY|CDR0000038142|PDQ|mesothelial sarcoma|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|mesothelial sarcoma, fibrous|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|mesothelial sarcoma, sarcomatous|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|mesothelioma, fibrous|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|mesothelioma, sarcomatous|9051/3
C0334513|T191|SY|CDR0000038142|PDQ|sarcoma, mesothelial|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|sarcoma, mesothelial, fibrous|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|sarcoma, mesothelial, sarcomatous|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|Sarcomatoid Mesothelioma|9051/3
C0334513|T191|SY|CDR0000039970|PDQ|sarcomatous mesothelial sarcoma|9051/3
C0334513|T191|PT|CDR0000039970|PDQ|sarcomatous mesothelioma|9051/3
C0334513|T191|SY|BBP3.|RCD|Fibrous mesothelioma|9051/3
C0334513|T191|PT|BBP3.|RCD|Malignant fibrous mesothelioma|9051/3
C1270206|T191|PT|388650006|SNOMEDCT_US|Desmoplastic mesothelioma|9051/3
C1270206|T191|SY|54443001|SNOMEDCT_US|Desmoplastic mesothelioma|9051/3
C0334513|T191|OAS|209241006|SNOMEDCT_US|Fibrous mesothelioma|9051/3
C0334513|T191|SY|54443001|SNOMEDCT_US|Fibrous mesothelioma|9051/3
C0334513|T191|PT|54443001|SNOMEDCT_US|Fibrous mesothelioma, malignant|9051/3
C0334513|T191|IS|54443001|SNOMEDCT_US|Fibrous mesothelioma, NOS|9051/3
C0334513|T191|OAP|209241006|SNOMEDCT_US|Malignant fibrous mesothelioma|9051/3
C0334513|T191|SY|54443001|SNOMEDCT_US|Sarcomatoid mesothelioma|9051/3
C0334513|T191|PT|399477001|SNOMEDCT_US|Sarcomatoid mesothelioma|9051/3
C0334513|T191|SY|54443001|SNOMEDCT_US|Spindled mesothelioma|9051/3
C0206675|T191|NP|0000023024|AOD|adenomatoid tumor|9052/0
C0206675|T191|PT|0000021013|CHV|adenomatoid tumor|9052/0
C0206675|T191|SY|0000021013|CHV|adenomatoid tumors|9052/0
C0206675|T191|ET|D19.9|ICD10CM|Benign mesothelioma NOS|9052/0
C0206675|T191|LLT|10061691|MDR|Benign mesothelioma|9052/0
C0206675|T191|PT|10061691|MDR|Benign mesothelioma|9052/0
C0206675|T191|LLT|10004291|MDR|Benign mesothelioma NOS|9052/0
C0206675|T191|HT|10027413|MDR|Mesotheliomas benign|9052/0
C0206675|T191|MH|D018254|MSH|Adenomatoid Tumor|9052/0
C0206675|T191|PM|D018254|MSH|Adenomatoid Tumors|9052/0
C0206675|T191|PM|D018254|MSH|Tumor, Adenomatoid|9052/0
C0206675|T191|PM|D018254|MSH|Tumors, Adenomatoid|9052/0
C0206675|T191|PT|C3762|NCI|Adenomatoid Tumor|9052/0
C0206675|T191|SY|C3762|NCI|Benign Localized Epithelial Mesothelioma|9052/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelial Neoplasm|9052/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelial Tumor|9052/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelioma|9052/0
C0206675|T191|SY|C3762|NCI|Benign Neoplasm of Mesothelium|9052/0
C0206675|T191|SY|C3762|NCI|Benign Neoplasm of the Mesothelium|9052/0
C0206675|T191|SY|C3762|NCI|Benign Tumor of Mesothelium|9052/0
C0206675|T191|SY|C3762|NCI|Benign Tumor of the Mesothelium|9052/0
C0206675|T191|SY|C3762|NCI|Mesothelioma, Benign|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Adenomatoid Tumor, Benign|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Localized Epithelial Mesothelioma|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelial Neoplasm|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelial Tumor|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelioma|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Neoplasm of Mesothelium|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Neoplasm of the Mesothelium|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Tumor of Mesothelium|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Tumor of the Mesothelium|9052/0
C0206675|T191|PT|C3762|NCI_CDISC|MESOTHELIOMA, BENIGN|9052/0
C0206675|T191|SY|C3762|NCI_CDISC|Mesothelioma, Benign|9052/0
C0206675|T191|PT|Xa9AD|RCD|Adenomatoid tumour|9052/0
C0334512|T191|AB|BBP4.|RCD|Benig epithelioid mesothelioma|9052/0
C0334512|T191|PT|BBP4.|RCD|Benign epithelioid mesothelioma|9052/0
C0206675|T191|PT|BBP0.|RCD|Benign mesothelioma|9052/0
C0206675|T191|PT|Xa9AD|RCDAE|Adenomatoid tumor|9052/0
C0206675|T191|OP|BBP8.|RCDSA|Adenomatoid tumor NOS|9052/0
C0206675|T191|OP|BBP8.|RCDSY|Adenomatoid tumour NOS|9052/0
C0206675|T191|PT|2348006|SNOMEDCT_US|Adenomatoid tumor|9052/0
C0206675|T191|IS|2348006|SNOMEDCT_US|Adenomatoid tumor, NOS|9052/0
C0206675|T191|PTGB|2348006|SNOMEDCT_US|Adenomatoid tumour|9052/0
C0334512|T191|SY|84919003|SNOMEDCT_US|Benign epithelioid mesothelioma|9052/0
C0206675|T191|SY|41183007|SNOMEDCT_US|Benign mesothelioma|9052/0
C0334512|T191|PT|84919003|SNOMEDCT_US|Epithelioid mesothelioma, benign|9052/0
C0334512|T191|SY|84919003|SNOMEDCT_US|Mesothelial papilloma|9052/0
C0206675|T191|PT|41183007|SNOMEDCT_US|Mesothelioma, benign|9052/0
C0334512|T191|IS|84919003|SNOMEDCT_US|Well differentiated papillary mesothelioma, benign|9052/0
C1337012|T191|SY|C7635|NCI|Benign/Intermediate Mesothelioma|9052/1
C1337012|T191|AB|C7635|NCI|WDPM|9052/1
C1337012|T191|PT|C7635|NCI|Well Differentiated Papillary Mesothelioma|9052/1
C1337012|T191|SY|C7635|NCI|Well-Differentiated Mesothelial Papillary Neoplasm|9052/1
C1337012|T191|SY|C7635|NCI|Well-Differentiated Mesothelial Papillary Tumor|9052/1
C1337012|T191|SY|C7635|NCI|Well-Differentiated Papillary Neoplasm of Mesothelium|9052/1
C1337012|T191|SY|C7635|NCI|Well-Differentiated Papillary Neoplasm of the Mesothelium|9052/1
C1337012|T191|SY|C7635|NCI|Well-Differentiated Papillary Tumor of Mesothelium|9052/1
C1337012|T191|SY|C7635|NCI|Well-Differentiated Papillary Tumor of the Mesothelium|9052/1
C1337012|T191|PT|734100004|SNOMEDCT_US|Well-differentiated papillary mesothelioma|9052/1
C0862312|T191|PT|MTHU026830|ICPC2ICD10ENG|epithelioid; mesothelioma|9052/3
C0862312|T191|PT|MTHU048947|ICPC2ICD10ENG|mesothelioma; epithelioid|9052/3
C0862312|T191|LLT|10015093|MDR|Epithelial malignant mesothelioma|9052/3
C0862312|T191|LLT|10073064|MDR|Epithelioid mesothelioma|9052/3
C0862312|T191|PT|10073064|MDR|Epithelioid mesothelioma|9052/3
C0862312|T191|SY|C7985|NCI|Epithelial Mesothelioma|9052/3
C0862312|T191|PT|C7985|NCI|Epithelioid Mesothelioma|9052/3
C0862312|T191|SY|C7985|NCI|Malignant Epithelial Mesothelioma|9052/3
C0862312|T191|DN|C7985|NCI_CTRP|Epithelioid Mesothelioma|9052/3
C0862312|T191|PT|CDR0000039969|PDQ|epithelial mesothelioma|9052/3
C0862312|T191|SY|CDR0000039969|PDQ|Epithelioid Mesothelioma|9052/3
C0862312|T191|SY|CDR0000039969|PDQ|Malignant Epithelial Mesothelioma|9052/3
C0862312|T191|SY|CDR0000039969|PDQ|mesothelioma, epithelial|9052/3
C0862312|T191|SY|BBP3.|RCD|Epithelioid mesothelioma|9052/3
C0862312|T191|OA|BBP5.|RCD|Malig epithelioid mesothelioma|9052/3
C0862312|T191|OP|BBP5.|RCD|Malignant epithelioid mesothelioma|9052/3
C0862312|T191|SY|65278006|SNOMEDCT_US|Epithelioid mesothelioma|9052/3
C0862312|T191|PT|65278006|SNOMEDCT_US|Epithelioid mesothelioma, malignant|9052/3
C0862312|T191|IS|65278006|SNOMEDCT_US|Epithelioid mesothelioma, NOS|9052/3
C0862312|T191|SY|65278006|SNOMEDCT_US|Malignant epithelioid mesothelioma|9052/3
C0334515|T191|PT|MTHU010710|ICPC2ICD10ENG|biphasic; mesothelioma|9053/3
C0334515|T191|PT|MTHU048938|ICPC2ICD10ENG|mesothelioma; biphasic|9053/3
C0334515|T191|LLT|10073062|MDR|Biphasic mesothelioma|9053/3
C0334515|T191|PT|10073062|MDR|Biphasic mesothelioma|9053/3
C0334515|T191|PT|C4282|NCI|Biphasic Mesothelioma|9053/3
C0334515|T191|SY|C4282|NCI|Malignant Biphasic Mesothelioma|9053/3
C0334515|T191|SY|C4282|NCI|Malignant Mixed Mesothelioma|9053/3
C0334515|T191|SY|C4282|NCI|Mixed Mesothelioma|9053/3
C0334515|T191|SY|BBP7.|RCD|Biphasic mesothelioma|9053/3
C0334515|T191|AB|BBP7.|RCD|Malign biphasic mesothelioma|9053/3
C0334515|T191|PT|BBP7.|RCD|Malignant biphasic mesothelioma|9053/3
C0334515|T191|SY|30383009|SNOMEDCT_US|Biphasic mesothelioma|9053/3
C0334515|T191|SY|30383009|SNOMEDCT_US|Malignant biphasic mesothelioma|9053/3
C0334515|T191|SY|30383009|SNOMEDCT_US|Mesothelioma, biphasic|9053/3
C0334515|T191|PT|30383009|SNOMEDCT_US|Mesothelioma, biphasic, malignant|9053/3
C0334515|T191|IS|30383009|SNOMEDCT_US|Mesothelioma, biphasic, NOS|9053/3
C0206675|T191|NP|0000023024|AOD|adenomatoid tumor|9054/0
C0206675|T191|PT|0000021013|CHV|adenomatoid tumor|9054/0
C0206675|T191|SY|0000021013|CHV|adenomatoid tumors|9054/0
C0206675|T191|ET|D19.9|ICD10CM|Benign mesothelioma NOS|9054/0
C0206675|T191|LLT|10061691|MDR|Benign mesothelioma|9054/0
C0206675|T191|PT|10061691|MDR|Benign mesothelioma|9054/0
C0206675|T191|LLT|10004291|MDR|Benign mesothelioma NOS|9054/0
C0206675|T191|HT|10027413|MDR|Mesotheliomas benign|9054/0
C0206675|T191|MH|D018254|MSH|Adenomatoid Tumor|9054/0
C0206675|T191|PM|D018254|MSH|Adenomatoid Tumors|9054/0
C0206675|T191|PM|D018254|MSH|Tumor, Adenomatoid|9054/0
C0206675|T191|PM|D018254|MSH|Tumors, Adenomatoid|9054/0
C0206675|T191|PT|C3762|NCI|Adenomatoid Tumor|9054/0
C0206675|T191|SY|C3762|NCI|Benign Localized Epithelial Mesothelioma|9054/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelial Neoplasm|9054/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelial Tumor|9054/0
C0206675|T191|SY|C3762|NCI|Benign Mesothelioma|9054/0
C0206675|T191|SY|C3762|NCI|Benign Neoplasm of Mesothelium|9054/0
C0206675|T191|SY|C3762|NCI|Benign Neoplasm of the Mesothelium|9054/0
C0206675|T191|SY|C3762|NCI|Benign Tumor of Mesothelium|9054/0
C0206675|T191|SY|C3762|NCI|Benign Tumor of the Mesothelium|9054/0
C0206675|T191|SY|C3762|NCI|Mesothelioma, Benign|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Adenomatoid Tumor, Benign|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Localized Epithelial Mesothelioma|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelial Neoplasm|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelial Tumor|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Mesothelioma|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Neoplasm of Mesothelium|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Neoplasm of the Mesothelium|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Tumor of Mesothelium|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Benign Tumor of the Mesothelium|9054/0
C0206675|T191|PT|C3762|NCI_CDISC|MESOTHELIOMA, BENIGN|9054/0
C0206675|T191|SY|C3762|NCI_CDISC|Mesothelioma, Benign|9054/0
C0206675|T191|PT|Xa9AD|RCD|Adenomatoid tumour|9054/0
C0206675|T191|PT|BBP0.|RCD|Benign mesothelioma|9054/0
C0206675|T191|PT|Xa9AD|RCDAE|Adenomatoid tumor|9054/0
C0206675|T191|OP|BBP8.|RCDSA|Adenomatoid tumor NOS|9054/0
C0206675|T191|OP|BBP8.|RCDSY|Adenomatoid tumour NOS|9054/0
C0206675|T191|PT|2348006|SNOMEDCT_US|Adenomatoid tumor|9054/0
C0206675|T191|IS|2348006|SNOMEDCT_US|Adenomatoid tumor, NOS|9054/0
C0206675|T191|PTGB|2348006|SNOMEDCT_US|Adenomatoid tumour|9054/0
C0206675|T191|SY|41183007|SNOMEDCT_US|Benign mesothelioma|9054/0
C0206675|T191|PT|41183007|SNOMEDCT_US|Mesothelioma, benign|9054/0
C0206680|T191|PT|MTHU020774|ICPC2ICD10ENG|cystic; mesothelioma|9055/0
C0206680|T191|PT|MTHU048946|ICPC2ICD10ENG|mesothelioma; cystic|9055/0
C0206680|T191|PM|D018261|MSH|Cystic Mesothelioma|9055/0
C0206680|T191|PM|D018261|MSH|Cystic Mesotheliomas|9055/0
C0206680|T191|MH|D018261|MSH|Mesothelioma, Cystic|9055/0
C0206680|T191|PM|D018261|MSH|Mesotheliomas, Cystic|9055/0
C0206680|T191|SY|C3765|NCI|Cystic Mesothelioma|9055/0
C0206680|T191|SY|C3765|NCI|Intermediate Mesothelioma|9055/0
C0206680|T191|PT|C3765|NCI|Multicystic Mesothelioma|9055/0
C0206680|T191|PT|X77ov|RCD|Cystic mesothelioma|9055/0
C0206680|T191|OAP|189836009|SNOMEDCT_US|Cystic mesothelioma|9055/0
C0206680|T191|OF|189836009|SNOMEDCT_US|Cystic mesothelioma|9055/0
C0206680|T191|PT|86562005|SNOMEDCT_US|Cystic mesothelioma|9055/0
C1266156|T191|SY|128901009|SNOMEDCT_US|Cystic mesothelioma, benign|9055/0
C1266156|T191|PT|128901009|SNOMEDCT_US|Multicystic mesothelioma, benign|9055/0
C0206680|T191|PT|MTHU020774|ICPC2ICD10ENG|cystic; mesothelioma|9055/1
C0206680|T191|PT|MTHU048946|ICPC2ICD10ENG|mesothelioma; cystic|9055/1
C0206680|T191|PM|D018261|MSH|Cystic Mesothelioma|9055/1
C0206680|T191|PM|D018261|MSH|Cystic Mesotheliomas|9055/1
C0206680|T191|MH|D018261|MSH|Mesothelioma, Cystic|9055/1
C0206680|T191|PM|D018261|MSH|Mesotheliomas, Cystic|9055/1
C0206680|T191|SY|C3765|NCI|Cystic Mesothelioma|9055/1
C0206680|T191|SY|C3765|NCI|Intermediate Mesothelioma|9055/1
C0206680|T191|PT|C3765|NCI|Multicystic Mesothelioma|9055/1
C0206680|T191|PT|X77ov|RCD|Cystic mesothelioma|9055/1
C0206680|T191|OF|189836009|SNOMEDCT_US|Cystic mesothelioma|9055/1
C0206680|T191|PT|86562005|SNOMEDCT_US|Cystic mesothelioma|9055/1
C0206680|T191|OAP|189836009|SNOMEDCT_US|Cystic mesothelioma|9055/1
C0013377|T191|SY|0000004207|CHV|disgerminoma|9060/3
C0013377|T191|PT|0000004207|CHV|dysgerminoma|9060/3
C0013377|T191|SY|0000004207|CHV|dysgerminomas|9060/3
C0013377|T191|ET|2016-0850|CSP|dysgerminoma|9060/3
C0013377|T191|PT|HP:0100621|HPO|Dysgerminoma|9060/3
C0013377|T191|PT|sh85038423|LCH_NW|Disgerminoma|9060/3
C0013377|T191|PT|271542|MEDCIN|dysgerminoma|9060/3
C0013377|T191|ET|D004407|MSH|Disgerminoma|9060/3
C0013377|T191|PM|D004407|MSH|Disgerminomas|9060/3
C0013377|T191|MH|D004407|MSH|Dysgerminoma|9060/3
C0013377|T191|PM|D004407|MSH|Dysgerminomas|9060/3
C0013377|T191|PT|C2996|NCI|Dysgerminoma|9060/3
C0013377|T191|PT|C2996|NCI_CDISC|DYSGERMINOMA, MALIGNANT|9060/3
C0013377|T191|PT|C2996|NCI_CPTAC|Dysgerminoma|9060/3
C0013377|T191|PT|C2996|NCI_CTRP|Dysgerminoma|9060/3
C0013377|T191|DN|C2996|NCI_CTRP|Dysgerminoma|9060/3
C0013377|T191|PT|CDR0000672835|NCI_NCI-GLOSS|dysgerminoma|9060/3
C0013377|T191|PT|C2996|NCI_NICHD|Dysgerminoma|9060/3
C0013377|T191|PT|BBQ0.|RCD|Dysgerminoma|9060/3
C0013377|T191|PT|60718004|SNOMEDCT_US|Dysgerminoma|9060/3
C0036631|T191|PT|0019989|CCPSS|SEMINOMA|9061/3
C0036631|T191|PT|0000011191|CHV|seminoma|9061/3
C0036631|T191|SY|0000011191|CHV|seminoma testicular cancer|9061/3
C0036631|T191|SY|0000011191|CHV|seminoma testis|9061/3
C0036631|T191|SY|0000011191|CHV|seminomas|9061/3
C0036631|T191|SY|0000011191|CHV|testicular seminoma|9061/3
C0036631|T191|PT|NOCODE|COSTAR|Seminoma|9061/3
C0036631|T191|PT|U000612|COSTAR|SEMINOMA OF TESTIS|9061/3
C0036631|T191|ET|2016-0850|CSP|seminoma|9061/3
C0036631|T191|GT|CARCINOMA|CST|SEMINOMA|9061/3
C0036631|T191|DI|U001835|DXP|TESTIS, SEMINOMA|9061/3
C0036631|T191|PT|HP:0100617|HPO|Testicular seminoma|9061/3
C0036631|T191|PT|Y78003|ICPC2P|Seminoma|9061/3
C0036631|T191|PTN|Y78003|ICPC2P|seminoma|9061/3
C0036631|T191|PT|10039956|MDR|Seminoma|9061/3
C0036631|T191|LLT|10039956|MDR|Seminoma|9061/3
C0036631|T191|LLT|10043353|MDR|Testicular seminoma pure NOS|9061/3
C0036631|T191|SY|339901|MEDCIN|malignant neoplasm seminoma|9061/3
C0036631|T191|PT|339901|MEDCIN|seminoma|9061/3
C0036631|T191|PT|31522|MEDCIN|seminoma of testis|9061/3
C0036631|T191|SY|31522|MEDCIN|testicular seminoma|9061/3
C0036631|T191|ET|434|MEDLINEPLUS|Seminoma|9061/3
C0036631|T191|MH|D018239|MSH|Seminoma|9061/3
C0036631|T191|PM|D018239|MSH|Seminomas|9061/3
C0036631|T191|PT|C9309|NCI|Seminoma|9061/3
C0036631|T191|SY|C7328|NCI|Seminoma of Testis|9061/3
C0036631|T191|SY|C7328|NCI|Seminoma of the Testis|9061/3
C0036631|T191|SY|C9309|NCI|Seminoma, Pure|9061/3
C0036631|T191|PT|C7328|NCI|Testicular Seminoma|9061/3
C0036631|T191|SY|C7328|NCI|Testicular Seminoma Pure|9061/3
C0036631|T191|SY|C9309|NCI_CDISC|Seminoma|9061/3
C0036631|T191|PT|C9309|NCI_CDISC|SEMINOMA, MALIGNANT|9061/3
C0036631|T191|SY|C9309|NCI_CDISC|Seminoma, Pure|9061/3
C0036631|T191|PT|C9309|NCI_CPTAC|Seminoma|9061/3
C0036631|T191|PT|10043353|NCI_CTEP-SDC|Testicular seminoma|9061/3
C0036631|T191|DN|C9309|NCI_CTRP|Seminoma|9061/3
C0036631|T191|PT|C9309|NCI_CTRP|Seminoma|9061/3
C0036631|T191|PT|C7328|NCI_CTRP|Testicular Seminoma|9061/3
C0036631|T191|DN|C7328|NCI_CTRP|Testicular Seminoma|9061/3
C0036631|T191|PT|CDR0000046577|NCI_NCI-GLOSS|seminoma|9061/3
C0036631|T191|PT|C9309|NCI_NICHD|Seminoma|9061/3
C0036631|T191|SY|CDR0000040003|PDQ|Seminoma of Testis|9061/3
C0036631|T191|SY|CDR0000040003|PDQ|seminoma of the testis|9061/3
C0036631|T191|SY|CDR0000040003|PDQ|seminoma, testicular|9061/3
C0036631|T191|SY|CDR0000040003|PDQ|testicle cancer, seminoma|9061/3
C0036631|T191|SY|CDR0000040003|PDQ|testicular cancer, seminoma|9061/3
C0036631|T191|PT|CDR0000040003|PDQ|testicular seminoma|9061/3
C0036631|T191|SY|CDR0000040003|PDQ|Testicular Seminoma Pure|9061/3
C0036631|T191|SY|CDR0000040003|PDQ|testis cancer, seminoma|9061/3
C0036631|T191|PT|R0121921|QMR|TESTICULAR SEMINOMA|9061/3
C0036631|T191|PT|Xa9AF|RCD|Seminoma|9061/3
C0036631|T191|PT|X78ip|RCD|Seminoma of testis|9061/3
C0036631|T191|OP|BBQ1z|RCDSY|Seminoma NOS|9061/3
C0036631|T191|OP|BBQ1.|RCDSY|Seminomas|9061/3
C4304144|T191|PT|720346009|SNOMEDCT_US|Primary seminoma|9061/3
C0036631|T191|PT|36741007|SNOMEDCT_US|Seminoma|9061/3
C0036631|T191|PT|443675005|SNOMEDCT_US|Seminoma|9061/3
C0036631|T191|PT|255107005|SNOMEDCT_US|Seminoma of testis|9061/3
C0036631|T191|OAS|188228003|SNOMEDCT_US|Seminoma of testis|9061/3
C0036631|T191|OAS|269603004|SNOMEDCT_US|Seminoma of testis|9061/3
C0036631|T191|OAS|154532006|SNOMEDCT_US|Seminoma of testis|9061/3
C0036631|T191|OAS|154532006|SNOMEDCT_US|Seminoma testis|9061/3
C0036631|T191|OAS|269603004|SNOMEDCT_US|Seminoma testis|9061/3
C0036631|T191|SY|36741007|SNOMEDCT_US|Seminoma, no ICD-O subtype|9061/3
C0036631|T191|SY|36741007|SNOMEDCT_US|Seminoma, no International Classification of Diseases for Oncology subtype|9061/3
C0036631|T191|IS|36741007|SNOMEDCT_US|Seminoma, NOS|9061/3
C0036631|T191|PT|1323|WHO|SEMINOMA|9061/3
C0334516|T191|SY|C39920|NCI|Anaplastic Seminoma|9062/3
C0334516|T191|SY|C39920|NCI|Atypical Seminoma|9062/3
C0334516|T191|PT|C39920|NCI|Testicular Seminoma with High Mitotic Index|9062/3
C0334516|T191|PT|BBQ10|RCD|Anaplastic seminoma|9062/3
C0334516|T191|SY|72907003|SNOMEDCT_US|Anaplastic seminoma|9062/3
C0334516|T191|SY|72907003|SNOMEDCT_US|Seminoma with high mitotic index|9062/3
C0334516|T191|PT|72907003|SNOMEDCT_US|Seminoma, anaplastic|9062/3
C0334517|T191|PT|10073118|MDR|Spermatocytic seminoma|9063/3
C0334517|T191|LLT|10073118|MDR|Spermatocytic seminoma|9063/3
C0334517|T191|OP|C39921|NCI|Spermatocytic Seminoma|9063/3
C0334517|T191|SY|C39921|NCI|Spermatocytic Tumor|9063/3
C0334517|T191|OP|C39921|NCI|Testicular Spermatocytic Seminoma|9063/3
C0334517|T191|PT|C39921|NCI|Testicular Spermatocytic Tumor|9063/3
C0334517|T191|PT|BBQ11|RCD|Spermatocytic seminoma|9063/3
C0334517|T191|SY|BBQ11|RCD|Spermatocytoma|9063/3
C0334517|T191|PT|9294008|SNOMEDCT_US|Spermatocytic seminoma|9063/3
C1302371|T191|PT|399399005|SNOMEDCT_US|Spermatocytic seminoma with sarcomatous component|9063/3
C0334517|T191|SY|9294008|SNOMEDCT_US|Spermatocytoma|9063/3
C1515286|T191|AB|C40345|NCI|GCNIS|9064/2
C1515286|T191|SY|C40345|NCI|Gonocytoma In Situ|9064/2
C1515286|T191|AB|C40345|NCI|IGCNU|9064/2
C1515286|T191|PT|C40345|NCI|Testicular Germ Cell Neoplasia In Situ|9064/2
C1515286|T191|SY|C40345|NCI|Testicular Intraepithelial Neoplasia|9064/2
C1515286|T191|SY|C40345|NCI|Testicular Intratubular Germ Cell Neoplasia of the Unclassified Type|9064/2
C1515286|T191|SY|C40345|NCI|Testicular Intratubular Germ Cell Neoplasia of Unclassified Type|9064/2
C1515286|T191|SY|C40345|NCI|Testicular Intratubular Germ Cell Neoplasia, Unclassified|9064/2
C1515286|T191|DN|C40345|NCI_CTRP|Testicular Intratubular Germ Cell Neoplasia, Unclassified|9064/2
C1266157|T191|SY|128902002|SNOMEDCT_US|Intratubular germ cell neoplasia|9064/2
C1266157|T191|PT|128902002|SNOMEDCT_US|Intratubular malignant germ cells|9064/2
C0206660|T191|PT|0000021003|CHV|germinoma|9064/3
C0206660|T191|PT|0000058162|CHV|germinoma|9064/3
C0206660|T191|SY|0000021003|CHV|germinomas|9064/3
C0206660|T191|PT|HP:0100620|HPO|Germinoma|9064/3
C0206660|T191|LLT|10018207|MDR|Germinoma|9064/3
C0206660|T191|PT|271541|MEDCIN|germinoma|9064/3
C0206660|T191|MH|D018237|MSH|Germinoma|9064/3
C0206660|T191|PM|D018237|MSH|Germinomas|9064/3
C0206660|T191|PN|NOCODE|MTH|Germinoma|9064/3
C1275403|T191|SY|C162139|NCI|Burnt-Out Germ Cell Tumor|9064/3
C0206660|T191|SY|TCGA|NCI|Germinoma|9064/3
C0206660|T191|PT|C3753|NCI|Germinoma|9064/3
C1275403|T191|PT|C162139|NCI|Regressed Testicular Germ Cell Tumor|9064/3
C0206660|T191|PT|C3753|NCI_CPTAC|Germinoma|9064/3
C0206660|T191|DN|C3753|NCI_CTRP|Germinoma|9064/3
C0206660|T191|PT|C3753|NCI_CTRP|Germinoma|9064/3
C0206660|T191|PT|C3753|NCI_NICHD|Germinoma|9064/3
C0206660|T191|PT|BBQ2.|RCD|Germinoma|9064/3
C1275403|T191|SY|399523002|SNOMEDCT_US|Burnt out germ cell tumor|9064/3
C1275403|T191|SYGB|399523002|SNOMEDCT_US|Burnt out germ cell tumour|9064/3
C0206660|T191|PT|28307001|SNOMEDCT_US|Germinoma|9064/3
C0206660|T191|OAP|154603000|SNOMEDCT_US|Germinoma|9064/3
C0206660|T191|OF|154603000|SNOMEDCT_US|Germinoma|9064/3
C1275403|T191|PT|399523002|SNOMEDCT_US|Regressed germ cell tumor|9064/3
C1275403|T191|PTGB|399523002|SNOMEDCT_US|Regressed germ cell tumour|9064/3
C1266158|T191|SY|271543|MEDCIN|nonseminomatous germ cell tumor|9065/3
C1266158|T191|PT|271543|MEDCIN|nonseminomatous germinoma|9065/3
C1266158|T191|CE|C537844|MSH|Non-seminomatous germ-cell tumors|9065/3
C1266158|T191|NM|C537844|MSH|Nonseminomatous germ cell tumor|9065/3
C1266158|T191|CE|C537844|MSH|NSGCT Nonseminomatous germ cell tumor|9065/3
C1266158|T191|PN|NOCODE|MTH|Nongerminomatous Germ Cell Tumor|9065/3
C1266158|T191|PT|C121619|NCI|Nongerminomatous Germ Cell Tumor|9065/3
C1266158|T191|SY|C121619|NCI|Nongerminomatous Germ Cell Tumor Including Central Nervous System|9065/3
C1336724|T191|SY|C9313|NCI|Testicular Germ Cell Tumor Non-Seminomatous|9065/3
C1336724|T191|PT|C9313|NCI|Testicular Non-Seminomatous Germ Cell Tumor|9065/3
C1336724|T191|DN|C9313|NCI_CTRP|Testicular Non-Seminomatous Germ Cell Tumor|9065/3
C1266158|T191|SY|C121619|NCI_NICHD|Non-dysgerminomatous Germ Cell Tumor|9065/3
C1266158|T191|SY|C121619|NCI_NICHD|Non-germinomatous Germ Cell Tumor|9065/3
C1266158|T191|SY|C121619|NCI_NICHD|Non-seminomatous Germ Cell Tumor|9065/3
C1266158|T191|PT|C121619|NCI_NICHD|Nongerminomatous Germ Cell Tumor|9065/3
C1266158|T191|PT|128766005|SNOMEDCT_US|Germ cell tumor, nonseminomatous|9065/3
C1266158|T191|PTGB|128766005|SNOMEDCT_US|Germ cell tumour, nonseminomatous|9065/3
C0206659|T191|PT|0000021002|CHV|embryonal carcinoma|9070/3
C0206659|T191|ET|2016-0850|CSP|embryonal carcinoma|9070/3
C0206659|T191|PT|271452|MEDCIN|embryonal carcinoma|9070/3
C0206659|T191|MH|D018236|MSH|Carcinoma, Embryonal|9070/3
C0206659|T191|PM|D018236|MSH|Carcinomas, Embryonal|9070/3
C0206659|T191|PM|D018236|MSH|Embryonal Carcinoma|9070/3
C0206659|T191|PM|D018236|MSH|Embryonal Carcinomas|9070/3
C0206659|T191|PN|NOCODE|MTH|Embryonal Carcinoma|9070/3
C0206659|T191|SY|TCGA|NCI|Embryonal Carcinoma|9070/3
C0206659|T191|PT|C3752|NCI|Embryonal Carcinoma|9070/3
C0206659|T191|PT|C3752|NCI_CDISC|CARCINOMA, EMBRYONAL, MALIGNANT|9070/3
C0206659|T191|SY|C3752|NCI_CDISC|Carcinoma, Embryonal, Malignant|9070/3
C0206659|T191|PT|C3752|NCI_CPTAC|Embryonal Carcinoma|9070/3
C0206659|T191|PT|C3752|NCI_CTRP|Embryonal Carcinoma|9070/3
C0206659|T191|DN|C3752|NCI_CTRP|Embryonal Carcinoma|9070/3
C0206659|T191|SY|Xa9AG|RCD|Embryonal adenocarcinoma|9070/3
C0206659|T191|PT|Xa9AG|RCD|Embryonal carcinoma|9070/3
C0206659|T191|OP|BBQ3.|RCDSY|Embryonal carcinoma NOS|9070/3
C0206659|T191|SY|28047004|SNOMEDCT_US|Embryonal adenocarcinoma|9070/3
C0206659|T191|PT|28047004|SNOMEDCT_US|Embryonal carcinoma|9070/3
C0206659|T191|IS|28047004|SNOMEDCT_US|Embryonal carcinoma, NOS|9070/3
C0014145|T191|SY|0000004455|CHV|endodermal sinus tumor|9071/3
C0014145|T191|SY|0000004455|CHV|endodermal sinus tumour|9071/3
C0014145|T191|SY|0000004455|CHV|orchioblastoma|9071/3
C0014145|T191|PT|0000004455|CHV|yolk sac tumor|9071/3
C0014145|T191|PT|MTHU055870|ICPC2ICD10ENG|orchioblastoma|9071/3
C0014145|T191|LLT|10062419|MDR|Endodermal sinus tumor site unspecified|9071/3
C0014145|T191|LLT|10014718|MDR|Endodermal sinus tumour site unspecified|9071/3
C0014145|T191|MTH_LLT|10048251|MDR|Yolk sac tumor site unspecified|9071/3
C0014145|T191|MTH_PT|10048251|MDR|Yolk sac tumor site unspecified|9071/3
C0014145|T191|LLT|10048251|MDR|Yolk sac tumour site unspecified|9071/3
C0014145|T191|PT|10048251|MDR|Yolk sac tumour site unspecified|9071/3
C0014145|T191|PT|271453|MEDCIN|yolk sac tumor|9071/3
C0014145|T191|MH|D018240|MSH|Endodermal Sinus Tumor|9071/3
C0014145|T191|PM|D018240|MSH|Endodermal Sinus Tumors|9071/3
C0014145|T191|PM|D018240|MSH|Tumor, Endodermal Sinus|9071/3
C0014145|T191|PM|D018240|MSH|Tumor, Yolk Sac|9071/3
C0014145|T191|PM|D018240|MSH|Tumors, Endodermal Sinus|9071/3
C0014145|T191|PM|D018240|MSH|Tumors, Yolk Sac|9071/3
C0014145|T191|ET|D018240|MSH|Yolk Sac Tumor|9071/3
C0014145|T191|PM|D018240|MSH|Yolk Sac Tumors|9071/3
C0014145|T191|PN|NOCODE|MTH|Yolk Sac Tumor|9071/3
C0014145|T191|SY|C3011|NCI|Endodermal Sinus Neoplasm|9071/3
C0014145|T191|SY|C3011|NCI|Endodermal Sinus Tumor|9071/3
C0014145|T191|SY|C3011|NCI|Yolk Sac Neoplasm|9071/3
C0014145|T191|PT|C3011|NCI|Yolk Sac Tumor|9071/3
C0014145|T191|SY|TCGA|NCI|Yolk Sac Tumor|9071/3
C0014145|T191|SY|C3011|NCI|Yolk Sac Tumour Site Unspecified|9071/3
C0014145|T191|SY|C3011|NCI_CDISC|Carcinoma, Yolk Sac|9071/3
C0014145|T191|SY|C3011|NCI_CDISC|Endodermal Sinus Neoplasm|9071/3
C0014145|T191|SY|C3011|NCI_CDISC|Endodermal Sinus Tumor|9071/3
C0014145|T191|SY|C3011|NCI_CDISC|Yolk Sac Neoplasm|9071/3
C0014145|T191|SY|C3011|NCI_CDISC|Yolk Sac Tumor Site Unspecified|9071/3
C0014145|T191|PT|C3011|NCI_CDISC|YOLK SAC TUMOR, MALIGNANT|9071/3
C0014145|T191|PT|C3011|NCI_CPTAC|Yolk Sac Tumor|9071/3
C0014145|T191|PT|C3011|NCI_CTRP|Yolk Sac Tumor|9071/3
C0014145|T191|DN|C3011|NCI_CTRP|Yolk Sac Tumor|9071/3
C0014145|T191|PT|BBQ4.|RCD|Endodermal sinus tumour|9071/3
C0014145|T191|SY|BBQ4.|RCD|Infantile embryonal carcinoma|9071/3
C0014145|T191|SY|BBQ4.|RCD|Orchioblastoma|9071/3
C0014145|T191|SY|BBQ4.|RCD|Polyvesicular vitelline tumour|9071/3
C0014145|T191|SY|BBQ4.|RCD|Yolk sac tumour|9071/3
C0014145|T191|PT|BBQ4.|RCDAE|Endodermal sinus tumor|9071/3
C0014145|T191|SY|BBQ4.|RCDAE|Polyvesicular vitelline tumor|9071/3
C0014145|T191|SY|BBQ4.|RCDAE|Yolk sac tumor|9071/3
C0014145|T191|SY|74409009|SNOMEDCT_US|Embryonal carcinoma, infantile|9071/3
C0014145|T191|PT|74409009|SNOMEDCT_US|Endodermal sinus tumor|9071/3
C0014145|T191|PTGB|74409009|SNOMEDCT_US|Endodermal sinus tumour|9071/3
C0014145|T191|SY|74409009|SNOMEDCT_US|Hepatoid yolk sac tumor|9071/3
C0014145|T191|SYGB|74409009|SNOMEDCT_US|Hepatoid yolk sac tumour|9071/3
C0014145|T191|SY|74409009|SNOMEDCT_US|Infantile embryonal carcinoma|9071/3
C0014145|T191|SY|74409009|SNOMEDCT_US|Orchioblastoma|9071/3
C0014145|T191|SY|74409009|SNOMEDCT_US|Polyvesicular vitelline tumor|9071/3
C0014145|T191|SYGB|74409009|SNOMEDCT_US|Polyvesicular vitelline tumour|9071/3
C0014145|T191|PT|404081005|SNOMEDCT_US|Yolk sac tumor|9071/3
C0014145|T191|SY|74409009|SNOMEDCT_US|Yolk sac tumor|9071/3
C0014145|T191|PTGB|404081005|SNOMEDCT_US|Yolk sac tumour|9071/3
C0014145|T191|SYGB|74409009|SNOMEDCT_US|Yolk sac tumour|9071/3
C0334518|T191|PT|271454|MEDCIN|polyembryoma|9072/3
C1880996|T191|PT|C66776|NCI|Gonadal Polyembryoma|9072/3
C1880996|T191|DN|C66776|NCI_CTRP|Gonadal Polyembryoma|9072/3
C0334518|T191|AB|BBQ5.|RCD|Embryonal ca - polyembryonal|9072/3
C0334518|T191|SY|BBQ5.|RCD|Embryonal carcinoma - polyembryonal type|9072/3
C0334518|T191|PT|BBQ5.|RCD|Polyembryoma|9072/3
C0334518|T191|SY|28325008|SNOMEDCT_US|Embryonal carcinoma - polyembryonal type|9072/3
C0334518|T191|SY|28325008|SNOMEDCT_US|Embryonal carcinoma, polyembryonal type|9072/3
C0334518|T191|PT|28325008|SNOMEDCT_US|Polyembryoma|9072/3
C0206661|T191|PT|0000021004|CHV|gonadoblastoma|9073/1
C0206661|T191|SY|0000021004|CHV|gonadoblastomas|9073/1
C0206661|T191|ET|2016-0850|CSP|gonadoblastoma|9073/1
C0206661|T191|PT|HP:0000150|HPO|Gonadoblastoma|9073/1
C0206661|T191|LLT|10018506|MDR|Gonadoblastoma|9073/1
C0206661|T191|MH|D018238|MSH|Gonadoblastoma|9073/1
C0206661|T191|PM|D018238|MSH|Gonadoblastomas|9073/1
C0206661|T191|PT|C3754|NCI|Gonadoblastoma|9073/1
C0206661|T191|PT|C3754|NCI_NICHD|Gonadoblastoma|9073/1
C0206661|T191|SY|BBQ6.|RCD|GBY - Gonadoblastoma|9073/1
C0206661|T191|PT|BBQ6.|RCD|Gonadoblastoma|9073/1
C0206661|T191|SY|BBQ6.|RCD|Gonocytoma|9073/1
C0206661|T191|SY|74751003|SNOMEDCT_US|GBY - Gonadoblastoma|9073/1
C0206661|T191|PT|74751003|SNOMEDCT_US|Gonadoblastoma|9073/1
C0206661|T191|SY|74751003|SNOMEDCT_US|Gonocytoma|9073/1
C1321219|T191|PT|406095005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumor, gonadoblastoma|9073/1
C1321219|T191|PTGB|406095005|SNOMEDCT_US|Mixed germ cell-sex cord-stromal tumour, gonadoblastoma|9073/1
C1879828|T191|PT|0012271|CCPSS|TERATOMA BENIGN|9080/0
C1368910|T191|PT|1009546|CCPSS|TERATOMA MATURE CYSTIC|9080/0
C1879828|T191|ET|D28|ICD10CM|benign teratoma|9080/0
C1879828|T191|LLT|10048460|MDR|Teratoma benign|9080/0
C1879828|T191|PT|10048460|MDR|Teratoma benign|9080/0
C1879828|T191|PM|D013724|MSH|Benign Teratoma|9080/0
C1879828|T191|PM|D013724|MSH|Benign Teratomas|9080/0
C1879828|T191|PEP|D013724|MSH|Teratoma, Benign|9080/0
C1879828|T191|ET|D013724|MSH|Teratoma, Cystic|9080/0
C1879828|T191|ET|D013724|MSH|Teratoma, Mature|9080/0
C1879828|T191|PM|D013724|MSH|Teratomas, Benign|9080/0
C1879828|T191|PN|NOCODE|MTH|Benign Teratoma|9080/0
C1368910|T191|PN|NOCODE|MTH|Mature Teratoma|9080/0
C1879828|T191|PT|C67107|NCI|Benign Teratoma|9080/0
C1368910|T191|SY|C9015|NCI|Grade 0 Teratoma|9080/0
C1368910|T191|PT|C9015|NCI|Mature Teratoma|9080/0
C1368910|T191|SY|TCGA|NCI|Mature Teratoma|9080/0
C1879828|T191|DN|C67107|NCI_CTRP|Benign Teratoma|9080/0
C1368910|T191|PT|CDR0000443575|NCI_NCI-GLOSS|mature teratoma|9080/0
C1879828|T191|PT|CDR0000561977|PDQ|benign teratoma|9080/0
C1879828|T191|SY|BBQ8.|RCD|Benign teratoma|9080/0
C1879828|T191|SY|BBQ8.|RCD|Cystic teratoma|9080/0
C1879828|T191|SY|BBQ8.|RCD|Differentiated teratoma|9080/0
C1368910|T191|SY|BBQ8.|RCD|Mature teratoma|9080/0
C1879828|T191|SY|42717009|SNOMEDCT_US|Benign teratoma|9080/0
C1879828|T191|SY|42717009|SNOMEDCT_US|Differentiated teratoma|9080/0
C1368910|T191|SY|42717009|SNOMEDCT_US|Mature teratoma|9080/0
C1368910|T191|IS|55818009|SNOMEDCT_US|Mature teratoma|9080/0
C1879828|T191|PT|42717009|SNOMEDCT_US|Teratoma, benign|9080/0
C1879828|T191|OAS|189119004|SNOMEDCT_US|Teratoma, benign|9080/0
C1879828|T191|SY|42717009|SNOMEDCT_US|Teratoma, differentiated|9080/0
C1879828|T191|PT|1823|WHO|TERATOMA BENIGN|9080/0
C0039538|T191|ET|0000004549|AOD|teratoma|9080/1
C0039538|T191|PT|0013786|CCPSS|TERATOMA|9080/1
C0039538|T191|SY|0000012107|CHV|teratoid tumor|9080/1
C0039538|T191|SY|0000012107|CHV|teratoid tumors|9080/1
C0039538|T191|PT|0000012107|CHV|teratoma|9080/1
C0039538|T191|SY|0000012107|CHV|teratomas|9080/1
C0039538|T191|PT|2000-4962|CSP|teratoma|9080/1
C0039538|T191|GT|NEOPL|CST|TERATOMA|9080/1
C0039538|T191|PT|HP:0009792|HPO|Teratoma|9080/1
C0039538|T191|PT|U004617|LCH|Teratoma|9080/1
C0039538|T191|PT|sh85133985|LCH_NW|Teratoma|9080/1
C0039538|T191|LLT|10043276|MDR|Teratoma|9080/1
C0039538|T191|PT|10043276|MDR|Teratoma|9080/1
C0039538|T191|LLT|10043277|MDR|Teratoma NOS|9080/1
C0039538|T191|PT|367879|MEDCIN|teratoma|9080/1
C0039538|T191|ET|D013724|MSH|Dysembryoma|9080/1
C0039538|T191|PM|D013724|MSH|Dysembryomas|9080/1
C0039538|T191|ET|D013724|MSH|Teratoid Tumor|9080/1
C0039538|T191|PM|D013724|MSH|Teratoid Tumors|9080/1
C0039538|T191|MH|D013724|MSH|Teratoma|9080/1
C0039538|T191|PM|D013724|MSH|Teratomas|9080/1
C0039538|T191|PM|D013724|MSH|Tumor, Teratoid|9080/1
C0039538|T191|PM|D013724|MSH|Tumors, Teratoid|9080/1
C0039538|T191|PN|NOCODE|MTH|Teratoma|9080/1
C0039538|T191|PT|C3403|NCI|Teratoma|9080/1
C0039538|T191|PT|C3403|NCI_CPTAC|Teratoma|9080/1
C0039538|T191|PT|C3403|NCI_CTRP|Teratoma|9080/1
C0039538|T191|DN|C3403|NCI_CTRP|Teratoma|9080/1
C0039538|T191|PT|CDR0000044248|NCI_NCI-GLOSS|teratoma|9080/1
C0039538|T191|PT|C3403|NCI_NICHD|Teratoma|9080/1
C0039538|T191|ET|CDR0000553672|PDQ|Teratoma|9080/1
C0039538|T191|PT|CDR0000553672|PDQ|teratoma|9080/1
C0039538|T191|PT|Xa9AH|RCD|Teratoma|9080/1
C0039538|T191|OP|BBQ71|RCDSY|Teratoma NOS|9080/1
C0039538|T191|OP|BBQ7.|RCDSY|Teratomas|9080/1
C0039538|T191|PT|36591000119102|SNOMEDCT_US|Teratoma|9080/1
C0039538|T191|PT|55818009|SNOMEDCT_US|Teratoma|9080/1
C0039538|T191|SY|55818009|SNOMEDCT_US|Teratoma, no ICD-O subtype|9080/1
C0039538|T191|SY|55818009|SNOMEDCT_US|Teratoma, no International Classification of Diseases for Oncology subtype|9080/1
C0039538|T191|IS|55818009|SNOMEDCT_US|Teratoma, NOS|9080/1
C0039538|T191|PT|1186|WHO|TERATOMA|9080/1
C0334520|T191|SY|0000030000|CHV|immature teratoma|9080/3
C0334520|T191|PT|0000030000|CHV|malignant teratoma|9080/3
C0334520|T191|SY|0000030000|CHV|teratoma malignant|9080/3
C0334520|T191|PT|271544|MEDCIN|malignant teratoma|9080/3
C0334520|T191|PM|D013724|MSH|Immature Teratoma|9080/3
C0334520|T191|PM|D013724|MSH|Immature Teratomas|9080/3
C0334520|T191|PM|D013724|MSH|Malignant Teratoma|9080/3
C0334520|T191|PM|D013724|MSH|Malignant Teratomas|9080/3
C0334520|T191|ET|D013724|MSH|Teratoma, Immature|9080/3
C0334520|T191|PEP|D013724|MSH|Teratoma, Malignant|9080/3
C0334520|T191|PM|D013724|MSH|Teratomas, Immature|9080/3
C0334520|T191|PM|D013724|MSH|Teratomas, Malignant|9080/3
C0334520|T191|PN|NOCODE|MTH|Teratoma, Malignant|9080/3
C0334520|T191|SY|C4286|NCI|Grade 2 Teratoma|9080/3
C0334520|T191|PT|C4286|NCI|Immature Teratoma|9080/3
C0334520|T191|SY|TCGA|NCI|Immature Teratoma|9080/3
C1302569|T191|SY|C7286|NCI|Monodermal Teratoma|9080/3
C1302569|T191|PT|C7286|NCI|Ovarian Monodermal Teratoma|9080/3
C0334520|T191|PT|CDR0000443576|NCI_NCI-GLOSS|immature teratoma|9080/3
C0334520|T191|SY|Xa9AI|RCD|Immature teratoma|9080/3
C0334520|T191|SY|Xa9AI|RCD|Malignant teratoblastoma|9080/3
C0334520|T191|PT|Xa9AI|RCD|Malignant teratoma|9080/3
C0334520|T191|SY|Xa9AI|RCDSY|Teratoma, malignant, NOS|9080/3
C0334520|T191|SY|19467007|SNOMEDCT_US|Embryonal teratoma|9080/3
C0334520|T191|IS|19467007|SNOMEDCT_US|Immature teratoma|9080/3
C0334520|T191|IS|19467007|SNOMEDCT_US|Immature teratoma, malignant|9080/3
C0334520|T191|SY|827161000|SNOMEDCT_US|Immature teratoma, malignant|9080/3
C0334520|T191|PT|827161000|SNOMEDCT_US|Malignant immature teratoma|9080/3
C0334520|T191|SY|19467007|SNOMEDCT_US|Malignant teratoblastoma|9080/3
C0334520|T191|OF|189847002|SNOMEDCT_US|Malignant teratoma|9080/3
C0334520|T191|PT|189847002|SNOMEDCT_US|Malignant teratoma|9080/3
C1302569|T191|PT|399632009|SNOMEDCT_US|Monodermal teratoma|9080/3
C4518229|T191|PT|733890000|SNOMEDCT_US|Postpubertal type teratoma|9080/3
C0334520|T191|SY|19467007|SNOMEDCT_US|Teratoblastoma, malignant|9080/3
C0334520|T191|PT|19467007|SNOMEDCT_US|Teratoma, malignant|9080/3
C0334520|T191|SY|19467007|SNOMEDCT_US|Teratoma, malignant, no ICD-O subtype|9080/3
C0334520|T191|SY|19467007|SNOMEDCT_US|Teratoma, malignant, no International Classification of Diseases for Oncology subtype|9080/3
C0334520|T191|IS|19467007|SNOMEDCT_US|Teratoma, malignant, NOS|9080/3
C0206664|T191|PT|0000021006|CHV|teratocarcinoma|9081/3
C0206664|T191|PT|sh85133982|LCH_NW|Teratocarcinoma|9081/3
C0206664|T191|PT|271545|MEDCIN|teratocarcinoma|9081/3
C0206664|T191|MH|D018243|MSH|Teratocarcinoma|9081/3
C0206664|T191|PM|D018243|MSH|Teratocarcinomas|9081/3
C0206664|T191|PT|C3756|NCI|Mixed Embryonal Carcinoma and Teratoma|9081/3
C0206664|T191|SY|C3756|NCI|Teratocarcinoma|9081/3
C0206664|T191|PT|CDR0000446558|NCI_NCI-GLOSS|teratocarcinoma|9081/3
C0206664|T191|AB|BBQ73|RCD|Mixed embryonal ca & teratoma|9081/3
C0206664|T191|SY|BBQ73|RCD|Mixed embryonal carcinoma and teratoma|9081/3
C0206664|T191|PT|BBQ73|RCD|Teratocarcinoma|9081/3
C0206664|T191|SY|67830002|SNOMEDCT_US|Mixed embryonal carcinoma and teratoma|9081/3
C0206664|T191|PT|67830002|SNOMEDCT_US|Teratocarcinoma|9081/3
C0334521|T191|SY|271546|MEDCIN|malignant undifferentiated teratoma|9082/3
C0334521|T191|PT|271546|MEDCIN|undifferentiated malignant teratoma|9082/3
C4722083|T191|PN|NOCODE|MTH|Grade 3 Teratoma|9082/3
C4722083|T191|SY|C4287|NCI|Grade 3 Teratoma|9082/3
C4722083|T191|PT|C4287|NCI|Malignant Teratoma|9082/3
C4722083|T191|PT|C4287|NCI_CDISC|TERATOMA, MALIGNANT|9082/3
C0334521|T191|SY|BBQ74|RCD|Malignant teratoma - anaplastic|9082/3
C0334521|T191|AB|BBQ74|RCD|Malignant teratoma - undiff|9082/3
C0334521|T191|PT|BBQ74|RCD|Malignant teratoma - undifferentiated|9082/3
C0334521|T191|AB|BBQ74|RCD|Malignant teratoma-anaplastic|9082/3
C0334521|T191|SY|83292005|SNOMEDCT_US|Malignant teratoma - anaplastic|9082/3
C0334521|T191|SY|83292005|SNOMEDCT_US|Malignant teratoma - undifferentiated|9082/3
C0334521|T191|SY|83292005|SNOMEDCT_US|Malignant teratoma, anaplastic|9082/3
C0334521|T191|PT|83292005|SNOMEDCT_US|Malignant teratoma, undifferentiated|9082/3
C0334522|T191|PT|271547|MEDCIN|intermediate malignant teratoma|9083/3
C0334522|T191|SY|271547|MEDCIN|malignant intermediate teratoma|9083/3
C0334522|T191|OP|C4288|NCI|Intermediate Immature Teratoma|9083/3
C0334522|T191|PT|C4288|NCI|Intermediate Immature Teratoma|9083/3
C0334522|T191|OP|C4288|NCI|Intermediate Malignant Teratoma|9083/3
C0334522|T191|AB|BBQ75|RCD|Malign teratoma-intermediate|9083/3
C0334522|T191|PT|BBQ75|RCD|Malignant teratoma - intermediate|9083/3
C0334522|T191|SY|21912003|SNOMEDCT_US|Malignant teratoma - intermediate|9083/3
C0334522|T191|PT|21912003|SNOMEDCT_US|Malignant teratoma, intermediate|9083/3
C0011649|T191|PT|1009398|CCPSS|DERMOID CYST|9084/0
C0011649|T191|SY|0000003805|CHV|benign teratoma|9084/0
C0011649|T191|SY|0000003805|CHV|cystic teratoma|9084/0
C0011649|T191|SY|0000003805|CHV|dermoid|9084/0
C0011649|T191|PT|0000003805|CHV|dermoid cyst|9084/0
C0011649|T191|SY|0000003805|CHV|dermoid cysts|9084/0
C0011649|T191|SY|0000003805|CHV|dermoids|9084/0
C0011649|T191|SY|0000003805|CHV|horn cyst|9084/0
C0011649|T191|SY|0000003805|CHV|mature cystic teratoma|9084/0
C0011649|T191|SY|0000003805|CHV|mature teratoma|9084/0
C0011649|T191|PT|NOCODE|COSTAR|Dermoid|9084/0
C0011649|T191|ET|2000-4962|CSP|dermoid cyst|9084/0
C0011649|T191|PT|HP:0025247|HPO|Dermoid cyst|9084/0
C0011649|T191|ET|K09.8|ICD10CM|Dermoid cyst|9084/0
C0011649|T191|PT|S79008|ICPC2P|Cyst;dermoid|9084/0
C0011649|T191|PTN|S79008|ICPC2P|dermoid cyst|9084/0
C0011649|T191|OP|S80002|ICPC2P|Dermoid cyst|9084/0
C0011649|T191|PT|10012522|MDR|Dermoid cyst|9084/0
C0011649|T191|LLT|10012522|MDR|Dermoid cyst|9084/0
C0011649|T191|LLT|10012523|MDR|Dermoid cyst NOS|9084/0
C0011649|T191|PM|D003884|MSH|Cyst, Dermoid|9084/0
C0011649|T191|PM|D003884|MSH|Cysts, Dermoid|9084/0
C0011649|T191|ET|D003884|MSH|Dermoid|9084/0
C0011649|T191|MH|D003884|MSH|Dermoid Cyst|9084/0
C0011649|T191|PM|D003884|MSH|Dermoid Cysts|9084/0
C0011649|T191|PM|D003884|MSH|Dermoids|9084/0
C0011649|T191|PN|NOCODE|MTH|Dermoid Cyst|9084/0
C0011649|T191|SY|C9011|NCI|Benign Cystic Teratoma|9084/0
C0011649|T191|SY|C9011|NCI|Dermoid|9084/0
C0011649|T191|PT|C9011|NCI|Dermoid Cyst|9084/0
C0011649|T191|SY|C9011|NCI|Dermoid Tumor|9084/0
C0011649|T191|SY|C9011|NCI|Mature Cystic Teratoma|9084/0
C0011649|T191|SY|C9011|NCI_CDISC|Benign Cystic Teratoma|9084/0
C0011649|T191|SY|C9011|NCI_CDISC|Dermoid|9084/0
C0011649|T191|PT|C9011|NCI_CDISC|DERMOID CYST, BENIGN|9084/0
C0011649|T191|SY|C9011|NCI_CDISC|Mature Cystic Teratoma|9084/0
C0011649|T191|DN|C9011|NCI_CTRP|Dermoid Cyst|9084/0
C0011649|T191|PT|CDR0000479002|NCI_NCI-GLOSS|dermoid cyst|9084/0
C0011649|T191|PT|C9011|NCI_NICHD|Dermoid Cyst|9084/0
C0011649|T191|SY|C9011|NCI_NICHD|Subcutaneous Cystic Teratoma|9084/0
C0011649|T191|IS|B7A1.|RCD|Dermoid|9084/0
C0011649|T191|OP|B7A1.|RCD|Dermoid cyst|9084/0
C0011649|T191|PT|BBQ8.|RCDSY|Dermoid cyst|9084/0
C0011649|T191|OP|417609007|SNOMEDCT_US|"Dermoid" tumor|9084/0
C0011649|T191|OP|417609007|SNOMEDCT_US|"Dermoid" tumour|9084/0
C0011649|T191|SY|417137001|SNOMEDCT_US|Dermoid|9084/0
C0011649|T191|IS|417609007|SNOMEDCT_US|Dermoid|9084/0
C0011649|T191|OAS|189117002|SNOMEDCT_US|Dermoid|9084/0
C0011649|T191|OAS|419952004|SNOMEDCT_US|Dermoid|9084/0
C0011649|T191|OAS|72277008|SNOMEDCT_US|Dermoid|9084/0
C0011649|T191|OAP|189117002|SNOMEDCT_US|Dermoid cyst|9084/0
C0011649|T191|OAP|419952004|SNOMEDCT_US|Dermoid cyst|9084/0
C0011649|T191|SY|416529009|SNOMEDCT_US|Dermoid cyst|9084/0
C0011649|T191|OAP|72277008|SNOMEDCT_US|Dermoid cyst|9084/0
C0011649|T191|OAS|269641006|SNOMEDCT_US|Dermoid cyst|9084/0
C0011649|T191|PT|123151001|SNOMEDCT_US|Dermoid cyst|9084/0
C0011649|T191|IS|123151001|SNOMEDCT_US|Dermoid cyst -RETIRED-|9084/0
C0011649|T191|OF|123151001|SNOMEDCT_US|Dermoid cyst -RETIRED-|9084/0
C0011649|T191|IS|72277008|SNOMEDCT_US|Dermoid cyst, NOS|9084/0
C0011649|T191|PT|417609007|SNOMEDCT_US|Dermoid tumor|9084/0
C0011649|T191|PTGB|417609007|SNOMEDCT_US|Dermoid tumour|9084/0
C0011649|T191|IS|72277008|SNOMEDCT_US|Dermoid, NOS|9084/0
C0011649|T191|OAS|72277008|SNOMEDCT_US|Mature cystic teratoma|9084/0
C0011649|T191|OAP|439575008|SNOMEDCT_US|Mature cystic teratoma|9084/0
C0011649|T191|IT|1823|WHO|DERMOID CYST|9084/0
C0334523|T191|PT|MTHU022656|ICPC2ICD10ENG|dermoid; cyst, with malignant transformation|9084/3
C0334523|T191|PT|MTHU047315|ICPC2ICD10ENG|malignant; transformation dermoid cyst|9084/3
C0334523|T191|PT|271548|MEDCIN|teratoma with malignant transformation|9084/3
C0334523|T191|SY|C4289|NCI|Dermoid Cyst with Malignant Transformation|9084/3
C0334523|T191|SY|C4289|NCI|Teratoma with Malignant Transformation|9084/3
C0334523|T191|PT|C4289|NCI|Teratoma with Somatic-Type Malignancy|9084/3
C0334523|T191|OP|BBQ9.|RCD|Dermoid cyst with malignant transformation|9084/3
C0334523|T191|OA|BBQ9.|RCD|Dermoid cyst+malign transform|9084/3
C0334523|T191|AB|Xa9AJ|RCD|Teratoma + malignant transform|9084/3
C0334523|T191|PT|Xa9AJ|RCD|Teratoma with malignant transformation|9084/3
C0334523|T191|IS|189849004|SNOMEDCT_US|:: Dermoid cyst with malignant transformation|9084/3
C0334523|T191|SY|88334008|SNOMEDCT_US|Dermoid cyst with malignant transformation|9084/3
C0334523|T191|SY|189849004|SNOMEDCT_US|Dermoid cyst with malignant transformation|9084/3
C0334523|T191|PT|189849004|SNOMEDCT_US|Dermoid cyst with secondary tumor|9084/3
C0334523|T191|SY|88334008|SNOMEDCT_US|Dermoid cyst with secondary tumor|9084/3
C0334523|T191|PTGB|189849004|SNOMEDCT_US|Dermoid cyst with secondary tumour|9084/3
C0334523|T191|SYGB|88334008|SNOMEDCT_US|Dermoid cyst with secondary tumour|9084/3
C4518371|T191|PT|734071003|SNOMEDCT_US|Germ cell neoplasm with somatic-type solid malignancy|9084/3
C0334523|T191|OAP|302854009|SNOMEDCT_US|Teratoma with malignant transformation|9084/3
C0334523|T191|PT|88334008|SNOMEDCT_US|Teratoma with malignant transformation|9084/3
C0334524|T191|PT|MTHU041362|ICPC2ICD10ENG|germ cell; tumor, mixed|9085/3
C0334524|T191|PT|MTHU031212|ICPC2ICD10ENG|mixed; germ cell tumor|9085/3
C0334524|T191|PT|MTHU077077|ICPC2ICD10ENG|tumor; germ cell, mixed|9085/3
C0334524|T191|PT|271549|MEDCIN|mixed germ cell tumor|9085/3
C0334524|T191|PN|NOCODE|MTH|Mixed Germ Cell Tumor|9085/3
C0334524|T191|SY|C4290|NCI|Combined Germ Cell Neoplasm|9085/3
C0334524|T191|SY|C4290|NCI|Combined Germ Cell Tumor|9085/3
C0334524|T191|SY|C4290|NCI|Mixed Germ Cell Neoplasm|9085/3
C0334524|T191|PT|C4290|NCI|Mixed Germ Cell Tumor|9085/3
C0334524|T191|SY|TCGA|NCI|Mixed Germ Cell Tumor|9085/3
C0334524|T191|PT|C9010|NCI|Mixed Teratoma and Seminoma|9085/3
C0334524|T191|PT|C4290|NCI_CPTAC|Mixed Germ Cell Tumor|9085/3
C0334524|T191|PT|C4290|NCI_CTRP|Mixed Germ Cell Tumor|9085/3
C0334524|T191|DN|C4290|NCI_CTRP|Mixed Germ Cell Tumor|9085/3
C0334524|T191|PT|X77ow|RCD|Mixed germ cell tumour|9085/3
C0334524|T191|PT|X77ow|RCDAE|Mixed germ cell tumor|9085/3
C0334524|T191|PT|32844007|SNOMEDCT_US|Mixed germ cell tumor|9085/3
C0334524|T191|OAP|189853002|SNOMEDCT_US|Mixed germ cell tumor|9085/3
C0334524|T191|OAP|189853002|SNOMEDCT_US|Mixed germ cell tumour|9085/3
C0334524|T191|OF|189853002|SNOMEDCT_US|Mixed germ cell tumour|9085/3
C0334524|T191|PTGB|32844007|SNOMEDCT_US|Mixed germ cell tumour|9085/3
C0334524|T191|SY|32844007|SNOMEDCT_US|Mixed teratoma and seminoma|9085/3
C4518245|T191|PT|733918007|SNOMEDCT_US|Prepubertal type mixed teratoma and yolk sac neoplasm|9085/3
C0038478|T191|SY|0000011788|CHV|ovary tumor thyroid|9090/0
C0038478|T191|PT|0000011788|CHV|struma ovarii|9090/0
C0038478|T191|SY|NOCODE|DXP|OVARIAN CANCER, STRUMA OVARII|9090/0
C0038478|T191|SY|NOCODE|DXP|OVARY, THYROID TUMOR|9090/0
C0038478|T191|DI|U001792|DXP|STRUMA OVARII|9090/0
C0038478|T191|PT|MTHU071029|ICPC2ICD10ENG|struma; ovarii|9090/0
C0038478|T191|LLT|10062581|MDR|Struma ovarii|9090/0
C0038478|T191|PT|31615|MEDCIN|benign struma ovarii of ovary|9090/0
C0038478|T191|SY|31615|MEDCIN|struma ovarii|9090/0
C0038478|T191|MH|D013330|MSH|Struma Ovarii|9090/0
C0038478|T191|PN|NOCODE|MTH|Struma Ovarii|9090/0
C0038478|T191|PT|C7468|NCI|Struma Ovarii|9090/0
C0038478|T191|PT|Xa9AK|RCD|Struma ovarii|9090/0
C0038478|T191|OP|BBQA0|RCDSY|Struma ovarii NOS|9090/0
C0038478|T191|PT|24327009|SNOMEDCT_US|Struma ovarii|9090/0
C0038478|T191|IS|24327009|SNOMEDCT_US|Struma ovarii, NOS|9090/0
C0334525|T191|PT|MTHU071030|ICPC2ICD10ENG|struma; ovarii, malignant|9090/3
C0334525|T191|PT|233172|MEDCIN|malignant struma ovarii|9090/3
C0334525|T191|PT|C4291|NCI|Malignant Struma Ovarii|9090/3
C0334525|T191|PT|BBQA1|RCD|Malignant struma ovarii|9090/3
C0334525|T191|SY|18854008|SNOMEDCT_US|Malignant struma ovarii|9090/3
C0334525|T191|PT|18854008|SNOMEDCT_US|Struma ovarii, malignant|9090/3
C0334526|T191|PT|MTHU014704|ICPC2ICD10ENG|carcinoid; strumal|9091/1
C0334526|T191|PT|MTHU014703|ICPC2ICD10ENG|carcinoid; with struma ovarii|9091/1
C0334526|T191|PT|MTHU071049|ICPC2ICD10ENG|struma ovarii; carcinoid|9091/1
C0334526|T191|PT|MTHU071031|ICPC2ICD10ENG|struma; ovarii, with carcinoid|9091/1
C0334526|T191|PT|MTHU070978|ICPC2ICD10ENG|strumal; carcinoid|9091/1
C0334526|T191|SY|C4292|NCI|Struma Ovarii and Carcinoid|9091/1
C0334526|T191|PT|C4292|NCI|Strumal Carcinoid|9091/1
C0334526|T191|SY|BBQA2|RCD|Struma ovarii and carcinoid|9091/1
C0334526|T191|PT|BBQA2|RCD|Strumal carcinoid|9091/1
C0334526|T191|SY|32071008|SNOMEDCT_US|Struma ovarii and carcinoid|9091/1
C0334526|T191|PT|32071008|SNOMEDCT_US|Strumal carcinoid|9091/1
C0020217|T191|PT|0026600|CCPSS|HYDATIDIFORM MOLE|9100/0
C0020217|T191|SY|0000006330|CHV|hydatid mole|9100/0
C0020217|T191|SY|0000006330|CHV|hydatidiform mole|9100/0
C0020217|T191|SY|0000006330|CHV|hydatidiform moles|9100/0
C0020217|T191|SY|0000006330|CHV|molar pregnancies|9100/0
C0020217|T191|PT|0000006330|CHV|molar pregnancy|9100/0
C0020217|T191|SY|0000006330|CHV|molars pregnancy|9100/0
C0020217|T191|SY|0000006330|CHV|mole hydatidiform|9100/0
C0020217|T191|SY|0000006330|CHV|mole pregnancy|9100/0
C0020217|T191|SY|0000006330|CHV|moles pregnancy|9100/0
C0020217|T191|SY|0000006330|CHV|pregnancy mole|9100/0
C0020217|T191|PT|NOCODE|COSTAR|Hydatidiform Mole|9100/0
C0020217|T191|PT|U000419|COSTAR|MOLAR PREGNANCY|9100/0
C0020217|T191|PT|2403-0989|CSP|hydatidiform mole|9100/0
C0020217|T191|ET|2403-0989|CSP|molar pregnancy|9100/0
C0020217|T191|ET|2403-0989|CSP|vesicular mole|9100/0
C0020217|T191|GT|NEOPL UTER|CST|HYDATIDIFORM MOLE|9100/0
C0020217|T191|FI|U002002|DXP|HYDATIDIFORM MOLE|9100/0
C0020217|T191|SY|NOCODE|DXP|MOLAR PREGNANCY|9100/0
C0020217|T191|SY|NOCODE|DXP|MOLE, HYDATID|9100/0
C0020217|T191|DI|U001195|DXP|MOLE, HYDATIDIFORM|9100/0
C0020217|T191|SY|NOCODE|DXP|PREGNANCY, MOLAR|9100/0
C0020217|T191|PT|HP:0032192|HPO|Hydatidiform mole|9100/0
C0020217|T191|PT|O01.0|ICD10|Classical hydatidiform mole|9100/0
C0020217|T191|HT|O01|ICD10|Hydatidiform mole|9100/0
C0020217|T191|PT|O01.9|ICD10|Hydatidiform mole, unspecified|9100/0
C0020217|T191|AB|O01.0|ICD10CM|Classical hydatidiform mole|9100/0
C0020217|T191|PT|O01.0|ICD10CM|Classical hydatidiform mole|9100/0
C0020217|T191|AB|O01|ICD10CM|Hydatidiform mole|9100/0
C0020217|T191|HT|O01|ICD10CM|Hydatidiform mole|9100/0
C0020217|T191|AB|O01.9|ICD10CM|Hydatidiform mole, unspecified|9100/0
C0020217|T191|PT|O01.9|ICD10CM|Hydatidiform mole, unspecified|9100/0
C0020217|T191|AB|630|ICD9CM|Hydatidiform mole|9100/0
C0020217|T191|PT|630|ICD9CM|Hydatidiform mole|9100/0
C0020217|T191|PT|MTHU041469|ICPC2ICD10ENG|classical; hydatidiform mole|9100/0
C0020217|T191|PT|MTHU035841|ICPC2ICD10ENG|hydatidiform mole|9100/0
C0020217|T191|PT|MTHU035844|ICPC2ICD10ENG|hydatidiform mole; classical|9100/0
C0020217|T191|PT|MTHU035849|ICPC2ICD10ENG|hydatidiform; mole|9100/0
C0020217|T191|PT|MTHU050164|ICPC2ICD10ENG|molar pregnancy|9100/0
C0020217|T191|PT|MTHU050183|ICPC2ICD10ENG|molar pregnancy; pregnancy|9100/0
C0020217|T191|PT|MTHU050142|ICPC2ICD10ENG|mole; hydatidiform|9100/0
C0020217|T191|PT|MTHU050145|ICPC2ICD10ENG|mole; hydatidiform, classical|9100/0
C0020217|T191|PT|MTHU050159|ICPC2ICD10ENG|mole; pregnancy, hydatidiform|9100/0
C0020217|T191|PT|MTHU050155|ICPC2ICD10ENG|mole; vesicular|9100/0
C0020217|T191|PT|MTHU083775|ICPC2ICD10ENG|pregnancy; hydatidiform mole|9100/0
C0020217|T191|PT|MTHU083873|ICPC2ICD10ENG|pregnancy; mole|9100/0
C0020217|T191|PT|MTHU083875|ICPC2ICD10ENG|pregnancy; mole, hydatidiform|9100/0
C0020217|T191|PT|MTHU080678|ICPC2ICD10ENG|vesicular; mole|9100/0
C0020217|T191|PT|W73002|ICPC2P|Hydatidiform mole|9100/0
C0020217|T191|PTN|W73002|ICPC2P|hydatidiform mole|9100/0
C0020217|T191|PT|U005660|LCH|Pregnancy, Molar|9100/0
C0020217|T191|PT|sh85106289|LCH_NW|Molar pregnancy|9100/0
C0020217|T191|LA|LA14685-4|LNC|Molar pregnancy|9100/0
C0549315|T191|LLT|10004272|MDR|Benign hydatidiform mole|9100/0
C0549315|T191|PT|10004272|MDR|Benign hydatidiform mole|9100/0
C0020217|T191|LLT|10020481|MDR|Hydatidiform mole|9100/0
C0549315|T191|LLT|10020482|MDR|Hydatidiform mole benign|9100/0
C0020217|T191|LLT|10020484|MDR|Hydatidiform mole NOS|9100/0
C0020217|T191|LLT|10065063|MDR|Molar pregnancy|9100/0
C0020217|T191|PT|30598|MEDCIN|hydatidiform mole|9100/0
C0020217|T191|SY|30598|MEDCIN|molar pregnancy|9100/0
C0020217|T191|ET|5534|MEDLINEPLUS|Molar Pregnancy|9100/0
C0020217|T191|ET|D006828|MSH|Hydatid Mole|9100/0
C0020217|T191|PM|D006828|MSH|Hydatid Moles|9100/0
C0020217|T191|MH|D006828|MSH|Hydatidiform Mole|9100/0
C0020217|T191|PM|D006828|MSH|Hydatidiform Moles|9100/0
C0020217|T191|DEV|D006828|MSH|MOLAR PREGN|9100/0
C0020217|T191|PM|D006828|MSH|Molar Pregnancies|9100/0
C0020217|T191|ET|D006828|MSH|Molar Pregnancy|9100/0
C0020217|T191|PM|D006828|MSH|Mole, Hydatid|9100/0
C0020217|T191|PM|D006828|MSH|Mole, Hydatidiform|9100/0
C0020217|T191|PM|D006828|MSH|Moles, Hydatid|9100/0
C0020217|T191|PM|D006828|MSH|Moles, Hydatidiform|9100/0
C0020217|T191|DEV|D006828|MSH|PREGN MOLAR|9100/0
C0020217|T191|PM|D006828|MSH|Pregnancies, Molar|9100/0
C0020217|T191|ET|D006828|MSH|Pregnancy, Molar|9100/0
C0020217|T191|PN|NOCODE|MTH|Hydatidiform Mole|9100/0
C0020217|T191|ET|630|MTHICD9|Vesicular mole|9100/0
C0020217|T191|SY|C3110|NCI|Hydatid Mole|9100/0
C0020217|T191|PT|C3110|NCI|Hydatidiform Mole|9100/0
C0020217|T191|SY|C3110|NCI|Molar Pregnancy|9100/0
C0020217|T191|DN|C3110|NCI_CTRP|Hydatidiform Mole|9100/0
C0020217|T191|PT|CDR0000446933|NCI_NCI-GLOSS|hydatidiform mole|9100/0
C0020217|T191|PT|CDR0000046747|NCI_NCI-GLOSS|molar pregnancy|9100/0
C0020217|T191|PT|C3110|NCI_NICHD|Hydatidiform Mole|9100/0
C0020217|T191|SY|CDR0000040675|PDQ|chorionic tumor|9100/0
C0020217|T191|SY|CDR0000040675|PDQ|gestational trophoblastic tumor, hydatidiform mole|9100/0
C0020217|T191|SY|CDR0000040675|PDQ|GTT, hydatidiform mole|9100/0
C0020217|T191|SY|CDR0000040675|PDQ|hydatid mole|9100/0
C0020217|T191|PSC|CDR0000040675|PDQ|hydatidiform mole|9100/0
C0020217|T191|SY|CDR0000040675|PDQ|hydatidiform mole GTT|9100/0
C0020217|T191|SY|CDR0000040675|PDQ|molar pregnancy|9100/0
C0020217|T191|SY|L000.|RCD|Classical hydatidiform mole|9100/0
C0020217|T191|SY|L000.|RCD|Hydatid mole|9100/0
C0020217|T191|PT|L000.|RCD|Hydatidiform mole|9100/0
C0020217|T191|OP|BBR0.|RCDSY|Hydatidiform mole NOS|9100/0
C0020217|T191|OAS|235323008|SNOMEDCT_US|Classical hydatidiform mole|9100/0
C0020217|T191|OAS|235323008|SNOMEDCT_US|Hydatid mole|9100/0
C0020217|T191|SY|417044008|SNOMEDCT_US|Hydatid mole|9100/0
C0020217|T191|SY|48430004|SNOMEDCT_US|Hydatid mole|9100/0
C0020217|T191|SY|417044008|SNOMEDCT_US|Hydatidiform mole|9100/0
C0020217|T191|OAP|156085008|SNOMEDCT_US|Hydatidiform mole|9100/0
C0020217|T191|PT|48430004|SNOMEDCT_US|Hydatidiform mole|9100/0
C0020217|T191|OAP|198611007|SNOMEDCT_US|Hydatidiform mole|9100/0
C0020217|T191|OAP|235323008|SNOMEDCT_US|Hydatidiform mole|9100/0
C0020217|T191|OAS|198610008|SNOMEDCT_US|Hydatidiform mole|9100/0
C0020217|T191|OF|156085008|SNOMEDCT_US|Hydatidiform mole|9100/0
C0549315|T191|PT|417044008|SNOMEDCT_US|Hydatidiform mole, benign|9100/0
C0549315|T191|PT|417271000|SNOMEDCT_US|Hydatidiform mole, benign|9100/0
C0020217|T191|SY|48430004|SNOMEDCT_US|Hydatidiform mole, no ICD-O subtype|9100/0
C0020217|T191|SY|48430004|SNOMEDCT_US|Hydatidiform mole, no International Classification of Diseases for Oncology subtype|9100/0
C0020217|T191|IS|48430004|SNOMEDCT_US|Hydatidiform mole, NOS|9100/0
C0020217|T191|PT|44782008|SNOMEDCT_US|Molar pregnancy|9100/0
C0020217|T191|IS|41491009|SNOMEDCT_US|Molar pregnancy with hydatid mole|9100/0
C0020217|T191|OAS|367455000|SNOMEDCT_US|Molar pregnancy with hydatid mole|9100/0
C0020217|T191|SY|417044008|SNOMEDCT_US|Molar pregnancy with hydatid mole|9100/0
C0020217|T191|OAP|41491009|SNOMEDCT_US|Molar pregnancy with hydatidiform mole|9100/0
C0020217|T191|OAP|367455000|SNOMEDCT_US|Molar pregnancy with hydatidiform mole|9100/0
C0020217|T191|IS|41491009|SNOMEDCT_US|Molar pregnancy with vesicular mole|9100/0
C0020217|T191|OAP|236118006|SNOMEDCT_US|Molar pregnancy with vesicular mole|9100/0
C0020217|T191|OAS|367455000|SNOMEDCT_US|Molar pregnancy with vesicular mole|9100/0
C0020217|T191|SY|417044008|SNOMEDCT_US|Molar pregnancy with vesicular mole|9100/0
C0020217|T191|IS|44782008|SNOMEDCT_US|Molar pregnancy, NOS|9100/0
C0020217|T191|OAP|123300001|SNOMEDCT_US|Mole|9100/0
C0020217|T191|IS|123300001|SNOMEDCT_US|Mole -RETIRED-|9100/0
C0020217|T191|OF|123300001|SNOMEDCT_US|Mole -RETIRED-|9100/0
C0020217|T191|SY|44782008|SNOMEDCT_US|Mole of pregnancy|9100/0
C0020217|T191|IS|44782008|SNOMEDCT_US|Mole of pregnancy, NOS|9100/0
C0020217|T191|IS|123300001|SNOMEDCT_US|Mole, NOS|9100/0
C0020217|T191|OAS|198610008|SNOMEDCT_US|Vesicular mole|9100/0
C0020217|T191|PT|0831|WHO|HYDATIDIFORM MOLE|9100/0
C0549315|T191|IT|0831|WHO|HYDATIDIFORM MOLE BENIGN|9100/0
C0008493|T191|SY|0000002908|CHV|chorioadenoma|9100/1
C0008493|T191|SY|0000002908|CHV|chorioadenoma destruens|9100/1
C0008493|T191|SY|0000002908|CHV|invasive hydatidiform mole|9100/1
C0008493|T191|PT|0000002908|CHV|invasive mole|9100/1
C0008493|T191|SY|0000002908|CHV|malignant mole|9100/1
C0008493|T191|SY|0000002908|CHV|malignant moles|9100/1
C0008493|T191|DI|U000347|DXP|CHORIOADENOMA DESTRUENS|9100/1
C0008493|T191|SY|NOCODE|DXP|MOLE, DESTRUCTIVE|9100/1
C0008493|T191|SY|NOCODE|DXP|MOLE, INVASIVE|9100/1
C0008493|T191|SY|NOCODE|DXP|MOLE, MALIGNANT|9100/1
C0008493|T191|ET|D39.2|ICD10CM|Chorioadenoma destruens|9100/1
C0008493|T191|ET|D39.2|ICD10CM|Invasive hydatidiform mole|9100/1
C0008493|T191|ET|D39.2|ICD10CM|Malignant hydatidiform mole|9100/1
C0008493|T191|PT|MTHU022699|ICPC2ICD10ENG|destructive; mole|9100/1
C0008493|T191|PT|MTHU035843|ICPC2ICD10ENG|hydatidiform mole; invasive|9100/1
C0008493|T191|PT|MTHU035845|ICPC2ICD10ENG|hydatidiform mole; malignant|9100/1
C0008493|T191|PT|MTHU040176|ICPC2ICD10ENG|invasive; hydatidiform mole|9100/1
C0008493|T191|PT|MTHU040177|ICPC2ICD10ENG|invasive; mole|9100/1
C0008493|T191|PT|MTHU047293|ICPC2ICD10ENG|malignant; hydatidiform mole|9100/1
C0008493|T191|PT|MTHU047301|ICPC2ICD10ENG|malignant; mole, hydatidiform|9100/1
C0008493|T191|PT|MTHU050140|ICPC2ICD10ENG|mole; destructive|9100/1
C0008493|T191|PT|MTHU050144|ICPC2ICD10ENG|mole; hydatidiform, invasive|9100/1
C0008493|T191|PT|MTHU050146|ICPC2ICD10ENG|mole; hydatidiform, malignant|9100/1
C0008493|T191|PT|MTHU050151|ICPC2ICD10ENG|mole; invasive|9100/1
C0008493|T191|PT|MTHU050152|ICPC2ICD10ENG|mole; malignant, hydatidiform mole|9100/1
C0008493|T191|PTN|S77010|ICPC2P|malignant mole|9100/1
C0008493|T191|PT|S77010|ICPC2P|Mole;malignant|9100/1
C0008493|T191|LLT|10020483|MDR|Hydatidiform mole malignant|9100/1
C0008493|T191|PT|10025598|MDR|Malignant hydatidiform mole|9100/1
C0008493|T191|LLT|10025598|MDR|Malignant hydatidiform mole|9100/1
C0008493|T191|PT|34981|MEDCIN|invasive hydatidiform mole|9100/1
C0008493|T191|ET|D002820|MSH|Chorioadenoma|9100/1
C0008493|T191|PM|D002820|MSH|Chorioadenomas|9100/1
C0008493|T191|MH|D002820|MSH|Hydatidiform Mole, Invasive|9100/1
C0008493|T191|PM|D002820|MSH|Hydatidiform Moles, Invasive|9100/1
C0008493|T191|PM|D002820|MSH|Invasive Hydatidiform Mole|9100/1
C0008493|T191|PM|D002820|MSH|Invasive Hydatidiform Moles|9100/1
C0008493|T191|ET|D002820|MSH|Invasive Mole|9100/1
C0008493|T191|PM|D002820|MSH|Invasive Moles|9100/1
C0008493|T191|PM|D002820|MSH|Mole, Invasive|9100/1
C0008493|T191|PM|D002820|MSH|Mole, Invasive Hydatidiform|9100/1
C0008493|T191|PM|D002820|MSH|Moles, Invasive|9100/1
C0008493|T191|PM|D002820|MSH|Moles, Invasive Hydatidiform|9100/1
C0008493|T191|ET|236.1|MTHICD9|Chorioadenoma|9100/1
C0008493|T191|ET|236.1|MTHICD9|Chorioadenoma destruens|9100/1
C0008493|T191|ET|236.1|MTHICD9|Invasive mole|9100/1
C0008493|T191|ET|236.1|MTHICD9|Malignant hydatid mole|9100/1
C0008493|T191|ET|236.1|MTHICD9|Malignant hydatidiform mole|9100/1
C0008493|T191|SY|C6985|NCI|Chorioadenoma|9100/1
C0008493|T191|SY|C6985|NCI|Chorioadenoma Destruens|9100/1
C0008493|T191|SY|C6985|NCI|Invasive Gestational Trophoblastic Neoplasm|9100/1
C0008493|T191|PT|C6985|NCI|Invasive Hydatidiform Mole|9100/1
C0008493|T191|SY|C6985|NCI|Invasive Mole|9100/1
C0008493|T191|DN|C6985|NCI_CTRP|Invasive Hydatidiform Mole|9100/1
C0008493|T191|PT|CDR0000458034|NCI_NCI-GLOSS|chorioadenoma destruens|9100/1
C0008493|T191|PT|CDR0000446955|NCI_NCI-GLOSS|invasive hydatidiform mole|9100/1
C0008493|T191|PT|C6985|NCI_NICHD|Invasive Hydatidiform Mole|9100/1
C0008493|T191|SY|CDR0000039967|PDQ|chorioadenoma|9100/1
C0008493|T191|PT|CDR0000039967|PDQ|chorioadenoma destruens|9100/1
C0008493|T191|SY|CDR0000039967|PDQ|gestational trophoblastic tumor, invasive mole|9100/1
C0008493|T191|SY|CDR0000039967|PDQ|GTT, invasive mole|9100/1
C0008493|T191|SY|CDR0000039967|PDQ|Invasive Gestational Trophoblastic Neoplasm|9100/1
C0008493|T191|SY|CDR0000039967|PDQ|Invasive Hydatidiform Mole|9100/1
C0008493|T191|SY|CDR0000039967|PDQ|invasive mole|9100/1
C0008493|T191|SY|XE2vj|RCD|Chorioadenoma|9100/1
C0008493|T191|SY|XE2vj|RCD|Chorioadenoma destruens|9100/1
C0008493|T191|SY|XE2vj|RCD|IM - Invasive mole|9100/1
C0008493|T191|SY|XE2vj|RCD|Invasive hydatidiform mole|9100/1
C0008493|T191|SY|XE2vj|RCD|Invasive mole|9100/1
C0008493|T191|SY|XE2vj|RCD|Invasive mole - placenta|9100/1
C0008493|T191|PT|XE2vj|RCD|Malignant hydatidiform mole|9100/1
C0008493|T191|SY|BBR1.|RCDSY|Chorioadenoma|9100/1
C0008493|T191|SY|BBR1.|RCDSY|Chorioadenoma destruens|9100/1
C0008493|T191|PT|BBR1.|RCDSY|Invasive hydatidiform mole|9100/1
C0008493|T191|SY|416669000|SNOMEDCT_US|Chorioadenoma|9100/1
C0008493|T191|SY|18799007|SNOMEDCT_US|Chorioadenoma|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Chorioadenoma|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Chorioadenoma destruens|9100/1
C0008493|T191|SY|416669000|SNOMEDCT_US|Chorioadenoma destruens|9100/1
C0008493|T191|SY|18799007|SNOMEDCT_US|Chorioadenoma destruens|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|IM - Invasive mole|9100/1
C0008493|T191|SY|416669000|SNOMEDCT_US|IM - Invasive mole|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Invasive hydatidiform mole|9100/1
C0008493|T191|PT|416669000|SNOMEDCT_US|Invasive hydatidiform mole|9100/1
C0008493|T191|PT|18799007|SNOMEDCT_US|Invasive hydatidiform mole|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Invasive mole|9100/1
C0008493|T191|SY|416669000|SNOMEDCT_US|Invasive mole|9100/1
C0008493|T191|SY|18799007|SNOMEDCT_US|Invasive mole|9100/1
C0008493|T191|OAS|189444004|SNOMEDCT_US|Invasive mole - placenta|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Invasive mole - placenta|9100/1
C0008493|T191|SY|416669000|SNOMEDCT_US|Invasive mole - placenta|9100/1
C0008493|T191|IS|18799007|SNOMEDCT_US|Invasive mole, NOS|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Malignant hydatidiform mole|9100/1
C0008493|T191|OF|154643005|SNOMEDCT_US|Malignant hydatidiform mole|9100/1
C0008493|T191|SY|18799007|SNOMEDCT_US|Malignant hydatidiform mole|9100/1
C0008493|T191|OAP|154643005|SNOMEDCT_US|Malignant hydatidiform mole|9100/1
C0008493|T191|OAS|189444004|SNOMEDCT_US|Malignant hydatidiform mole|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Molar pregnancy with chorioadenoma|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Molar pregnancy with chorioadenoma destruens|9100/1
C0008493|T191|OAP|74153005|SNOMEDCT_US|Molar pregnancy with invasive hydatidiform mole|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Molar pregnancy with invasive mole|9100/1
C0008493|T191|OAS|74153005|SNOMEDCT_US|Molar pregnancy with malignant hydatidiform mole|9100/1
C0008497|T191|PT|1006588|CCPSS|CHORIOCARCINOMA|9100/3
C0008497|T191|PT|0000041850|CHV|chorioblastoma|9100/3
C0008497|T191|PT|0000002910|CHV|choriocarcinoma|9100/3
C0008497|T191|SY|0000002910|CHV|chorioepithelioma|9100/3
C0008497|T191|SY|0000002910|CHV|chorionepithelioma|9100/3
C0008497|T191|PT|U000136|COSTAR|CHORIOCARCINOMA|9100/3
C0008497|T191|ET|2000-4323|CSP|chordocarcinoma|9100/3
C0008497|T191|ET|2000-4323|CSP|chordoepithelioma|9100/3
C0008497|T191|ET|2403-0675|CSP|chorioblastoma|9100/3
C0008497|T191|PT|2403-0675|CSP|choriocarcinoma|9100/3
C0008497|T191|ET|2403-0675|CSP|chorioepithelioma|9100/3
C0008497|T191|PT|HP:0100768|HPO|Choriocarcinoma|9100/3
C0008497|T191|ET|C58|ICD10CM|choriocarcinoma NOS|9100/3
C0008497|T191|ET|C58|ICD10CM|chorionepithelioma NOS|9100/3
C0008497|T191|PT|MTHU016400|ICPC2ICD10ENG|choriocarcinoma|9100/3
C0008497|T191|PTN|W72002|ICPC2P|chorioepithelioma|9100/3
C0008497|T191|PT|W72002|ICPC2P|Chorioepithelioma|9100/3
C0008497|T191|PT|U000999|LCH|Choriocarcinoma|9100/3
C0008497|T191|PT|sh85024747|LCH_NW|Choriocarcinoma|9100/3
C0008497|T191|LLT|10008757|MDR|Choriocarcinoma|9100/3
C0008497|T191|PT|10008757|MDR|Choriocarcinoma|9100/3
C0008497|T191|LLT|10008759|MDR|Choriocarcinoma NOS|9100/3
C0008497|T191|PT|271551|MEDCIN|choriocarcinoma|9100/3
C0008497|T191|MH|D002822|MSH|Choriocarcinoma|9100/3
C0008497|T191|PM|D002822|MSH|Choriocarcinomas|9100/3
C0008497|T191|PN|NOCODE|MTH|Choriocarcinoma|9100/3
C0008497|T191|ET|181|MTHICD9|Choriocarcinoma NOS|9100/3
C0008497|T191|ET|181|MTHICD9|Chorioepithelioma NOS|9100/3
C0008497|T191|SY|TCGA|NCI|Choriocarcinoma|9100/3
C0008497|T191|PT|C2948|NCI|Choriocarcinoma|9100/3
C0008497|T191|SY|C2948|NCI|Chorioepithelioma|9100/3
C0349557|T191|PT|C4646|NCI|Gestational Choriocarcinoma|9100/3
C0008497|T191|PT|C2948|NCI_CDISC|CHORIOCARCINOMA, MALIGNANT|9100/3
C0008497|T191|SY|C2948|NCI_CDISC|Chorioepithelioma|9100/3
C0008497|T191|PT|C2948|NCI_CPTAC|Choriocarcinoma|9100/3
C0008497|T191|DN|C2948|NCI_CTRP|Choriocarcinoma|9100/3
C0008497|T191|PT|C2948|NCI_CTRP|Choriocarcinoma|9100/3
C0008497|T191|PT|CDR0000554834|NCI_NCI-GLOSS|chorioblastoma|9100/3
C0008497|T191|PT|CDR0000046753|NCI_NCI-GLOSS|choriocarcinoma|9100/3
C0008497|T191|PT|CDR0000554835|NCI_NCI-GLOSS|chorioepithelioma|9100/3
C0008497|T191|PT|CDR0000554836|NCI_NCI-GLOSS|chorionic carcinoma|9100/3
C0008497|T191|OP|B420.|RCD|Choriocarcinoma|9100/3
C0008497|T191|IS|B420.|RCD|Chorioepithelioma|9100/3
C0008497|T191|IS|B420.|RCD|Chorionepithelioma|9100/3
C0349557|T191|PT|X78Y1|RCD|Gestational choriocarcinoma|9100/3
C0008497|T191|PT|BBR2.|RCDSY|Choriocarcinoma|9100/3
C0008497|T191|SY|BBR2.|RCDSY|Chorioepithelioma|9100/3
C1275855|T191|SY|399380001|SNOMEDCT_US|Biphasic choriocarcinoma|9100/3
C0008497|T191|OAS|189444004|SNOMEDCT_US|Choriocarcinoma|9100/3
C0008497|T191|PT|188188009|SNOMEDCT_US|Choriocarcinoma|9100/3
C0008497|T191|PT|44769000|SNOMEDCT_US|Choriocarcinoma|9100/3
C1275855|T191|PT|399380001|SNOMEDCT_US|Choriocarcinoma, biphasic|9100/3
C1275871|T191|PT|399669007|SNOMEDCT_US|Choriocarcinoma, monophasic|9100/3
C0008497|T191|SY|44769000|SNOMEDCT_US|Choriocarcinoma, no ICD-O subtype|9100/3
C0008497|T191|SY|44769000|SNOMEDCT_US|Choriocarcinoma, no International Classification of Diseases for Oncology subtype|9100/3
C0008497|T191|IS|44769000|SNOMEDCT_US|Choriocarcinoma, NOS|9100/3
C0008497|T191|SY|188188009|SNOMEDCT_US|Chorioepithelioma|9100/3
C0008497|T191|SY|44769000|SNOMEDCT_US|Chorioepithelioma|9100/3
C0008497|T191|SY|44769000|SNOMEDCT_US|Chorionepithelioma|9100/3
C0008497|T191|SY|188188009|SNOMEDCT_US|Chorionepithelioma|9100/3
C0349557|T191|PT|417057000|SNOMEDCT_US|Gestational choriocarcinoma|9100/3
C0349557|T191|OAS|1884006|SNOMEDCT_US|Gestational choriocarcinoma|9100/3
C0349557|T191|PT|417570003|SNOMEDCT_US|Gestational choriocarcinoma|9100/3
C0349557|T191|SY|417570003|SNOMEDCT_US|Gestational chorioepithelioma|9100/3
C0349557|T191|SY|417570003|SNOMEDCT_US|Gestational chorionepithelioma|9100/3
C0349557|T191|OAP|1884006|SNOMEDCT_US|Molar pregnancy with choriocarcinoma|9100/3
C0349557|T191|OAS|1884006|SNOMEDCT_US|Molar pregnancy with chorioepithelioma|9100/3
C0349557|T191|OAS|1884006|SNOMEDCT_US|Molar pregnancy with chorionepithelioma|9100/3
C1275871|T191|SY|399669007|SNOMEDCT_US|Monophasic choriocarcinoma|9100/3
C0008497|T191|SY|44769000|SNOMEDCT_US|Syncytioma|9100/3
C1298201|T191|PT|10071532|MDR|Metastatic choriocarcinoma|9100/6
C1298201|T191|LLT|10071532|MDR|Metastatic choriocarcinoma|9100/6
C1298201|T191|PT|370079006|SNOMEDCT_US|Choriocarcinoma, metastatic|9100/6
C0334527|T191|PT|271552|MEDCIN|choriocarcinoma combined with other germ cell elements|9101/3
C0334527|T191|PT|C66777|NCI|Choriocarcinoma Combined with Other Germ Cell Elements|9101/3
C0334527|T191|AB|Xa9AQ|RCD|Chorioca + germ cell elements|9101/3
C0334527|T191|AB|Xa9AQ|RCD|Chorioca with embryonal ca|9101/3
C0334527|T191|SY|Xa9AQ|RCD|Choriocarcinoma combined with embryonal carcinoma|9101/3
C0334527|T191|PT|Xa9AQ|RCD|Choriocarcinoma combined with germ cell elements|9101/3
C0600067|T191|OP|BBR3.|RCD|Choriocarcinoma combined with teratoma|9101/3
C0600067|T191|OA|BBR3.|RCD|Choriocarcinoma with teratoma|9101/3
C0334527|T191|SY|8734000|SNOMEDCT_US|Choriocarcinoma combined with embryonal carcinoma|9101/3
C0334527|T191|SY|8734000|SNOMEDCT_US|Choriocarcinoma combined with germ cell elements|9101/3
C0334527|T191|PT|8734000|SNOMEDCT_US|Choriocarcinoma combined with other germ cell elements|9101/3
C0600067|T191|PT|189857001|SNOMEDCT_US|Choriocarcinoma combined with teratoma|9101/3
C0600067|T191|SY|8734000|SNOMEDCT_US|Choriocarcinoma combined with teratoma|9101/3
C0334528|T191|PT|MTHU047311|ICPC2ICD10ENG|malignant; teratoma, trophoblastic, unspecified site|9102/3
C0334528|T191|PT|MTHU073784|ICPC2ICD10ENG|teratoma; malignant, trophoblastic, unspecified site|9102/3
C0334528|T191|SY|271550|MEDCIN|malignant trophoblastic teratoma|9102/3
C0334528|T191|PT|271550|MEDCIN|trophoblastic malignant teratoma|9102/3
C0334528|T191|PN|NOCODE|MTH|Malignant Trophoblastic Teratoma|9102/3
C0334528|T191|OP|C66778|NCI|Malignant Trophoblastic Teratoma|9102/3
C0334528|T191|PT|C66778|NCI|Malignant Trophoblastic Teratoma|9102/3
C0334528|T191|AB|BBR4.|RCD|Trophoblastic malign teratoma|9102/3
C0334528|T191|PT|BBR4.|RCD|Trophoblastic malignant teratoma|9102/3
C0334528|T191|PT|65646006|SNOMEDCT_US|Malignant teratoma, trophoblastic|9102/3
C0334528|T191|SY|65646006|SNOMEDCT_US|Trophoblastic malignant teratoma|9102/3
C0334529|T191|PT|O01.1|ICD10|Incomplete and partial hydatidiform mole|9103/0
C0334529|T191|AB|O01.1|ICD10CM|Incomplete and partial hydatidiform mole|9103/0
C0334529|T191|PT|O01.1|ICD10CM|Incomplete and partial hydatidiform mole|9103/0
C0334529|T191|PT|MTHU035846|ICPC2ICD10ENG|hydatidiform mole; partial|9103/0
C0334529|T191|PT|MTHU050147|ICPC2ICD10ENG|mole; hydatidiform, incomplete|9103/0
C0334529|T191|PT|MTHU050148|ICPC2ICD10ENG|mole; hydatidiform, partial|9103/0
C0334529|T191|PT|MTHU058008|ICPC2ICD10ENG|partial; hydatidiform mole|9103/0
C0334529|T191|PEP|D006828|MSH|Hydatidiform Mole, Partial|9103/0
C0334529|T191|PM|D006828|MSH|Hydatidiform Moles, Partial|9103/0
C0334529|T191|PM|D006828|MSH|Mole, Partial Hydatidiform|9103/0
C0334529|T191|PM|D006828|MSH|Moles, Partial Hydatidiform|9103/0
C0334529|T191|PM|D006828|MSH|Partial Hydatidiform Mole|9103/0
C0334529|T191|PM|D006828|MSH|Partial Hydatidiform Moles|9103/0
C0334529|T191|SY|C4293|NCI|Incomplete Hydatid Mole|9103/0
C0334529|T191|SY|C4293|NCI|Incomplete Hydatidiform Mole|9103/0
C0334529|T191|SY|C4293|NCI|Incomplete Molar Pregnancy|9103/0
C0334529|T191|SY|C4293|NCI|Partial Hydatid Mole|9103/0
C0334529|T191|PT|C4293|NCI|Partial Hydatidiform Mole|9103/0
C0334529|T191|SY|C4293|NCI|Partial Molar Pregnancy|9103/0
C0334529|T191|SY|C4293|NCI|Partial Mole|9103/0
C0334529|T191|SY|C4293|NCI_NICHD|Incomplete Hydatidiform Mole|9103/0
C0334529|T191|PT|C4293|NCI_NICHD|Partial Hydatidiform Mole|9103/0
C0334529|T191|PT|X40B5|RCD|Incomplete hydatidiform mole|9103/0
C0334529|T191|SY|X40B5|RCD|Partial hydatidiform mole|9103/0
C0334529|T191|AB|X40B5|RCD|PHM - Partial hydatid mole|9103/0
C0334529|T191|SY|X40B5|RCD|PHM - Partial hydatidiform mole|9103/0
C0334529|T191|OP|BBR5.|RCDSY|Partial hydatidiform mole|9103/0
C0334529|T191|OAP|198612000|SNOMEDCT_US|Incomplete hydatidiform mole|9103/0
C0334529|T191|OF|198612000|SNOMEDCT_US|Incomplete hydatidiform mole|9103/0
C0334529|T191|SY|237250000|SNOMEDCT_US|Incomplete hydatidiform mole|9103/0
C0334529|T191|PT|237250000|SNOMEDCT_US|Partial hydatidiform mole|9103/0
C0334529|T191|PT|51793002|SNOMEDCT_US|Partial hydatidiform mole|9103/0
C0334529|T191|SY|51793002|SNOMEDCT_US|Partial mole|9103/0
C0334529|T191|SY|237250000|SNOMEDCT_US|PHM - Partial hydatidiform mole|9103/0
C0206666|T191|PT|MTHU077139|ICPC2ICD10ENG|tumor; placental site trophoblastic|9104/1
C0206666|T191|PM|D018245|MSH|Placental Site Trophoblastic Tumor|9104/1
C0206666|T191|PM|D018245|MSH|Placental Trophoblastic Tumor|9104/1
C0206666|T191|PM|D018245|MSH|Placental Trophoblastic Tumors|9104/1
C0206666|T191|ET|D018245|MSH|Placental-Site Trophoblastic Tumor|9104/1
C0206666|T191|PM|D018245|MSH|Placental-Site Trophoblastic Tumors|9104/1
C0206666|T191|ET|D018245|MSH|Trophoblastic Tumor, Placental|9104/1
C0206666|T191|MH|D018245|MSH|Trophoblastic Tumor, Placental Site|9104/1
C0206666|T191|PM|D018245|MSH|Trophoblastic Tumor, Placental-Site|9104/1
C0206666|T191|PM|D018245|MSH|Trophoblastic Tumors, Placental|9104/1
C0206666|T191|PM|D018245|MSH|Trophoblastic Tumors, Placental-Site|9104/1
C0206666|T191|PM|D018245|MSH|Tumor, Placental Trophoblastic|9104/1
C0206666|T191|PM|D018245|MSH|Tumor, Placental-Site Trophoblastic|9104/1
C0206666|T191|PM|D018245|MSH|Tumors, Placental Trophoblastic|9104/1
C0206666|T191|PM|D018245|MSH|Tumors, Placental-Site Trophoblastic|9104/1
C0206666|T191|SY|C3757|NCI|Placental Site Gestational Trophoblastic Tumor|9104/1
C0206666|T191|SY|C3757|NCI|Placental-Site Gestational Trophoblastic Neoplasm|9104/1
C0206666|T191|PT|C3757|NCI|Placental-Site Gestational Trophoblastic Tumor|9104/1
C0206666|T191|SY|C3757|NCI|Placental-Site GTT|9104/1
C0206666|T191|SY|CDR0000041357|PDQ|gestational trophoblastic tumor, placental site|9104/1
C0206666|T191|SY|CDR0000041357|PDQ|gestational trophoblastic tumor, placental-site|9104/1
C0206666|T191|SY|CDR0000041357|PDQ|GTT, placental site|9104/1
C0206666|T191|SY|CDR0000041357|PDQ|GTT, placental-site|9104/1
C0206666|T191|SY|CDR0000041357|PDQ|placental site gestational trophoblastic tumor|9104/1
C0206666|T191|SY|CDR0000041357|PDQ|placental site GTT|9104/1
C0206666|T191|PSC|CDR0000041357|PDQ|placental-site gestational trophoblastic tumor|9104/1
C0206666|T191|SY|CDR0000041357|PDQ|placental-site GTT|9104/1
C0206666|T191|AB|X40B9|RCD|Placental site trophob tumour|9104/1
C0206666|T191|PT|X40B9|RCD|Placental site trophoblastic tumour|9104/1
C0206666|T191|AB|X40B9|RCDAE|Placental site trophob tumor|9104/1
C0206666|T191|PT|X40B9|RCDAE|Placental site trophoblastic tumor|9104/1
C0206666|T191|OP|BBR6.|RCDSA|Placental site trophoblastic tumor|9104/1
C0206666|T191|OP|BBR6.|RCDSY|Placental site trophoblastic tumour|9104/1
C0206666|T191|OA|BBR6.|RCDSY|Placental trophoblast tumur|9104/1
C0206666|T191|PT|75320001|SNOMEDCT_US|Placental site trophoblastic tumor|9104/1
C0206666|T191|PT|237252008|SNOMEDCT_US|Placental site trophoblastic tumor|9104/1
C0206666|T191|PTGB|75320001|SNOMEDCT_US|Placental site trophoblastic tumour|9104/1
C0206666|T191|PTGB|237252008|SNOMEDCT_US|Placental site trophoblastic tumour|9104/1
C1266159|T191|PT|271553|MEDCIN|malignant epithelioid trophoblastic tumor|9105/3
C1266159|T191|PT|C6900|NCI|Epithelioid Trophoblastic Tumor|9105/3
C1266159|T191|DN|C6900|NCI_CTRP|Epithelioid Trophoblastic Tumor|9105/3
C1266159|T191|PT|CDR0000709370|PDQ|epithelioid trophoblastic tumor|9105/3
C1266159|T191|PT|609515005|SNOMEDCT_US|Epithelioid trophoblastic tumor|9105/3
C1266159|T191|PTGB|609515005|SNOMEDCT_US|Epithelioid trophoblastic tumour|9105/3
C1266159|T191|PT|128767001|SNOMEDCT_US|Trophoblastic tumor, epithelioid|9105/3
C1266159|T191|PTGB|128767001|SNOMEDCT_US|Trophoblastic tumour, epithelioid|9105/3
C0334530|T191|PT|C4294|NCI|Benign Mesonephroma|9110/0
C0334530|T191|SY|C4294|NCI|Mesonephric Adenoma|9110/0
C1514905|T191|PT|C40018|NCI|Rete Ovarii Adenoma|9110/0
C0334530|T191|SY|C4294|NCI|Wolffian Duct Adenoma|9110/0
C1514905|T191|PT|C40018|NCI_CDISC|ADENOMA, RETE OVARII, BENIGN|9110/0
C0334530|T191|PT|BBS0.|RCD|Benign mesonephroma|9110/0
C0334530|T191|SY|BBS0.|RCD|Mesonephric adenoma|9110/0
C0334530|T191|SY|BBS0.|RCD|Wolffian duct adenoma|9110/0
C1514905|T191|PT|703654008|SNOMEDCT_US|Adenoma of rete ovarii|9110/0
C0334530|T191|SY|72889001|SNOMEDCT_US|Benign mesonephroma|9110/0
C0334530|T191|SY|72889001|SNOMEDCT_US|Mesonephric adenoma|9110/0
C0334530|T191|PT|72889001|SNOMEDCT_US|Mesonephroma, benign|9110/0
C0334530|T191|SY|72889001|SNOMEDCT_US|Wolffian duct adenoma|9110/0
C0334531|T191|PN|NOCODE|MTH|Mesonephric tumor|9110/1
C0334531|T191|PT|C4295|NCI|Mesonephric Neoplasm|9110/1
C0334531|T191|SY|C4295|NCI|Mesonephric Tumor|9110/1
C0334531|T191|SY|C4295|NCI|Mesonephroma|9110/1
C0334531|T191|SY|C4295|NCI|Wolffian Duct Neoplasm|9110/1
C0334531|T191|SY|C4295|NCI|Wolffian Duct Tumor|9110/1
C0334531|T191|PT|CDR0000335092|NCI_NCI-GLOSS|mesonephroma|9110/1
C0334531|T191|SY|BBS..|RCD|Mesonephric tumour|9110/1
C0334531|T191|SY|BBS..|RCDAE|Mesonephric tumor|9110/1
C0334531|T191|OP|BBS1.|RCDSA|Mesonephric tumor|9110/1
C0334531|T191|OP|BBS1.|RCDSY|Mesonephric tumour|9110/1
C0334531|T191|SY|127577004|SNOMEDCT_US|Mesonephric neoplasm|9110/1
C0334531|T191|OAP|13071008|SNOMEDCT_US|Mesonephric tumor|9110/1
C5230997|T191|SY|817967001|SNOMEDCT_US|Mesonephric tumor uncertain whether benign or malignant|9110/1
C0334531|T191|OAP|13071008|SNOMEDCT_US|Mesonephric tumour|9110/1
C5230997|T191|SYGB|817967001|SNOMEDCT_US|Mesonephric tumour uncertain whether benign or malignant|9110/1
C0334531|T191|OAS|13071008|SNOMEDCT_US|Wolffian duct tumor|9110/1
C5230997|T191|SY|817967001|SNOMEDCT_US|Wolffian duct tumor uncertain whether benign or malignant|9110/1
C0334531|T191|OAS|13071008|SNOMEDCT_US|Wolffian duct tumour|9110/1
C5230997|T191|SYGB|817967001|SNOMEDCT_US|Wolffian duct tumour uncertain whether benign or malignant|9110/1
C5230997|T191|PT|817967001|SNOMEDCT_US|Wolffian tumor uncertain whether benign or malignant|9110/1
C5230997|T191|PTGB|817967001|SNOMEDCT_US|Wolffian tumour uncertain whether benign or malignant|9110/1
C0025490|T191|SY|0000007990|CHV|mesonephric adenocarcinoma|9110/3
C0025490|T191|PT|0000007990|CHV|mesonephroma|9110/3
C0025490|T191|PT|MTHU048924|ICPC2ICD10ENG|mesonephroma|9110/3
C0025490|T191|PT|271554|MEDCIN|malignant mesonephroma|9110/3
C0025490|T191|MH|D008649|MSH|Mesonephroma|9110/3
C0025490|T191|PM|D008649|MSH|Mesonephromas|9110/3
C0025490|T191|PN|NOCODE|MTH|Mesonephroma|9110/3
C0025490|T191|SY|C4072|NCI|Malignant Mesonephroma|9110/3
C0025490|T191|PT|C4072|NCI|Mesonephric Adenocarcinoma|9110/3
C3840223|T191|PT|C40017|NCI|Rete Ovarii Adenocarcinoma|9110/3
C0025490|T191|PT|BBS2.|RCD|Malignant mesonephroma|9110/3
C0025490|T191|SY|BBS2.|RCD|Mesonephric adenocarcinoma|9110/3
C0025490|T191|PT|BBS..|RCD|Mesonephroma|9110/3
C0025490|T191|SY|BBS2.|RCD|Wolffian duct carcinoma|9110/3
C0025490|T191|OP|BBSz.|RCDSY|Mesonephroma NOS|9110/3
C3840223|T191|PT|703655009|SNOMEDCT_US|Adenocarcinoma of rete ovarii|9110/3
C0025490|T191|SY|2221008|SNOMEDCT_US|Malignant mesonephroma|9110/3
C0025490|T191|SY|2221008|SNOMEDCT_US|Mesonephric adenocarcinoma|9110/3
C0025490|T191|IS|2221008|SNOMEDCT_US|Mesonephroma|9110/3
C0025490|T191|PT|2221008|SNOMEDCT_US|Mesonephroma, malignant|9110/3
C0025490|T191|IS|2221008|SNOMEDCT_US|Mesonephroma, NOS|9110/3
C0025490|T191|SY|2221008|SNOMEDCT_US|Wolffian duct carcinoma|9110/3
C0018916|T191|ET|0000004564|AOD|hemangioma|9120/0
C0018916|T191|PT|0053526|CCPSS|HEMANGIOMA|9120/0
C0018916|T191|PT|0000037071|CHV|benign hemangioma|9120/0
C0018916|T191|SY|0000037071|CHV|benign hemangiomas|9120/0
C0677608|T191|PT|0000042638|CHV|chorioangioma|9120/0
C0677608|T191|SY|0000042638|CHV|chorioangiomas|9120/0
C0018916|T191|SY|0000005936|CHV|haemangioma|9120/0
C0018916|T191|SY|0000058170|CHV|haemangioma|9120/0
C0018916|T191|SY|0000005936|CHV|haemangiomas|9120/0
C0018916|T191|SY|0000058170|CHV|haemangiomas|9120/0
C0018916|T191|PT|0000058170|CHV|hemangioma|9120/0
C0018916|T191|PT|0000005936|CHV|hemangioma|9120/0
C0018916|T191|SY|0000005936|CHV|hemangiomas|9120/0
C0677608|T191|SY|0000042638|CHV|placental chorioangioma|9120/0
C0018916|T191|PT|349|COSTAR|HEMANGIOMA|9120/0
C0018916|T191|PT|2007-1757|CSP|hemangioma|9120/0
C0018916|T191|GT|ANOMALY VASCUL|CST|HEMANGIOMA|9120/0
C0018916|T191|FI|U001925|DXP|HEMANGIOMA|9120/0
C0677608|T191|PT|HP:0100883|HPO|Chorangioma|9120/0
C0018916|T191|PT|HP:0001028|HPO|Hemangioma|9120/0
C0018916|T191|ET|HP:0001028|HPO|Hemangiomata|9120/0
C0677608|T191|SY|HP:0100883|HPO|Placental hamartoma|9120/0
C0018916|T191|SY|HP:0001028|HPO|Strawberry mark|9120/0
C0018916|T191|PT|D18.0|ICD10|Haemangioma, any site|9120/0
C0018916|T191|PT|D18.0|ICD10AE|Hemangioma, any site|9120/0
C0018916|T191|ET|D18.0|ICD10CM|Angioma NOS|9120/0
C0018916|T191|AB|D18.0|ICD10CM|Hemangioma|9120/0
C0018916|T191|HT|D18.0|ICD10CM|Hemangioma|9120/0
C0018916|T191|PT|D18.00|ICD10CM|Hemangioma unspecified site|9120/0
C0018916|T191|AB|D18.00|ICD10CM|Hemangioma unspecified site|9120/0
C0018916|T191|AB|228.00|ICD9CM|Hemangioma NOS|9120/0
C0018916|T191|PT|228.00|ICD9CM|Hemangioma of unspecified site|9120/0
C0018916|T191|HT|228.0|ICD9CM|Hemangioma, any site|9120/0
C0677608|T191|PT|MTHU006383|ICPC2ICD10ENG|angioma; placenta|9120/0
C0677608|T191|PT|MTHU016399|ICPC2ICD10ENG|chorioangioma|9120/0
C0018916|T191|PT|MTHU033761|ICPC2ICD10ENG|hemangioma|9120/0
C0677608|T191|PT|MTHU059775|ICPC2ICD10ENG|placenta; angioma|9120/0
C0018916|T191|PT|S81009|ICPC2P|Haemangioma|9120/0
C0018916|T191|PTN|S81009|ICPC2P|haemangioma|9120/0
C0018916|T191|OP|K99045|ICPC2P|Haemangioma|9120/0
C0018916|T191|OPN|K99045|ICPC2P|haemangioma|9120/0
C0018916|T191|MTH_PT|S81009|ICPC2P|Hemangioma|9120/0
C0018916|T191|MTH_PTN|S81009|ICPC2P|hemangioma|9120/0
C0018916|T191|MTH_OP|K99045|ICPC2P|Hemangioma|9120/0
C0018916|T191|MTH_OPN|K99045|ICPC2P|hemangioma|9120/0
C0018916|T191|PT|U002126|LCH|Hemangioma|9120/0
C0018916|T191|PT|sh85060117|LCH_NW|Hemangiomas|9120/0
C0018916|T191|LPN|LP266918-4|LNC|Hemangioma|9120/0
C0018916|T191|PT|10018814|MDR|Haemangioma|9120/0
C0018916|T191|LLT|10018814|MDR|Haemangioma|9120/0
C0018916|T191|LLT|10018819|MDR|Haemangioma NOS|9120/0
C0018916|T191|LLT|10055903|MDR|Haemangioma of unspecified site|9120/0
C0018916|T191|OL|10018824|MDR|Haemangioma, any site|9120/0
C0018916|T191|LLT|10019386|MDR|Hemangioma|9120/0
C0018916|T191|MTH_PT|10018814|MDR|Hemangioma|9120/0
C0018916|T191|LLT|10019393|MDR|Hemangioma NOS|9120/0
C0018916|T191|LLT|10019401|MDR|Hemangioma of unspecified site|9120/0
C0018916|T191|MTH_OL|10018824|MDR|Hemangioma, any site|9120/0
C0018916|T191|OL|10019405|MDR|Hemangioma, any site|9120/0
C0677608|T191|LLT|10056718|MDR|Placental chorioangioma|9120/0
C0677608|T191|PT|10056718|MDR|Placental chorioangioma|9120/0
C0018916|T191|PT|97903|MEDCIN|hemangioma|9120/0
C0018916|T191|PT|10395|MEDCIN|hemangioma|9120/0
C0018916|T191|SY|5402|MEDLINEPLUS|Hemangioma|9120/0
C0018916|T191|ET|3585|MEDLINEPLUS|Hemangioma|9120/0
C0018916|T191|ET|5402|MEDLINEPLUS|Hemangioma|9120/0
C0018916|T191|ET|533|MEDLINEPLUS|Hemangioma|9120/0
C0677608|T191|ET|D006391|MSH|Chorangioma|9120/0
C0677608|T191|PM|D006391|MSH|Chorangiomas|9120/0
C0677608|T191|PEP|D006391|MSH|Chorioangioma|9120/0
C0677608|T191|PM|D006391|MSH|Chorioangiomas|9120/0
C0018916|T191|MH|D006391|MSH|Hemangioma|9120/0
C0018916|T191|PM|D006391|MSH|Hemangiomas|9120/0
C0677608|T191|PN|NOCODE|MTH|Chorioangioma|9120/0
C0018916|T191|PN|NOCODE|MTH|Hemangioma|9120/0
C0018916|T191|SY|C3085|NCI|Angioma|9120/0
C0677608|T191|SY|C4868|NCI|Angioma of Placenta|9120/0
C0677608|T191|SY|C4868|NCI|Angioma of the Placenta|9120/0
C0018916|T191|SY|C3085|NCI|Benign Angioma|9120/0
C0018916|T191|SY|C3085|NCI|Benign Hemangioma|9120/0
C0677608|T191|SY|C4868|NCI|Chorangioma|9120/0
C0677608|T191|SY|C4868|NCI|Chorangioma of the Placenta|9120/0
C0677608|T191|SY|C4868|NCI|Chorangioma Placentae|9120/0
C0677608|T191|SY|C4868|NCI|Chorioangioma|9120/0
C0018916|T191|PT|C3085|NCI|Hemangioma|9120/0
C0677608|T191|SY|C4868|NCI|Hemangioma of Placenta|9120/0
C0677608|T191|SY|C4868|NCI|Hemangioma of the Placenta|9120/0
C0677608|T191|SY|C4868|NCI|Placental Angioma|9120/0
C0677608|T191|PT|C4868|NCI|Placental Hemangioma|9120/0
C0018916|T191|SY|C3085|NCI_CDISC|Angioma|9120/0
C0018916|T191|SY|C3085|NCI_CDISC|Benign Angioma|9120/0
C0018916|T191|SY|C3085|NCI_CDISC|Benign Hemangioma|9120/0
C0018916|T191|PT|C3085|NCI_CDISC|HEMANGIOMA, BENIGN|9120/0
C0018916|T191|PT|C3085|NCI_CPTAC|Hemangioma|9120/0
C0018916|T191|DN|C3085|NCI_CTRP|Hemangioma|9120/0
C0677608|T191|PT|C4868|NCI_NICHD|Chorangioma|9120/0
C0677608|T191|SY|C4868|NCI_NICHD|Chorangioma of the Placenta|9120/0
C0677608|T191|SY|C4868|NCI_NICHD|Chorangioma Placentae|9120/0
C0677608|T191|SY|C4868|NCI_NICHD|Chorioangioma|9120/0
C0018916|T191|PT|C3085|NCI_NICHD|Hemangioma|9120/0
C0677608|T191|SY|C4868|NCI_NICHD|Placental Hemangioma|9120/0
C0018916|T191|SY|CDR0000665618|PDQ|Benign Angioma|9120/0
C0018916|T191|SY|CDR0000665618|PDQ|Benign Hemangioma|9120/0
C0018916|T191|PT|CDR0000665618|PDQ|hemangioma|9120/0
C0018916|T191|SY|XE1wE|RCD|Angioma|9120/0
C0018916|T191|OP|X78VN|RCD|Angioma - benign|9120/0
C0018916|T191|PT|X77p0|RCD|Benign haemangioma|9120/0
C0677608|T191|PT|X40Bl|RCD|Chorioangioma|9120/0
C0018916|T191|PT|XE1wE|RCD|Haemangioma|9120/0
C0018916|T191|PT|XaBBE|RCD|Haemangioma - morphology|9120/0
C0018916|T191|OP|B7J0z|RCD|Haemangioma NOS|9120/0
C0018916|T191|OP|B7J00|RCD|Haemangioma of unspecified site|9120/0
C0018916|T191|OA|B7J00|RCD|Haemangioma unspecified site|9120/0
C0018916|T191|PT|X77p0|RCDAE|Benign hemangioma|9120/0
C0018916|T191|PT|XE1wE|RCDAE|Hemangioma|9120/0
C0018916|T191|PT|XaBBE|RCDAE|Hemangioma - morphology|9120/0
C0018916|T191|OP|B7J0z|RCDAE|Hemangioma NOS|9120/0
C0018916|T191|OP|B7J00|RCDAE|Hemangioma of unspecified site|9120/0
C0018916|T191|OA|B7J00|RCDAE|Hemangioma unspecified site|9120/0
C0018916|T191|OP|BBT0.|RCDSA|Hemangioma NOS|9120/0
C0018916|T191|OP|BBT0.|RCDSY|Haemangioma NOS|9120/0
C0018916|T191|SY|2099007|SNOMEDCT_US|Angioma|9120/0
C0018916|T191|OAS|154625006|SNOMEDCT_US|Angioma|9120/0
C0018916|T191|OAS|269646001|SNOMEDCT_US|Angioma|9120/0
C0018916|T191|OAP|254822005|SNOMEDCT_US|Angioma - benign|9120/0
C0018916|T191|OAS|189192007|SNOMEDCT_US|Angioma - benign|9120/0
C0018916|T191|IS|2099007|SNOMEDCT_US|Angioma, NOS|9120/0
C0018916|T191|PTGB|253053003|SNOMEDCT_US|Benign haemangioma|9120/0
C0018916|T191|PT|253053003|SNOMEDCT_US|Benign hemangioma|9120/0
C0677608|T191|SY|237268002|SNOMEDCT_US|Chorangioma|9120/0
C0677608|T191|PT|699948001|SNOMEDCT_US|Chorangioma|9120/0
C0677608|T191|SY|2099007|SNOMEDCT_US|Chorioangioma|9120/0
C0677608|T191|PT|237268002|SNOMEDCT_US|Chorioangioma|9120/0
C0677608|T191|SY|699948001|SNOMEDCT_US|Chorioangioma|9120/0
C0018916|T191|OAP|367337005|SNOMEDCT_US|Haemangioma|9120/0
C0018916|T191|OAS|269646001|SNOMEDCT_US|Haemangioma|9120/0
C0018916|T191|OAS|189193002|SNOMEDCT_US|Haemangioma|9120/0
C0018916|T191|PTGB|400210000|SNOMEDCT_US|Haemangioma|9120/0
C0018916|T191|OAS|154625006|SNOMEDCT_US|Haemangioma|9120/0
C0018916|T191|PTGB|2099007|SNOMEDCT_US|Haemangioma|9120/0
C0018916|T191|OF|367337005|SNOMEDCT_US|Haemangioma|9120/0
C0018916|T191|SYGB|2099007|SNOMEDCT_US|Haemangioma - morphology|9120/0
C0018916|T191|OAP|189199003|SNOMEDCT_US|Haemangioma NOS|9120/0
C0018916|T191|OAP|189194008|SNOMEDCT_US|Haemangioma of unspecified site|9120/0
C0018916|T191|OAP|93474003|SNOMEDCT_US|Haemangioma of unspecified site|9120/0
C0018916|T191|IS|2099007|SNOMEDCT_US|Haemangioma, NOS|9120/0
C0018916|T191|IS|2099007|SNOMEDCT_US|Haemangioma, site unspecified|9120/0
C0018916|T191|OAP|367337005|SNOMEDCT_US|Hemangioma|9120/0
C0018916|T191|OAS|154625006|SNOMEDCT_US|Hemangioma|9120/0
C0018916|T191|PT|2099007|SNOMEDCT_US|Hemangioma|9120/0
C0018916|T191|OAS|189193002|SNOMEDCT_US|Hemangioma|9120/0
C0018916|T191|PT|400210000|SNOMEDCT_US|Hemangioma|9120/0
C0018916|T191|OAS|269646001|SNOMEDCT_US|Hemangioma|9120/0
C0018916|T191|SY|2099007|SNOMEDCT_US|Hemangioma - morphology|9120/0
C0018916|T191|OAP|189199003|SNOMEDCT_US|Hemangioma NOS|9120/0
C0018916|T191|OAP|93474003|SNOMEDCT_US|Hemangioma of unspecified site|9120/0
C0018916|T191|OAP|189194008|SNOMEDCT_US|Hemangioma of unspecified site|9120/0
C0018916|T191|SY|2099007|SNOMEDCT_US|Hemangioma, no ICD-O subtype|9120/0
C0018916|T191|SY|2099007|SNOMEDCT_US|Hemangioma, no International Classification of Diseases for Oncology subtype|9120/0
C0018916|T191|IS|2099007|SNOMEDCT_US|Hemangioma, NOS|9120/0
C0018916|T191|IS|2099007|SNOMEDCT_US|Hemangioma, site unspecified|9120/0
C1304507|T191|PTGB|699606005|SNOMEDCT_US|Sinusoidal haemangioma|9120/0
C1304507|T191|PTGB|403965008|SNOMEDCT_US|Sinusoidal haemangioma|9120/0
C1304507|T191|PT|699606005|SNOMEDCT_US|Sinusoidal hemangioma|9120/0
C1304507|T191|PT|403965008|SNOMEDCT_US|Sinusoidal hemangioma|9120/0
C0018923|T191|ET|0000004565|AOD|angiosarcoma|9120/3
C0018923|T191|NP|0000023030|AOD|malignant hemangioendothelioma|9120/3
C0018923|T191|PT|0000005940|CHV|angiosarcoma|9120/3
C0018923|T191|SY|0000005940|CHV|angiosarcomas|9120/3
C0018923|T191|SY|0000005940|CHV|haemangiosarcoma|9120/3
C0018923|T191|SY|0000005940|CHV|hemangiosarcoma|9120/3
C0018923|T191|SY|0000005940|CHV|hemangiosarcomas|9120/3
C0018923|T191|PT|NOCODE|COSTAR|Hemangiosarcoma|9120/3
C0018923|T191|PT|2007-1041|CSP|angiosarcoma|9120/3
C0018923|T191|ET|2007-1041|CSP|hemangiosarcoma|9120/3
C0018923|T191|PT|HP:0200058|HPO|Angiosarcoma|9120/3
C0018923|T191|PT|sh85005032|LCH_NW|Angiosarcoma|9120/3
C0018923|T191|LA|LA26515-9|LNC|Angiosarcoma|9120/3
C0018923|T191|LLT|10002476|MDR|Angiosarcoma|9120/3
C0018923|T191|PT|10002476|MDR|Angiosarcoma|9120/3
C0018923|T191|LLT|10002479|MDR|Angiosarcoma NOS|9120/3
C0018923|T191|LLT|10050367|MDR|Haemangioendothelioma malignant|9120/3
C0018923|T191|LLT|10018827|MDR|Haemangiosarcoma|9120/3
C0018923|T191|LLT|10018828|MDR|Haemangiosarcoma NOS|9120/3
C0018923|T191|LLT|10060540|MDR|Hemangioendothelioma malignant|9120/3
C0018923|T191|LLT|10019407|MDR|Hemangiosarcoma|9120/3
C0018923|T191|MTH_LLT|10018828|MDR|Hemangiosarcoma NOS|9120/3
C0018923|T191|PT|36080|MEDCIN|angiosarcoma|9120/3
C0018923|T191|PT|271555|MEDCIN|malignant hemangioendothelioma|9120/3
C0018923|T191|ET|D006394|MSH|Angiosarcoma|9120/3
C0018923|T191|PM|D006394|MSH|Angiosarcomas|9120/3
C0018923|T191|MH|D006394|MSH|Hemangiosarcoma|9120/3
C0018923|T191|PM|D006394|MSH|Hemangiosarcomas|9120/3
C0018923|T191|PN|NOCODE|MTH|Hemangiosarcoma|9120/3
C0018923|T191|PT|C3088|NCI|Angiosarcoma|9120/3
C0018923|T191|OP|C3088|NCI|Hemangiosarcoma|9120/3
C0018923|T191|OP|C3088|NCI|Malignant Angioendothelioma|9120/3
C0018923|T191|OP|C3088|NCI|Malignant Hemangioendothelioma|9120/3
C0018923|T191|SY|C3088|NCI_CDISC|Hemangiosarcoma|9120/3
C0018923|T191|PT|C3088|NCI_CDISC|HEMANGIOSARCOMA, MALIGNANT|9120/3
C0018923|T191|PT|C3088|NCI_CPTAC|Angiosarcoma|9120/3
C0018923|T191|DN|C3088|NCI_CTRP|Angiosarcoma|9120/3
C0018923|T191|PT|C3088|NCI_CTRP|Angiosarcoma|9120/3
C0018923|T191|PT|CDR0000046532|NCI_NCI-GLOSS|angiosarcoma|9120/3
C0018923|T191|PT|CDR0000335069|NCI_NCI-GLOSS|hemangiosarcoma|9120/3
C0018923|T191|SY|BBT1.|RCD|Angiosarcoma|9120/3
C0018923|T191|SY|BBT71|RCD|Haemangioendothelial sarcoma|9120/3
C0018923|T191|PT|BBT1.|RCD|Haemangiosarcoma|9120/3
C0018923|T191|AB|BBT71|RCD|Malign haemangioendothelioma|9120/3
C0018923|T191|PT|BBT71|RCD|Malignant haemangioendothelioma|9120/3
C0018923|T191|PT|BBT1.|RCDAE|Hemangiosarcoma|9120/3
C0018923|T191|AB|BBT71|RCDAE|Malign hemangioendothelioma|9120/3
C0018923|T191|PT|BBT71|RCDAE|Malignant hemangioendothelioma|9120/3
C0018923|T191|SY|39000009|SNOMEDCT_US|Angiosarcoma|9120/3
C0018923|T191|PT|403977003|SNOMEDCT_US|Angiosarcoma|9120/3
C0018923|T191|SYGB|33176006|SNOMEDCT_US|Haemangioendothelial sarcoma|9120/3
C0018923|T191|PTGB|33176006|SNOMEDCT_US|Haemangioendothelioma, malignant|9120/3
C0018923|T191|PTGB|39000009|SNOMEDCT_US|Haemangiosarcoma|9120/3
C0018923|T191|SY|33176006|SNOMEDCT_US|Hemangioendothelial sarcoma|9120/3
C0018923|T191|PT|33176006|SNOMEDCT_US|Hemangioendothelioma, malignant|9120/3
C0018923|T191|PT|39000009|SNOMEDCT_US|Hemangiosarcoma|9120/3
C0018923|T191|SYGB|403977003|SNOMEDCT_US|Malignant haemangioendothelioma|9120/3
C0018923|T191|SYGB|33176006|SNOMEDCT_US|Malignant haemangioendothelioma|9120/3
C0018923|T191|SY|403977003|SNOMEDCT_US|Malignant hemangioendothelioma|9120/3
C0018923|T191|SY|33176006|SNOMEDCT_US|Malignant hemangioendothelioma|9120/3
C0018920|T191|SY|0000023599|CHV|cavernous haemangioma|9121/0
C0018920|T191|SY|0000005937|CHV|cavernous haemangioma|9121/0
C0018920|T191|SY|0000023599|CHV|cavernous hemangioma|9121/0
C0018920|T191|PT|0000005937|CHV|cavernous hemangioma|9121/0
C0018920|T191|SY|0000005937|CHV|cavernous hemangiomas|9121/0
C0018920|T191|SY|0000005937|CHV|hemangioma cavernous|9121/0
C0018920|T191|PT|NOCODE|COSTAR|Cavernous Hemangioma|9121/0
C0018920|T191|DI|U000784|DXP|HEMANGIOMA, CAVERNOUS|9121/0
C0018920|T191|SY|NOCODE|DXP|HEMANGIOMA, MATURE|9121/0
C0018920|T191|SY|HP:0001048|HPO|Cavernous angioma|9121/0
C0018920|T191|SY|HP:0001048|HPO|Cavernous haemangioma|9121/0
C0018920|T191|PT|HP:0001048|HPO|Cavernous hemangioma|9121/0
C0018920|T191|SY|HP:0001048|HPO|Collection of dilated blood vessels that forms mass|9121/0
C0018920|T191|ET|D18.0|ICD10CM|Cavernous nevus|9121/0
C0018920|T191|PT|MTHU015297|ICPC2ICD10ENG|cavernous; hemangioma|9121/0
C0018920|T191|PT|MTHU015301|ICPC2ICD10ENG|cavernous; nevus|9121/0
C0018920|T191|PT|MTHU033765|ICPC2ICD10ENG|hemangioma; cavernous|9121/0
C0018920|T191|PT|MTHU033762|ICPC2ICD10ENG|hemangioma; strawberry|9121/0
C0018920|T191|PT|MTHU051508|ICPC2ICD10ENG|nevus; cavernous|9121/0
C0018920|T191|PT|MTHU001645|ICPC2ICD10ENG|strawberry; hemangioma|9121/0
C0018920|T191|PTN|S81006|ICPC2P|cavernous naevus|9121/0
C0018920|T191|MTH_PTN|S81006|ICPC2P|cavernous nevus|9121/0
C0018920|T191|PT|S81006|ICPC2P|Naevus;cavernous|9121/0
C0018920|T191|MTH_PT|S81006|ICPC2P|Nevus;cavernous|9121/0
C0018920|T191|LLT|10071746|MDR|Cavernoma|9121/0
C0018920|T191|LLT|10055899|MDR|Haemangioma cavernous|9121/0
C0018920|T191|LLT|10019390|MDR|Hemangioma cavernous|9121/0
C0018920|T191|PT|33261|MEDCIN|cavernous hemangioma|9121/0
C0018920|T191|PT|10399|MEDCIN|cavernous hemangioma|9121/0
C0018920|T191|SY|10399|MEDCIN|hemangioma cavernous|9121/0
C0018920|T191|ET|D006392|MSH|Cavernous Hemangioma|9121/0
C0018920|T191|PM|D006392|MSH|Cavernous Hemangiomas|9121/0
C0018920|T191|MH|D006392|MSH|Hemangioma, Cavernous|9121/0
C0018920|T191|PM|D006392|MSH|Hemangioma, Strawberry|9121/0
C0018920|T191|PM|D006392|MSH|Hemangiomas, Cavernous|9121/0
C0018920|T191|PM|D006392|MSH|Hemangiomas, Strawberry|9121/0
C0018920|T191|PM|D006392|MSH|Strawberry Hemangioma|9121/0
C0018920|T191|ET|D006392|MSH|Strawberry Hemangiomas|9121/0
C0018920|T191|PN|NOCODE|MTH|Hemangioma, Cavernous|9121/0
C0018920|T191|SY|C3086|NCI|Cavernoma|9121/0
C0018920|T191|SY|C3086|NCI|Cavernous Angioma|9121/0
C0018920|T191|PT|C3086|NCI|Cavernous Hemangioma|9121/0
C0018920|T191|SY|PH311|RCD|Cavernous angioma of skin|9121/0
C0018920|T191|SY|PH311|RCD|Cavernous haemangioma|9121/0
C0018920|T191|SY|PH311|RCD|Cavernous naevus|9121/0
C0018920|T191|SY|PH311|RCD|Cavernous naevus of skin|9121/0
C0018920|T191|PT|PH312|RCD|Strawberry haemangioma|9121/0
C0018920|T191|SY|PH311|RCDAE|Cavernous hemangioma|9121/0
C0018920|T191|SY|PH311|RCDAE|Cavernous nevus|9121/0
C0018920|T191|SY|PH311|RCDAE|Cavernous nevus of skin|9121/0
C0018920|T191|PT|PH312|RCDAE|Strawberry hemangioma|9121/0
C0018920|T191|PT|BBT2.|RCDSA|Cavernous hemangioma|9121/0
C0018920|T191|PT|BBT2.|RCDSY|Cavernous haemangioma|9121/0
C0018920|T191|IS|416824008|SNOMEDCT_US|Cavernous angioma of skin|9121/0
C0018920|T191|OAS|67668002|SNOMEDCT_US|Cavernous angioma of skin|9121/0
C0018920|T191|OAS|67668002|SNOMEDCT_US|Cavernous haemangioma|9121/0
C0018920|T191|PTGB|416824008|SNOMEDCT_US|Cavernous haemangioma|9121/0
C0018920|T191|PTGB|33377007|SNOMEDCT_US|Cavernous haemangioma|9121/0
C0018920|T191|PT|416824008|SNOMEDCT_US|Cavernous hemangioma|9121/0
C0018920|T191|PT|33377007|SNOMEDCT_US|Cavernous hemangioma|9121/0
C0018920|T191|OAS|67668002|SNOMEDCT_US|Cavernous hemangioma|9121/0
C0018920|T191|OAS|67668002|SNOMEDCT_US|Cavernous naevus|9121/0
C0018920|T191|OAS|189192007|SNOMEDCT_US|Cavernous naevus|9121/0
C0018920|T191|SYGB|416824008|SNOMEDCT_US|Cavernous naevus|9121/0
C0018920|T191|IS|416824008|SNOMEDCT_US|Cavernous naevus of skin|9121/0
C0018920|T191|OAS|67668002|SNOMEDCT_US|Cavernous naevus of skin|9121/0
C0018920|T191|OAS|67668002|SNOMEDCT_US|Cavernous nevus|9121/0
C0018920|T191|OAS|189192007|SNOMEDCT_US|Cavernous nevus|9121/0
C0018920|T191|SY|416824008|SNOMEDCT_US|Cavernous nevus|9121/0
C0018920|T191|IS|416824008|SNOMEDCT_US|Cavernous nevus of skin|9121/0
C0018920|T191|OAS|67668002|SNOMEDCT_US|Cavernous nevus of skin|9121/0
C0018920|T191|SYGB|56975005|SNOMEDCT_US|Strawberry haemangioma|9121/0
C0018920|T191|OAP|157014007|SNOMEDCT_US|Strawberry haemangioma|9121/0
C0018920|T191|OAP|254781005|SNOMEDCT_US|Strawberry haemangioma|9121/0
C0018920|T191|OF|157014007|SNOMEDCT_US|Strawberry haemangioma|9121/0
C0018920|T191|OF|254781005|SNOMEDCT_US|Strawberry haemangioma|9121/0
C0018920|T191|SY|56975005|SNOMEDCT_US|Strawberry hemangioma|9121/0
C0018920|T191|OAP|157014007|SNOMEDCT_US|Strawberry hemangioma|9121/0
C0018920|T191|OAP|254781005|SNOMEDCT_US|Strawberry hemangioma|9121/0
C0334532|T191|SY|0000030001|CHV|hemangioma venous|9122/0
C0334532|T191|SY|0000030001|CHV|hemangiomas venous|9122/0
C0334532|T191|PT|0000030001|CHV|venous hemangioma|9122/0
C0334532|T191|PT|MTHU033776|ICPC2ICD10ENG|hemangioma; venous|9122/0
C0334532|T191|PT|MTHU079502|ICPC2ICD10ENG|venous; hemangioma|9122/0
C0334532|T191|SY|C4296|NCI|Venous Angioma|9122/0
C0334532|T191|PT|C4296|NCI|Venous Hemangioma|9122/0
C0334532|T191|PT|BBT3.|RCD|Venous haemangioma|9122/0
C0334532|T191|PT|BBT3.|RCDAE|Venous hemangioma|9122/0
C1304506|T191|PTGB|699607001|SNOMEDCT_US|Microvenular haemangioma|9122/0
C1304506|T191|PTGB|403964007|SNOMEDCT_US|Microvenular haemangioma|9122/0
C1304506|T191|PT|699607001|SNOMEDCT_US|Microvenular hemangioma|9122/0
C1304506|T191|PT|403964007|SNOMEDCT_US|Microvenular hemangioma|9122/0
C0334532|T191|PTGB|56468002|SNOMEDCT_US|Venous haemangioma|9122/0
C0334532|T191|PTGB|403968005|SNOMEDCT_US|Venous haemangioma|9122/0
C0334532|T191|PT|56468002|SNOMEDCT_US|Venous hemangioma|9122/0
C0334532|T191|PT|403968005|SNOMEDCT_US|Venous hemangioma|9122/0
C0334533|T191|SY|0000030002|CHV|arterial hemangioma|9123/0
C0334533|T191|SY|0000030002|CHV|arteriovenous haemangioma|9123/0
C0334533|T191|PT|0000030002|CHV|arteriovenous malformation|9123/0
C0334533|T191|SY|0000030002|CHV|arteriovenous malformations|9123/0
C0334533|T191|SY|0000030002|CHV|cirsoid aneurysm|9123/0
C0334533|T191|ET|I77.0|ICD10CM|Aneurysmal varix|9123/0
C0334533|T191|PT|MTHU006287|ICPC2ICD10ENG|aneurysm; racemose|9123/0
C0334533|T191|PT|MTHU006318|ICPC2ICD10ENG|aneurysmal; varix|9123/0
C0334533|T191|PT|MTHU008118|ICPC2ICD10ENG|arteriovenous; hemangioma|9123/0
C0334533|T191|PT|MTHU033763|ICPC2ICD10ENG|hemangioma; arteriovenous|9123/0
C0334533|T191|PT|MTHU033774|ICPC2ICD10ENG|hemangioma; racemose|9123/0
C0334533|T191|PT|MTHU063545|ICPC2ICD10ENG|racemose; aneurysm|9123/0
C0334533|T191|PT|MTHU063544|ICPC2ICD10ENG|racemose; hemangioma|9123/0
C0334533|T191|PT|MTHU079204|ICPC2ICD10ENG|varix; aneurysmal|9123/0
C0334533|T191|LLT|10055898|MDR|Haemangioma arterial|9123/0
C0334533|T191|LLT|10019389|MDR|Hemangioma arterial|9123/0
C0334533|T191|PN|NOCODE|MTH|Arteriovenous hemangioma|9123/0
C0334533|T191|SY|C2882|NCI|Arteriovenous Angioma|9123/0
C0334533|T191|SY|C2882|NCI|Arteriovenous Hemangioma|9123/0
C0334533|T191|PT|C2882|NCI|Arteriovenous Hemangioma/Malformation|9123/0
C0334533|T191|SY|C2882|NCI|Arteriovenous Malformation|9123/0
C0334533|T191|SY|C2882|NCI|Racemose Angioma|9123/0
C0334533|T191|SY|C2882|NCI|Racemose Hemangioma|9123/0
C0334533|T191|PT|C2882|NCI_NICHD|Arteriovenous Hemangioma|9123/0
C0334533|T191|SY|BBT4.|RCD|Arteriovenous haemangioma|9123/0
C0334533|T191|OP|X2049|RCD|Cirsoid aneurysm|9123/0
C0334533|T191|PT|BBT4.|RCD|Racemose haemangioma|9123/0
C0334533|T191|SY|BBT4.|RCDAE|Arteriovenous hemangioma|9123/0
C0334533|T191|PT|BBT4.|RCDAE|Racemose hemangioma|9123/0
C0334533|T191|SY|14156004|SNOMEDCT_US|Aneurysmal varix|9123/0
C0334533|T191|SYGB|11071001|SNOMEDCT_US|Arteriovenous haemangioma|9123/0
C0334533|T191|PTGB|403966009|SNOMEDCT_US|Arteriovenous haemangioma|9123/0
C0334533|T191|PT|403966009|SNOMEDCT_US|Arteriovenous hemangioma|9123/0
C0334533|T191|SY|11071001|SNOMEDCT_US|Arteriovenous hemangioma|9123/0
C0334533|T191|IS|403966009|SNOMEDCT_US|Arteriovenous malformation|9123/0
C0334533|T191|OAS|204480002|SNOMEDCT_US|Cirsoid aneurysm|9123/0
C0334533|T191|PT|233982006|SNOMEDCT_US|Cirsoid aneurysm|9123/0
C0334533|T191|SY|14156004|SNOMEDCT_US|Cirsoid aneurysm|9123/0
C0334533|T191|IS|403966009|SNOMEDCT_US|Cirsoid aneurysm|9123/0
C0334533|T191|SY|14156004|SNOMEDCT_US|Diffuse arterial ectasia|9123/0
C0334533|T191|PT|14156004|SNOMEDCT_US|Racemose aneurysm|9123/0
C0334533|T191|SY|11071001|SNOMEDCT_US|Racemose angioma|9123/0
C0334533|T191|PTGB|11071001|SNOMEDCT_US|Racemose haemangioma|9123/0
C0334533|T191|PT|11071001|SNOMEDCT_US|Racemose hemangioma|9123/0
C0334533|T191|SY|14156004|SNOMEDCT_US|Venous racemose aneurysm|9123/0
C0334534|T191|ET|0000004599|AOD|Kupffer cell sarcoma|9124/3
C0345907|T191|SY|0000031026|CHV|angiosarcoma liver|9124/3
C0345907|T191|PT|0000031026|CHV|angiosarcoma of liver|9124/3
C0345907|T191|PT|C22.3|ICD10|Angiosarcoma of liver|9124/3
C0345907|T191|AB|C22.3|ICD10CM|Angiosarcoma of liver|9124/3
C0345907|T191|PT|C22.3|ICD10CM|Angiosarcoma of liver|9124/3
C0334534|T191|ET|C22.3|ICD10CM|Kupffer cell sarcoma|9124/3
C0345907|T191|PT|MTHU006399|ICPC2ICD10ENG|angiosarcoma; liver|9124/3
C0334534|T191|PT|MTHU042235|ICPC2ICD10ENG|Kupffer cell sarcoma|9124/3
C0334534|T191|PT|MTHU042234|ICPC2ICD10ENG|Kupffer cell; sarcoma|9124/3
C0345907|T191|PT|MTHU044922|ICPC2ICD10ENG|liver; angiosarcoma|9124/3
C0334534|T191|PT|MTHU065917|ICPC2ICD10ENG|sarcoma; Kupffer cell|9124/3
C0345907|T191|LLT|10067388|MDR|Hepatic angiosarcoma|9124/3
C0345907|T191|PT|10067388|MDR|Hepatic angiosarcoma|9124/3
C0345907|T191|PT|353432|MEDCIN|Angiosarcoma of liver|9124/3
C0345907|T191|PT|31586|MEDCIN|hemangiosarcoma of liver|9124/3
C0345907|T191|SY|31586|MEDCIN|hepatic hemangiosarcoma|9124/3
C0345907|T191|SY|353432|MEDCIN|liver neoplasm malignant angiosarcoma|9124/3
C0334534|T191|PN|NOCODE|MTH|Kupffer cell sarcoma|9124/3
C0345907|T191|SY|C4438|NCI|Angiosarcoma of Liver|9124/3
C0345907|T191|SY|C4438|NCI|Angiosarcoma of the Liver|9124/3
C0345907|T191|SY|C4438|NCI|Hemangiosarcoma of Liver|9124/3
C0345907|T191|SY|C4438|NCI|Hemangiosarcoma of the Liver|9124/3
C0345907|T191|SY|C4438|NCI|Hepatic Angiosarcoma|9124/3
C0345907|T191|SY|C4438|NCI|Hepatic Hemangiosarcoma|9124/3
C0345907|T191|PT|C4438|NCI|Liver Angiosarcoma|9124/3
C0345907|T191|SY|C4438|NCI|Liver Hemangiosarcoma|9124/3
C0345907|T191|SY|C4438|NCI|Primary Angiosarcoma of Liver|9124/3
C0345907|T191|SY|C4438|NCI|Primary Angiosarcoma of the Liver|9124/3
C0345907|T191|PT|C4438|NCI_CPTAC|Liver Angiosarcoma|9124/3
C0345907|T191|PT|X78P0|RCD|Angiosarcoma of liver|9124/3
C0334534|T191|PT|BBT5.|RCD|Kupffer cell sarcoma|9124/3
C0345907|T191|SY|X78P0|RCD|Primary angiosarcoma of liver|9124/3
C0345907|T191|OAP|187770005|SNOMEDCT_US|Angiosarcoma of liver|9124/3
C0345907|T191|OF|187770005|SNOMEDCT_US|Angiosarcoma of liver|9124/3
C0345907|T191|PT|109844006|SNOMEDCT_US|Angiosarcoma of liver|9124/3
C0334534|T191|PT|69317001|SNOMEDCT_US|Kupffer cell sarcoma|9124/3
C0345907|T191|SY|109844006|SNOMEDCT_US|Primary angiosarcoma of liver|9124/3
C0205788|T191|SY|HP:0032060|HPO|Angiolymphoid hyperplasia with eosinophilia|9125/0
C0205788|T191|PT|HP:0032060|HPO|Epithelioid hemangioma|9125/0
C0205788|T191|PT|MTHU026832|ICPC2ICD10ENG|epithelioid; hemangioma|9125/0
C0205788|T191|PT|MTHU033767|ICPC2ICD10ENG|hemangioma; epithelioid|9125/0
C0205788|T191|PT|MTHU033768|ICPC2ICD10ENG|hemangioma; histiocytoid|9125/0
C0205788|T191|PT|MTHU035169|ICPC2ICD10ENG|histiocytoid; hemangioma|9125/0
C0205788|T191|LLT|10048637|MDR|Angiolymphoid hyperplasia with eosinophilia|9125/0
C0205788|T191|PT|10048637|MDR|Angiolymphoid hyperplasia with eosinophilia|9125/0
C0205788|T191|PEP|D006391|MSH|Hemangioma, Histiocytoid|9125/0
C0205788|T191|PM|D006391|MSH|Hemangiomas, Histiocytoid|9125/0
C0205788|T191|PM|D006391|MSH|Histiocytoid Hemangioma|9125/0
C0205788|T191|PM|D006391|MSH|Histiocytoid Hemangiomas|9125/0
C0205788|T191|PN|NOCODE|MTH|Histiocytoid hemangioma|9125/0
C0205788|T191|SY|C4298|NCI|Angiolymphoid Hyperplasia with Eosinophilia|9125/0
C0205788|T191|PT|C4298|NCI|Epithelioid Hemangioma|9125/0
C0205788|T191|SY|C4298|NCI|Histiocytoid Hemangioma|9125/0
C0205788|T191|PT|CDR0000779852|PDQ|adult epithelioid hemangioma|9125/0
C0205788|T191|SY|CDR0000779852|PDQ|angiolymphoid hyperplasia with eosinophilia|9125/0
C0205788|T191|SY|CDR0000779852|PDQ|epithelioid hemangioma|9125/0
C0205788|T191|SY|CDR0000779852|PDQ|histiocytoid hemangioma|9125/0
C0205788|T191|PT|X77p1|RCD|Epithelioid haemangioma|9125/0
C0205788|T191|PT|X77p2|RCD|Histiocytoid haemangioma|9125/0
C0205788|T191|PT|X77p1|RCDAE|Epithelioid hemangioma|9125/0
C0205788|T191|PT|X77p2|RCDAE|Histiocytoid hemangioma|9125/0
C0205788|T191|PT|125574005|SNOMEDCT_US|Angiolymphoid hyperplasia with eosinophilia|9125/0
C5230993|T191|PT|817950008|SNOMEDCT_US|Cutaneous epithelioid angiomatoid nodule|9125/0
C5230993|T191|SY|817950008|SNOMEDCT_US|Cutaneous epithelioid angiomatous nodule|9125/0
C0205788|T191|PTGB|33929001|SNOMEDCT_US|Epithelioid haemangioma|9125/0
C0205788|T191|OAP|189869009|SNOMEDCT_US|Epithelioid haemangioma|9125/0
C0205788|T191|OF|189869009|SNOMEDCT_US|Epithelioid haemangioma|9125/0
C0205788|T191|OAP|189869009|SNOMEDCT_US|Epithelioid hemangioma|9125/0
C0205788|T191|PT|33929001|SNOMEDCT_US|Epithelioid hemangioma|9125/0
C0205788|T191|OAP|253054009|SNOMEDCT_US|Histiocytoid haemangioma|9125/0
C0205788|T191|OF|189870005|SNOMEDCT_US|Histiocytoid haemangioma|9125/0
C0205788|T191|SYGB|33929001|SNOMEDCT_US|Histiocytoid haemangioma|9125/0
C0205788|T191|OAP|189870005|SNOMEDCT_US|Histiocytoid haemangioma|9125/0
C0205788|T191|OAP|69159005|SNOMEDCT_US|Histiocytoid haemangioma|9125/0
C0205788|T191|IS|69159005|SNOMEDCT_US|Histiocytoid haemangioma -RETIRED-|9125/0
C0205788|T191|OAP|69159005|SNOMEDCT_US|Histiocytoid hemangioma|9125/0
C0205788|T191|SY|33929001|SNOMEDCT_US|Histiocytoid hemangioma|9125/0
C0205788|T191|OAP|253054009|SNOMEDCT_US|Histiocytoid hemangioma|9125/0
C0205788|T191|OAP|189870005|SNOMEDCT_US|Histiocytoid hemangioma|9125/0
C0205788|T191|OF|69159005|SNOMEDCT_US|Histiocytoid hemangioma -RETIRED-|9125/0
C0205788|T191|IS|69159005|SNOMEDCT_US|Histiocytoid hemangioma -RETIRED-|9125/0
C0334536|T191|PT|MTHU006360|ICPC2ICD10ENG|angioendothelioma; benign|9130/0
C0334536|T191|PT|MTHU010308|ICPC2ICD10ENG|benign; angioendothelioma|9130/0
C0334536|T191|PT|MTHU010314|ICPC2ICD10ENG|benign; hemangioendothelioma|9130/0
C0334536|T191|PT|MTHU033757|ICPC2ICD10ENG|hemangioendothelioma; benign|9130/0
C0334539|T191|PT|MTHU040141|ICPC2ICD10ENG|intravascular; bronchial alveolar tumor|9130/0
C0334539|T191|PT|MTHU077075|ICPC2ICD10ENG|tumor; intravascular bronchial alveolar|9130/0
C0334536|T191|OP|C66779|NCI|Benign Hemangioendothelioma|9130/0
C0334536|T191|PT|C66779|NCI|Benign Hemangioendothelioma|9130/0
C0334536|T191|PT|BBT70|RCD|Benign haemangioendothelioma|9130/0
C0334539|T191|AB|X77p5|RCD|Intravasc bronchial alveol tum|9130/0
C0334539|T191|PT|X77p5|RCD|Intravascular bronchial alveolar tumour|9130/0
C0334536|T191|PT|BBT70|RCDAE|Benign hemangioendothelioma|9130/0
C0334539|T191|PT|X77p5|RCDAE|Intravascular bronchial alveolar tumor|9130/0
C0334539|T191|AB|X77p5|RCDSY|Intravas bronch alveol tumr|9130/0
C0334536|T191|SYGB|31104000|SNOMEDCT_US|Benign haemangioendothelioma|9130/0
C0334536|T191|SY|31104000|SNOMEDCT_US|Benign hemangioendothelioma|9130/0
C0334536|T191|PTGB|31104000|SNOMEDCT_US|Haemangioendothelioma, benign|9130/0
C0334536|T191|PT|31104000|SNOMEDCT_US|Hemangioendothelioma, benign|9130/0
C0334539|T191|OAP|189873007|SNOMEDCT_US|Intravascular bronchial alveolar tumor|9130/0
C0334539|T191|OAP|85170001|SNOMEDCT_US|Intravascular bronchial alveolar tumor|9130/0
C0334539|T191|PT|253055005|SNOMEDCT_US|Intravascular bronchial alveolar tumor|9130/0
C0334539|T191|IS|85170001|SNOMEDCT_US|Intravascular bronchial alveolar tumor -RETIRED-|9130/0
C0334539|T191|OF|85170001|SNOMEDCT_US|Intravascular bronchial alveolar tumor -RETIRED-|9130/0
C0334539|T191|OAP|189873007|SNOMEDCT_US|Intravascular bronchial alveolar tumour|9130/0
C0334539|T191|OAP|85170001|SNOMEDCT_US|Intravascular bronchial alveolar tumour|9130/0
C0334539|T191|OF|189873007|SNOMEDCT_US|Intravascular bronchial alveolar tumour|9130/0
C0334539|T191|PTGB|253055005|SNOMEDCT_US|Intravascular bronchial alveolar tumour|9130/0
C0334539|T191|IS|85170001|SNOMEDCT_US|Intravascular bronchial alveolar tumour -RETIRED-|9130/0
C0018915|T191|NP|0000023029|AOD|hemangioendothelioma|9130/1
C0018915|T191|SY|0000005935|CHV|haemangioendothelioma|9130/1
C0018915|T191|PT|0000005935|CHV|hemangioendothelioma|9130/1
C0018915|T191|SY|0000005935|CHV|hemangioendotheliomas|9130/1
C0018915|T191|ET|2007-1757|CSP|hemangioendothelioma|9130/1
C0018915|T191|ET|2007-1757|CSP|vascular endothelioma|9130/1
C0018915|T191|PT|MTHU006359|ICPC2ICD10ENG|angioendothelioma|9130/1
C0018915|T191|PT|355050|MEDCIN|hemangioendothelioma|9130/1
C0018915|T191|SY|355050|MEDCIN|neoplasm - soft tissue types blood vessel hemangioendothelioma|9130/1
C0018915|T191|ET|D006390|MSH|Endothelioma, Vascular|9130/1
C0018915|T191|PM|D006390|MSH|Endotheliomas, Vascular|9130/1
C0018915|T191|PM|D006390|MSH|Hemangio Endothelioma|9130/1
C0018915|T191|ET|D006390|MSH|Hemangio-Endothelioma|9130/1
C0018915|T191|PM|D006390|MSH|Hemangio-Endotheliomas|9130/1
C0018915|T191|MH|D006390|MSH|Hemangioendothelioma|9130/1
C0018915|T191|PM|D006390|MSH|Hemangioendotheliomas|9130/1
C0018915|T191|PM|D006390|MSH|Vascular Endothelioma|9130/1
C0018915|T191|PM|D006390|MSH|Vascular Endotheliomas|9130/1
C0018915|T191|SY|C3084|NCI|Angioendothelioma|9130/1
C0018915|T191|PT|C3084|NCI|Hemangioendothelioma|9130/1
C0018915|T191|PT|C3084|NCI_NICHD|Hemangioendothelioma|9130/1
C0018915|T191|SY|BBT7.|RCD|Angioendothelioma|9130/1
C0018915|T191|SY|BBT7.|RCD|Haemangioendothelioma|9130/1
C0018915|T191|SY|BBT7.|RCDAE|Hemangioendothelioma|9130/1
C0018915|T191|OP|BBT7z|RCDSA|Hemangioendothelioma NOS|9130/1
C0018915|T191|OP|BBT7z|RCDSY|Haemangioendothelioma NOS|9130/1
C0018915|T191|SY|66229009|SNOMEDCT_US|Angioendothelioma|9130/1
C0018915|T191|PTGB|66229009|SNOMEDCT_US|Haemangioendothelioma|9130/1
C0018915|T191|PTGB|403980002|SNOMEDCT_US|Haemangioendothelioma|9130/1
C0018915|T191|IS|66229009|SNOMEDCT_US|Haemangioendothelioma, NOS|9130/1
C0018915|T191|PT|66229009|SNOMEDCT_US|Hemangioendothelioma|9130/1
C0018915|T191|PT|403980002|SNOMEDCT_US|Hemangioendothelioma|9130/1
C0018915|T191|IS|66229009|SNOMEDCT_US|Hemangioendothelioma, NOS|9130/1
C2959809|T191|PTGB|447203005|SNOMEDCT_US|Infantile haemangioendothelioma, type I|9130/1
C2959809|T191|PT|447203005|SNOMEDCT_US|Infantile hemangioendothelioma, type I|9130/1
C0018923|T191|ET|0000004565|AOD|angiosarcoma|9130/3
C0018923|T191|NP|0000023030|AOD|malignant hemangioendothelioma|9130/3
C0018923|T191|PT|0000005940|CHV|angiosarcoma|9130/3
C0018923|T191|SY|0000005940|CHV|angiosarcomas|9130/3
C0206732|T191|PT|0000021056|CHV|epithelioid hemangioendothelioma|9130/3
C0018923|T191|SY|0000005940|CHV|haemangiosarcoma|9130/3
C0018923|T191|SY|0000005940|CHV|hemangiosarcoma|9130/3
C0018923|T191|SY|0000005940|CHV|hemangiosarcomas|9130/3
C0018923|T191|PT|NOCODE|COSTAR|Hemangiosarcoma|9130/3
C0018923|T191|PT|2007-1041|CSP|angiosarcoma|9130/3
C0018923|T191|ET|2007-1041|CSP|hemangiosarcoma|9130/3
C0018923|T191|PT|HP:0200058|HPO|Angiosarcoma|9130/3
C0018923|T191|PT|sh85005032|LCH_NW|Angiosarcoma|9130/3
C0018923|T191|LA|LA26515-9|LNC|Angiosarcoma|9130/3
C0018923|T191|LLT|10002476|MDR|Angiosarcoma|9130/3
C0018923|T191|PT|10002476|MDR|Angiosarcoma|9130/3
C0018923|T191|LLT|10002479|MDR|Angiosarcoma NOS|9130/3
C0206732|T191|LLT|10079874|MDR|Epithelioid haemangioendothelioma|9130/3
C0206732|T191|LLT|10079873|MDR|Epithelioid hemangioendothelioma|9130/3
C0018923|T191|LLT|10050367|MDR|Haemangioendothelioma malignant|9130/3
C0018923|T191|LLT|10018827|MDR|Haemangiosarcoma|9130/3
C0018923|T191|LLT|10018828|MDR|Haemangiosarcoma NOS|9130/3
C0018923|T191|LLT|10060540|MDR|Hemangioendothelioma malignant|9130/3
C0018923|T191|LLT|10019407|MDR|Hemangiosarcoma|9130/3
C0018923|T191|MTH_LLT|10018828|MDR|Hemangiosarcoma NOS|9130/3
C0018923|T191|PT|36080|MEDCIN|angiosarcoma|9130/3
C0206732|T191|PT|355058|MEDCIN|epithelioid hemangioendothelioma|9130/3
C0018923|T191|PT|271555|MEDCIN|malignant hemangioendothelioma|9130/3
C0206732|T191|SY|355058|MEDCIN|neoplasm - soft tissue blood vessel hemangioendothelioma epithelioid|9130/3
C0018923|T191|ET|D006394|MSH|Angiosarcoma|9130/3
C0018923|T191|PM|D006394|MSH|Angiosarcomas|9130/3
C0206732|T191|PM|D018323|MSH|Epithelioid Hemangioendothelioma|9130/3
C0206732|T191|PM|D018323|MSH|Epithelioid Hemangioendotheliomas|9130/3
C0206732|T191|MH|D018323|MSH|Hemangioendothelioma, Epithelioid|9130/3
C0206732|T191|PM|D018323|MSH|Hemangioendotheliomas, Epithelioid|9130/3
C0018923|T191|MH|D006394|MSH|Hemangiosarcoma|9130/3
C0018923|T191|PM|D006394|MSH|Hemangiosarcomas|9130/3
C0206732|T191|PN|NOCODE|MTH|Epithelioid hemangioendothelioma|9130/3
C0018923|T191|PN|NOCODE|MTH|Hemangiosarcoma|9130/3
C0018923|T191|PT|C3088|NCI|Angiosarcoma|9130/3
C0206732|T191|SY|C3800|NCI|Epithelioid Angioendothelioma|9130/3
C0206732|T191|SY|C3800|NCI|Epithelioid Angiosarcoma|9130/3
C0206732|T191|PT|C3800|NCI|Epithelioid Hemangioendothelioma|9130/3
C0018923|T191|OP|C3088|NCI|Hemangiosarcoma|9130/3
C0018923|T191|OP|C3088|NCI|Malignant Angioendothelioma|9130/3
C0018923|T191|OP|C3088|NCI|Malignant Hemangioendothelioma|9130/3
C0018923|T191|SY|C3088|NCI_CDISC|Hemangiosarcoma|9130/3
C0018923|T191|PT|C3088|NCI_CDISC|HEMANGIOSARCOMA, MALIGNANT|9130/3
C0018923|T191|PT|C3088|NCI_CPTAC|Angiosarcoma|9130/3
C0018923|T191|DN|C3088|NCI_CTRP|Angiosarcoma|9130/3
C0018923|T191|PT|C3088|NCI_CTRP|Angiosarcoma|9130/3
C0018923|T191|PT|CDR0000046532|NCI_NCI-GLOSS|angiosarcoma|9130/3
C0018923|T191|PT|CDR0000335069|NCI_NCI-GLOSS|hemangiosarcoma|9130/3
C0018923|T191|SY|BBT1.|RCD|Angiosarcoma|9130/3
C0206732|T191|AB|X77p4|RCD|Epithel haemangioendothelioma|9130/3
C0206732|T191|PT|X77p4|RCD|Epithelioid haemangioendothelioma|9130/3
C0018923|T191|SY|BBT71|RCD|Haemangioendothelial sarcoma|9130/3
C0018923|T191|PT|BBT1.|RCD|Haemangiosarcoma|9130/3
C0018923|T191|AB|BBT71|RCD|Malign haemangioendothelioma|9130/3
C0018923|T191|PT|BBT71|RCD|Malignant haemangioendothelioma|9130/3
C0206732|T191|AB|X77p4|RCDAE|Epithel hemangioendothelioma|9130/3
C0206732|T191|PT|X77p4|RCDAE|Epithelioid hemangioendothelioma|9130/3
C0018923|T191|PT|BBT1.|RCDAE|Hemangiosarcoma|9130/3
C0018923|T191|AB|BBT71|RCDAE|Malign hemangioendothelioma|9130/3
C0018923|T191|PT|BBT71|RCDAE|Malignant hemangioendothelioma|9130/3
C0206732|T191|OP|BBTJ.|RCDSA|Epithelioid hemangioendothelioma NOS|9130/3
C0206732|T191|OA|BBTJ.|RCDSY|Epithe haemngioendothelioma|9130/3
C0206732|T191|OP|BBTJ.|RCDSY|Epithelioid haemangioendothelioma NOS|9130/3
C0018923|T191|PT|403977003|SNOMEDCT_US|Angiosarcoma|9130/3
C0018923|T191|SY|39000009|SNOMEDCT_US|Angiosarcoma|9130/3
C0206732|T191|OAP|84290008|SNOMEDCT_US|Epithelioid haemangioendothelioma|9130/3
C0206732|T191|PTGB|403981003|SNOMEDCT_US|Epithelioid haemangioendothelioma|9130/3
C0206732|T191|OAP|84290008|SNOMEDCT_US|Epithelioid hemangioendothelioma|9130/3
C0206732|T191|PT|403981003|SNOMEDCT_US|Epithelioid hemangioendothelioma|9130/3
C0206732|T191|IS|84290008|SNOMEDCT_US|Epithelioid hemangioendothelioma, NOS|9130/3
C0018923|T191|SYGB|33176006|SNOMEDCT_US|Haemangioendothelial sarcoma|9130/3
C0018923|T191|PTGB|33176006|SNOMEDCT_US|Haemangioendothelioma, malignant|9130/3
C0018923|T191|PTGB|39000009|SNOMEDCT_US|Haemangiosarcoma|9130/3
C0018923|T191|SY|33176006|SNOMEDCT_US|Hemangioendothelial sarcoma|9130/3
C0018923|T191|PT|33176006|SNOMEDCT_US|Hemangioendothelioma, malignant|9130/3
C0018923|T191|PT|39000009|SNOMEDCT_US|Hemangiosarcoma|9130/3
C0018923|T191|SYGB|403977003|SNOMEDCT_US|Malignant haemangioendothelioma|9130/3
C0018923|T191|SYGB|33176006|SNOMEDCT_US|Malignant haemangioendothelioma|9130/3
C0018923|T191|SY|403977003|SNOMEDCT_US|Malignant hemangioendothelioma|9130/3
C0018923|T191|SY|33176006|SNOMEDCT_US|Malignant hemangioendothelioma|9130/3
C0085653|T191|PT|1009419|CCPSS|GRANULOMA PYOGENIC|9131/0
C0206733|T191|SY|0000021057|CHV|angiomas strawberry|9131/0
C0206733|T191|SY|0000021057|CHV|birthmarks strawberry|9131/0
C0206733|T191|SY|0000015722|CHV|capillary angioma|9131/0
C0206733|T191|SY|0000021057|CHV|capillary haemangioma|9131/0
C0206733|T191|PT|0000021057|CHV|capillary hemangioma|9131/0
C0206733|T191|SY|0000021057|CHV|capillary hemangiomas|9131/0
C0085653|T191|SY|0000015711|CHV|capillary lobular hemangioma|9131/0
C0085653|T191|SY|0000015711|CHV|granuloma pyogenic|9131/0
C0085653|T191|SY|0000015711|CHV|granuloma pyogenicum|9131/0
C0085653|T191|SY|0000015711|CHV|granulomas pyogenic|9131/0
C0206733|T191|SY|0000021057|CHV|hemangioma simplex|9131/0
C0206733|T191|SY|0000021057|CHV|hemangioma strawberry|9131/0
C0206733|T191|SY|0000021057|CHV|hemangiomas infantile|9131/0
C0206733|T191|SY|0000021057|CHV|hemangiomas strawberry|9131/0
C0206733|T191|SY|0000021057|CHV|infantile hemangioma|9131/0
C0206733|T191|SY|0000021057|CHV|juvenile hemangioma|9131/0
C0085653|T191|SY|0000015711|CHV|lobular capillary hemangioma|9131/0
C0206733|T191|SY|0000021057|CHV|mark strawberry|9131/0
C0206733|T191|SY|0000021057|CHV|marks strawberry|9131/0
C0206733|T191|SY|0000021057|CHV|nevus capillary|9131/0
C0206733|T191|SY|0000021057|CHV|plexiform hemangioma|9131/0
C0085653|T191|PT|0000015711|CHV|pyogenic granuloma|9131/0
C0206733|T191|SY|0000021057|CHV|strawberry angioma|9131/0
C0206733|T191|SY|0000021057|CHV|strawberry birthmark|9131/0
C0206733|T191|SY|0000021057|CHV|strawberry hemangioma|9131/0
C0206733|T191|SY|0000021057|CHV|strawberry mark|9131/0
C0206733|T191|SY|0000021057|CHV|strawberry naevus|9131/0
C0206733|T191|SY|0000021057|CHV|strawberry nevus|9131/0
C0206733|T191|PT|NOCODE|COSTAR|Capillary Hemangioma|9131/0
C0085653|T191|PT|U000575|COSTAR|PYOGENIC GRANULOMA|9131/0
C0206733|T191|GT|ANOMALY VASCUL|CST|STRAWBERRY MARK|9131/0
C0206733|T191|SY|HP:0005306|HPO|Capillary hemangioma|9131/0
C0206733|T191|PT|HP:0005306|HPO|Capillary hemangioma|9131/0
C0206733|T191|SY|HP:0005306|HPO|Strawberry birthmark|9131/0
C0085653|T191|ET|K13.4|ICD10CM|Granuloma pyogenicum|9131/0
C0206733|T191|ET|Q82.5|ICD10CM|Strawberry Nevus|9131/0
C0206733|T191|PT|MTHU006372|ICPC2ICD10ENG|angiomatous; nevus|9131/0
C0206733|T191|PT|MTHU014660|ICPC2ICD10ENG|capillary; hemangioma|9131/0
C0206733|T191|PT|MTHU014663|ICPC2ICD10ENG|capillary; nevus|9131/0
C0085653|T191|PT|MTHU032806|ICPC2ICD10ENG|granuloma; pyogenic|9131/0
C0085653|T191|PT|MTHU032824|ICPC2ICD10ENG|granuloma; telangiectaticum|9131/0
C0206733|T191|PT|MTHU033764|ICPC2ICD10ENG|hemangioma; capillary|9131/0
C0206733|T191|PT|MTHU033769|ICPC2ICD10ENG|hemangioma; infantile|9131/0
C0206733|T191|PT|MTHU033771|ICPC2ICD10ENG|hemangioma; juvenile|9131/0
C0206733|T191|PT|MTHU033773|ICPC2ICD10ENG|hemangioma; plexiform|9131/0
C0206733|T191|PT|MTHU033775|ICPC2ICD10ENG|hemangioma; simplex|9131/0
C0206733|T191|PT|MTHU037880|ICPC2ICD10ENG|infantile; hemangioma|9131/0
C0206733|T191|PT|MTHU040685|ICPC2ICD10ENG|juvenile; hemangioma|9131/0
C0206733|T191|PT|MTHU051505|ICPC2ICD10ENG|nevus; angiomatous|9131/0
C0206733|T191|PT|MTHU051507|ICPC2ICD10ENG|nevus; capillary|9131/0
C0206733|T191|PT|MTHU051503|ICPC2ICD10ENG|nevus; strawberry|9131/0
C0206733|T191|PT|MTHU060147|ICPC2ICD10ENG|plexiform; hemangioma|9131/0
C0085653|T191|PT|MTHU063427|ICPC2ICD10ENG|pyogenic; granuloma|9131/0
C0206733|T191|PT|MTHU067895|ICPC2ICD10ENG|simplex; hemangioma|9131/0
C0206733|T191|PT|MTHU001646|ICPC2ICD10ENG|strawberry; nevus|9131/0
C0085653|T191|PT|MTHU073641|ICPC2ICD10ENG|telangiectaticum; granuloma|9131/0
C0206733|T191|PT|S81004|ICPC2P|Mark;raspberry|9131/0
C0206733|T191|PT|S81005|ICPC2P|Mark;strawberry|9131/0
C0206733|T191|PTN|S81004|ICPC2P|raspberry mark|9131/0
C0206733|T191|PTN|S81005|ICPC2P|strawberry mark|9131/0
C0206733|T191|LLT|10007197|MDR|Capillary naevus|9131/0
C0206733|T191|LLT|10062789|MDR|Capillary nevus|9131/0
C0085653|T191|LLT|10078020|MDR|Granuloma telangiectaticum|9131/0
C0206733|T191|LLT|10055906|MDR|Haemangioma simplex|9131/0
C0206733|T191|LLT|10019404|MDR|Hemangioma simplex|9131/0
C0085653|T191|LLT|10037649|MDR|Pyogenic granuloma|9131/0
C0085653|T191|PT|10037649|MDR|Pyogenic granuloma|9131/0
C0206733|T191|LLT|10042171|MDR|Strawberry mark|9131/0
C0206733|T191|LLT|10042172|MDR|Strawberry naevus|9131/0
C0206733|T191|LLT|10062803|MDR|Strawberry nevus|9131/0
C0206733|T191|PT|10396|MEDCIN|capillary hemangioma|9131/0
C0206733|T191|SY|10396|MEDCIN|hemangioma capillary|9131/0
C0206733|T191|PT|261561|MEDCIN|strawberry nevus|9131/0
C0206733|T191|PT|272076|MEDCIN|strawberry nevus|9131/0
C0206733|T191|SY|261561|MEDCIN|strawberry nevus was observed|9131/0
C0206733|T191|SY|5402|MEDLINEPLUS|Strawberry mark|9131/0
C0206733|T191|PM|D018324|MSH|Capillary Hemangioma|9131/0
C0085653|T191|PM|D017789|MSH|Capillary Hemangioma, Lobular|9131/0
C0206733|T191|PM|D018324|MSH|Capillary Hemangiomas|9131/0
C0085653|T191|ET|D017789|MSH|Granuloma Pyogenicum|9131/0
C0085653|T191|ET|D017789|MSH|Granuloma Telangiecticum|9131/0
C0085653|T191|MH|D017789|MSH|Granuloma, Pyogenic|9131/0
C0206733|T191|MH|D018324|MSH|Hemangioma, Capillary|9131/0
C0085653|T191|ET|D017789|MSH|Hemangioma, Lobular Capillary|9131/0
C0206733|T191|PM|D018324|MSH|Hemangiomas, Capillary|9131/0
C0085653|T191|PM|D017789|MSH|Lobular Capillary Hemangioma|9131/0
C0085653|T191|PM|D017789|MSH|Pyogenic Granuloma|9131/0
C0085653|T191|PN|NOCODE|MTH|Pyogenic granuloma|9131/0
C0206733|T191|PN|NOCODE|MTH|Strawberry nevus of skin|9131/0
C0085653|T191|ET|686.1|MTHICD9|Granuloma, suppurative|9131/0
C0085653|T191|ET|686.1|MTHICD9|Granuloma, telangiectaticum|9131/0
C0206733|T191|ET|757.32|MTHICD9|Strawberry nevus|9131/0
C0206733|T191|SY|C7457|NCI|Capillary Angioma|9131/0
C0206733|T191|PT|C7457|NCI|Capillary Hemangioma|9131/0
C0085653|T191|SY|C3480|NCI|Granulation Tissue-Type Hemangioma|9131/0
C0085653|T191|SY|C3480|NCI|Granuloma Pyogenicum|9131/0
C0085653|T191|SY|C3480|NCI|Granuloma Telangiecticum|9131/0
C0085653|T191|SY|C3480|NCI|Granulomata Pyogenicum|9131/0
C0085653|T191|SY|C3480|NCI|Hemangiomatous Granulation Tissue|9131/0
C0085653|T191|PT|C3480|NCI|Lobular Hemangioma|9131/0
C0085653|T191|SY|C3480|NCI|Pyogenic Granuloma|9131/0
C0085653|T191|SY|C3480|NCI_NICHD|Lobular Capillary Hemangioma|9131/0
C0085653|T191|PT|C3480|NCI_NICHD|Pyogenic Granuloma|9131/0
C0085653|T191|PT|CDR0000779854|PDQ|adult lobular hemangioma|9131/0
C0085653|T191|SY|CDR0000779854|PDQ|granulation tissue-type hemangioma|9131/0
C0085653|T191|SY|CDR0000779854|PDQ|granuloma pyogenicum|9131/0
C0085653|T191|SY|CDR0000779854|PDQ|granuloma telangiecticum|9131/0
C0085653|T191|SY|CDR0000779854|PDQ|granulomata pyogenicum|9131/0
C0085653|T191|SY|CDR0000779854|PDQ|hemangiomatous granulation tissue|9131/0
C0085653|T191|SY|CDR0000779854|PDQ|lobular hemangioma|9131/0
C0085653|T191|SY|CDR0000779854|PDQ|pyogenic granuloma|9131/0
C0206733|T191|SY|X78DE|RCD|Angiomatous naevus|9131/0
C0206733|T191|SY|G7710|RCD|Capillary angioma|9131/0
C0206733|T191|PT|BBT8.|RCD|Capillary haemangioma|9131/0
C0206733|T191|SY|PH312|RCD|Capillary haemangioma of skin|9131/0
C0206733|T191|SY|BBT8.|RCD|Capillary naevus|9131/0
C0206733|T191|SY|PH312|RCD|Capillary naevus of skin|9131/0
C0206733|T191|PT|X78DE|RCD|Congenital vascular naevus|9131/0
C0206733|T191|SY|BBT8.|RCD|Haemangioma simplex|9131/0
C0206733|T191|SY|BBT8.|RCD|Infantile haemangioma|9131/0
C0206733|T191|SY|BBT8.|RCD|Juvenile haemangioma|9131/0
C0206733|T191|SY|BBT8.|RCD|Plexiform haemangioma|9131/0
C0085653|T191|OP|M071z|RCD|Pyogenic granuloma NOS|9131/0
C0085653|T191|OP|M0710|RCD|Pyogenic granuloma unspecified|9131/0
C0206733|T191|SY|PH312|RCD|Strawberry angioma|9131/0
C0206733|T191|SY|PH312|RCD|Strawberry birthmark|9131/0
C0206733|T191|SY|PH312|RCD|Strawberry mark|9131/0
C0206733|T191|SY|PH312|RCD|Strawberry naevus|9131/0
C0206733|T191|SY|X78DE|RCDAE|Angiomatous nevus|9131/0
C0206733|T191|PT|BBT8.|RCDAE|Capillary hemangioma|9131/0
C0206733|T191|SY|PH312|RCDAE|Capillary hemangioma of skin|9131/0
C0206733|T191|SY|BBT8.|RCDAE|Capillary nevus|9131/0
C0206733|T191|SY|PH312|RCDAE|Capillary nevus of skin|9131/0
C0206733|T191|PT|X78DE|RCDAE|Congenital vascular nevus|9131/0
C0206733|T191|SY|BBT8.|RCDAE|Hemangioma simplex|9131/0
C0206733|T191|SY|BBT8.|RCDAE|Infantile hemangioma|9131/0
C0206733|T191|SY|BBT8.|RCDAE|Juvenile hemangioma|9131/0
C0206733|T191|SY|BBT8.|RCDAE|Plexiform hemangioma|9131/0
C0206733|T191|SY|PH312|RCDAE|Strawberry nevus|9131/0
C0206733|T191|SYGB|83343001|SNOMEDCT_US|Angiomatous naevus|9131/0
C0206733|T191|SYGB|254206003|SNOMEDCT_US|Angiomatous naevus|9131/0
C0206733|T191|SYGB|56975005|SNOMEDCT_US|Angiomatous naevus of skin|9131/0
C0206733|T191|SY|83343001|SNOMEDCT_US|Angiomatous nevus|9131/0
C0206733|T191|SY|254206003|SNOMEDCT_US|Angiomatous nevus|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Angiomatous nevus of skin|9131/0
C0206733|T191|SY|195382003|SNOMEDCT_US|Capillary angioma|9131/0
C0206733|T191|PTGB|83343001|SNOMEDCT_US|Capillary haemangioma|9131/0
C0206733|T191|PTGB|402867006|SNOMEDCT_US|Capillary haemangioma|9131/0
C0085653|T191|SYGB|17372009|SNOMEDCT_US|Capillary haemangioma of granulation tissue type|9131/0
C0206733|T191|SYGB|56975005|SNOMEDCT_US|Capillary haemangioma of skin|9131/0
C0206733|T191|PT|83343001|SNOMEDCT_US|Capillary hemangioma|9131/0
C0206733|T191|PT|402867006|SNOMEDCT_US|Capillary hemangioma|9131/0
C0085653|T191|SY|17372009|SNOMEDCT_US|Capillary hemangioma of granulation tissue type|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Capillary hemangioma of skin|9131/0
C0206733|T191|SYGB|83343001|SNOMEDCT_US|Capillary naevus|9131/0
C0206733|T191|SYGB|56975005|SNOMEDCT_US|Capillary naevus of skin|9131/0
C0206733|T191|SY|83343001|SNOMEDCT_US|Capillary nevus|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Capillary nevus of skin|9131/0
C0206733|T191|SY|254206003|SNOMEDCT_US|Congenital vascular hamartoma|9131/0
C0206733|T191|OAS|205560007|SNOMEDCT_US|Congenital vascular naevus|9131/0
C0206733|T191|PTGB|254206003|SNOMEDCT_US|Congenital vascular naevus|9131/0
C0206733|T191|PT|254206003|SNOMEDCT_US|Congenital vascular nevus|9131/0
C0206733|T191|OAS|205560007|SNOMEDCT_US|Congenital vascular nevus|9131/0
C0085653|T191|PT|17372009|SNOMEDCT_US|Granuloma pyogenicum|9131/0
C0085653|T191|SY|17372009|SNOMEDCT_US|Granuloma telangiectaticum|9131/0
C0085653|T191|IS|17372009|SNOMEDCT_US|Granulomatous polyp|9131/0
C0206733|T191|SYGB|83343001|SNOMEDCT_US|Haemangioma simplex|9131/0
C0206733|T191|SY|83343001|SNOMEDCT_US|Hemangioma simplex|9131/0
C0206733|T191|SYGB|83343001|SNOMEDCT_US|Infantile haemangioma|9131/0
C0206733|T191|SY|83343001|SNOMEDCT_US|Infantile hemangioma|9131/0
C0206733|T191|SYGB|83343001|SNOMEDCT_US|Juvenile haemangioma|9131/0
C0206733|T191|SY|83343001|SNOMEDCT_US|Juvenile hemangioma|9131/0
C0085653|T191|SYGB|17372009|SNOMEDCT_US|Lobular capillary haemangioma|9131/0
C0085653|T191|SY|17372009|SNOMEDCT_US|Lobular capillary hemangioma|9131/0
C0085653|T191|SY|39629007|SNOMEDCT_US|PG - Pyogenic granuloma|9131/0
C0206733|T191|SYGB|83343001|SNOMEDCT_US|Plexiform haemangioma|9131/0
C0206733|T191|SY|83343001|SNOMEDCT_US|Plexiform hemangioma|9131/0
C0206733|T191|SY|83343001|SNOMEDCT_US|Port wine stain|9131/0
C0085653|T191|OAS|267838007|SNOMEDCT_US|Pyogenic granuloma|9131/0
C0085653|T191|OF|200722003|SNOMEDCT_US|Pyogenic granuloma|9131/0
C0085653|T191|OF|395604005|SNOMEDCT_US|Pyogenic granuloma|9131/0
C0085653|T191|OAP|395604005|SNOMEDCT_US|Pyogenic granuloma|9131/0
C0085653|T191|PT|200722003|SNOMEDCT_US|Pyogenic granuloma|9131/0
C0085653|T191|OAS|156323008|SNOMEDCT_US|Pyogenic granuloma|9131/0
C0085653|T191|SY|17372009|SNOMEDCT_US|Pyogenic granuloma|9131/0
C0085653|T191|OAP|200725001|SNOMEDCT_US|Pyogenic granuloma NOS|9131/0
C0085653|T191|OAP|200720006|SNOMEDCT_US|Pyogenic granuloma unspecified|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Raspberry mark of skin|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Strawberry angioma|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Strawberry birthmark|9131/0
C0206733|T191|SYGB|56975005|SNOMEDCT_US|Strawberry haemangioma of skin|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Strawberry hemangioma of skin|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Strawberry mark|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Strawberry mark of skin|9131/0
C0206733|T191|SYGB|56975005|SNOMEDCT_US|Strawberry naevus|9131/0
C0206733|T191|PTGB|56975005|SNOMEDCT_US|Strawberry naevus of skin|9131/0
C0206733|T191|SY|56975005|SNOMEDCT_US|Strawberry nevus|9131/0
C0206733|T191|PT|56975005|SNOMEDCT_US|Strawberry nevus of skin|9131/0
C0206733|T191|IS|56975005|SNOMEDCT_US|Strawberry nevus of skin, NOS|9131/0
C0085653|T191|PT|1680|WHO|PYOGENIC GRANULOMA|9131/0
C0206733|T191|IT|0764|WHO|STRAWBERRY MARK|9131/0
C0205789|T191|PT|0000020717|CHV|intramuscular haemangioma|9132/0
C0205789|T191|SY|0000020717|CHV|intramuscular hemangioma|9132/0
C0205789|T191|PT|MTHU033770|ICPC2ICD10ENG|hemangioma; intramuscular|9132/0
C0205789|T191|PT|MTHU040072|ICPC2ICD10ENG|intramuscular; hemangioma|9132/0
C0205789|T191|PEP|D006391|MSH|Hemangioma, Intramuscular|9132/0
C0205789|T191|PM|D006391|MSH|Hemangiomas, Intramuscular|9132/0
C0205789|T191|PM|D006391|MSH|Intramuscular Hemangioma|9132/0
C0205789|T191|PM|D006391|MSH|Intramuscular Hemangiomas|9132/0
C0205789|T191|SY|C3699|NCI|Intramuscular Angioma|9132/0
C0205789|T191|PT|C3699|NCI|Intramuscular Hemangioma|9132/0
C0205789|T191|PT|BBT9.|RCD|Intramuscular haemangioma|9132/0
C0205789|T191|PT|BBT9.|RCDAE|Intramuscular hemangioma|9132/0
C0205789|T191|SY|54249004|SNOMEDCT_US|Intramuscular angioma|9132/0
C0205789|T191|PTGB|54249004|SNOMEDCT_US|Intramuscular haemangioma|9132/0
C0205789|T191|PT|54249004|SNOMEDCT_US|Intramuscular hemangioma|9132/0
C0206732|T191|PT|0000021056|CHV|epithelioid hemangioendothelioma|9133/1
C0206732|T191|LLT|10079874|MDR|Epithelioid haemangioendothelioma|9133/1
C0206732|T191|LLT|10079873|MDR|Epithelioid hemangioendothelioma|9133/1
C0206732|T191|PT|355058|MEDCIN|epithelioid hemangioendothelioma|9133/1
C0206732|T191|SY|355058|MEDCIN|neoplasm - soft tissue blood vessel hemangioendothelioma epithelioid|9133/1
C0206732|T191|PM|D018323|MSH|Epithelioid Hemangioendothelioma|9133/1
C0206732|T191|PM|D018323|MSH|Epithelioid Hemangioendotheliomas|9133/1
C0206732|T191|MH|D018323|MSH|Hemangioendothelioma, Epithelioid|9133/1
C0206732|T191|PM|D018323|MSH|Hemangioendotheliomas, Epithelioid|9133/1
C0206732|T191|PN|NOCODE|MTH|Epithelioid hemangioendothelioma|9133/1
C0206732|T191|SY|C3800|NCI|Epithelioid Angioendothelioma|9133/1
C0206732|T191|SY|C3800|NCI|Epithelioid Angiosarcoma|9133/1
C0206732|T191|PT|C3800|NCI|Epithelioid Hemangioendothelioma|9133/1
C0206732|T191|AB|X77p4|RCD|Epithel haemangioendothelioma|9133/1
C0206732|T191|PT|X77p4|RCD|Epithelioid haemangioendothelioma|9133/1
C0206732|T191|AB|X77p4|RCDAE|Epithel hemangioendothelioma|9133/1
C0206732|T191|PT|X77p4|RCDAE|Epithelioid hemangioendothelioma|9133/1
C0206732|T191|OP|BBTJ.|RCDSA|Epithelioid hemangioendothelioma NOS|9133/1
C0206732|T191|OA|BBTJ.|RCDSY|Epithe haemngioendothelioma|9133/1
C0206732|T191|OP|BBTJ.|RCDSY|Epithelioid haemangioendothelioma NOS|9133/1
C0206732|T191|PTGB|403981003|SNOMEDCT_US|Epithelioid haemangioendothelioma|9133/1
C0206732|T191|OAP|84290008|SNOMEDCT_US|Epithelioid haemangioendothelioma|9133/1
C0206732|T191|PT|403981003|SNOMEDCT_US|Epithelioid hemangioendothelioma|9133/1
C0206732|T191|OAP|84290008|SNOMEDCT_US|Epithelioid hemangioendothelioma|9133/1
C0206732|T191|IS|84290008|SNOMEDCT_US|Epithelioid hemangioendothelioma, NOS|9133/1
C0206732|T191|PT|0000021056|CHV|epithelioid hemangioendothelioma|9133/3
C0206732|T191|LLT|10079874|MDR|Epithelioid haemangioendothelioma|9133/3
C0206732|T191|LLT|10079873|MDR|Epithelioid hemangioendothelioma|9133/3
C0206732|T191|PT|355058|MEDCIN|epithelioid hemangioendothelioma|9133/3
C0334538|T191|PT|271556|MEDCIN|malignant epithelioid hemangioendothelioma|9133/3
C0206732|T191|SY|355058|MEDCIN|neoplasm - soft tissue blood vessel hemangioendothelioma epithelioid|9133/3
C0206732|T191|PM|D018323|MSH|Epithelioid Hemangioendothelioma|9133/3
C0206732|T191|PM|D018323|MSH|Epithelioid Hemangioendotheliomas|9133/3
C0206732|T191|MH|D018323|MSH|Hemangioendothelioma, Epithelioid|9133/3
C0206732|T191|PM|D018323|MSH|Hemangioendotheliomas, Epithelioid|9133/3
C0206732|T191|PN|NOCODE|MTH|Epithelioid hemangioendothelioma|9133/3
C0334538|T191|PN|NOCODE|MTH|Epithelioid hemangioendothelioma, malignant|9133/3
C0206732|T191|SY|C3800|NCI|Epithelioid Angioendothelioma|9133/3
C0206732|T191|SY|C3800|NCI|Epithelioid Angiosarcoma|9133/3
C0206732|T191|PT|C3800|NCI|Epithelioid Hemangioendothelioma|9133/3
C0206732|T191|AB|X77p4|RCD|Epithel haemangioendothelioma|9133/3
C0206732|T191|PT|X77p4|RCD|Epithelioid haemangioendothelioma|9133/3
C0334538|T191|AB|X77p3|RCD|Mal epith haemangioendotheliom|9133/3
C0334538|T191|PT|X77p3|RCD|Malignant epithelioid haemangioendothelioma|9133/3
C0206732|T191|AB|X77p4|RCDAE|Epithel hemangioendothelioma|9133/3
C0206732|T191|PT|X77p4|RCDAE|Epithelioid hemangioendothelioma|9133/3
C0334538|T191|PT|X77p3|RCDAE|Malignant epithelioid hemangioendothelioma|9133/3
C0206732|T191|OP|BBTJ.|RCDSA|Epithelioid hemangioendothelioma NOS|9133/3
C0334538|T191|SY|X77p3|RCDSA|Epithelioid hemangioendothelioma, malignant|9133/3
C0206732|T191|OA|BBTJ.|RCDSY|Epithe haemngioendothelioma|9133/3
C0206732|T191|OP|BBTJ.|RCDSY|Epithelioid haemangioendothelioma NOS|9133/3
C0334538|T191|SY|X77p3|RCDSY|Epithelioid haemangioendothelioma, malignant|9133/3
C0334538|T191|AB|X77p3|RCDSY|Epithld haemngendthel, malg|9133/3
C0334538|T191|PTGB|54124005|SNOMEDCT_US|Epithelioid haemangioendothelioma|9133/3
C0206732|T191|OAP|84290008|SNOMEDCT_US|Epithelioid haemangioendothelioma|9133/3
C0206732|T191|PTGB|403981003|SNOMEDCT_US|Epithelioid haemangioendothelioma|9133/3
C0334538|T191|SYGB|54124005|SNOMEDCT_US|Epithelioid haemangioendothelioma, malignant|9133/3
C0334538|T191|PT|54124005|SNOMEDCT_US|Epithelioid hemangioendothelioma|9133/3
C0206732|T191|PT|403981003|SNOMEDCT_US|Epithelioid hemangioendothelioma|9133/3
C0206732|T191|OAP|84290008|SNOMEDCT_US|Epithelioid hemangioendothelioma|9133/3
C0334538|T191|SY|54124005|SNOMEDCT_US|Epithelioid hemangioendothelioma, malignant|9133/3
C0206732|T191|IS|84290008|SNOMEDCT_US|Epithelioid hemangioendothelioma, NOS|9133/3
C0334538|T191|OAP|189872002|SNOMEDCT_US|Malignant epithelioid haemangioendothelioma|9133/3
C0334538|T191|OF|189872002|SNOMEDCT_US|Malignant epithelioid haemangioendothelioma|9133/3
C0334538|T191|OAP|189872002|SNOMEDCT_US|Malignant epithelioid hemangioendothelioma|9133/3
C0346087|T191|PT|0000031044|CHV|dabska tumor|9135/1
C0346087|T191|PN|NOCODE|MTH|Endovascular papillary angioendothelioma|9135/1
C0346087|T191|SY|C7526|NCI|Dabska Tumor|9135/1
C0346087|T191|SY|C7526|NCI|Malignant Endothelial Papillary Angioendothelioma|9135/1
C0346087|T191|SY|C7526|NCI|Papillary Endovascular Angioendothelioma|9135/1
C0346087|T191|PT|C7526|NCI|Papillary Intralymphatic Angioendothelioma|9135/1
C0346087|T191|AB|C7526|NCI|PILA|9135/1
C0346087|T191|SY|128768006|SNOMEDCT_US|Dabska tumor|9135/1
C0346087|T191|SYGB|128768006|SNOMEDCT_US|Dabska tumour|9135/1
C0346087|T191|PT|128768006|SNOMEDCT_US|Endovascular papillary angioendothelioma|9135/1
C0346087|T191|SY|128768006|SNOMEDCT_US|Papillary intralymphatic angioendomethelioma|9135/1
C1304508|T191|PN|NOCODE|MTH|Spindle cell hemangioma|9136/0
C1304508|T191|AB|C4754|NCI|SCH|9136/0
C1304508|T191|SY|C4754|NCI|Spindle -Cell Hemangioma|9136/0
C1304508|T191|SY|C4754|NCI|Spindle Cell Hemangioendothelioma|9136/0
C1304508|T191|PT|C4754|NCI|Spindle Cell Hemangioma|9136/0
C1304508|T191|PT|CDR0000779851|PDQ|adult spindle cell hemangioma|9136/0
C1304508|T191|AB|CDR0000779851|PDQ|SCH|9136/0
C1304508|T191|SY|CDR0000779851|PDQ|spindle cell hemangioendothelioma|9136/0
C1304508|T191|SY|CDR0000779851|PDQ|Spindle Cell Hemangioma|9136/0
C1304508|T191|SY|CDR0000779851|PDQ|spindle-cell hemangioma|9136/0
C1304508|T191|AB|Xa0Za|RCD|Spindle cell haemangendothelom|9136/0
C1304508|T191|PT|Xa0Za|RCD|Spindle cell haemangioendothelioma|9136/0
C1304508|T191|PT|Xa0Za|RCDAE|Spindle cell hemangioendothelioma|9136/0
C1304508|T191|SY|128769003|SNOMEDCT_US|Spindle cell angioendothelioma|9136/0
C1304508|T191|OAP|134304005|SNOMEDCT_US|Spindle cell haemangioendothelioma|9136/0
C1304508|T191|PTGB|128769003|SNOMEDCT_US|Spindle cell haemangioendothelioma|9136/0
C1304508|T191|PTGB|403967000|SNOMEDCT_US|Spindle cell haemangioma|9136/0
C1304508|T191|SYGB|128769003|SNOMEDCT_US|Spindle cell haemangioma|9136/0
C1304508|T191|PT|128769003|SNOMEDCT_US|Spindle cell hemangioendothelioma|9136/0
C1304508|T191|OAP|134304005|SNOMEDCT_US|Spindle cell hemangioendothelioma|9136/0
C1304508|T191|PT|403967000|SNOMEDCT_US|Spindle cell hemangioma|9136/0
C1304508|T191|SY|128769003|SNOMEDCT_US|Spindle cell hemangioma|9136/0
C1304513|T191|PT|355053|MEDCIN|Composite hemangioendothelioma|9136/1
C1304513|T191|SY|355053|MEDCIN|neoplasm - soft tissue blood vessel hemangioendothelioma composite|9136/1
C1304512|T191|SY|355051|MEDCIN|neoplasm - soft tissue blood vessel hemangioendothelioma retiform|9136/1
C1304512|T191|PT|355051|MEDCIN|Retiform hemangioendothelioma|9136/1
C1304508|T191|PN|NOCODE|MTH|Spindle cell hemangioma|9136/1
C1304513|T191|PT|C45475|NCI|Composite Hemangioendothelioma|9136/1
C3840252|T191|SY|C121668|NCI|Epithelioid Sarcoma-Like Hemangioendothelioma|9136/1
C1304512|T191|SY|C27511|NCI|Hobnail Hemangioendothelioma|9136/1
C3840252|T191|PT|C121668|NCI|Pseudomyogenic Hemangioendothelioma|9136/1
C1304512|T191|PT|C27511|NCI|Retiform Hemangioendothelioma|9136/1
C1304508|T191|AB|C4754|NCI|SCH|9136/1
C1304508|T191|SY|C4754|NCI|Spindle -Cell Hemangioma|9136/1
C1304508|T191|SY|C4754|NCI|Spindle Cell Hemangioendothelioma|9136/1
C1304508|T191|PT|C4754|NCI|Spindle Cell Hemangioma|9136/1
C1304513|T191|PT|CDR0000779859|PDQ|adult composite hemangioendothelioma|9136/1
C1304512|T191|PT|CDR0000779857|PDQ|adult retiform hemangioendothelioma|9136/1
C1304508|T191|PT|CDR0000779851|PDQ|adult spindle cell hemangioma|9136/1
C1304513|T191|SY|CDR0000779859|PDQ|composite hemangioendothelioma|9136/1
C1304512|T191|SY|CDR0000779857|PDQ|hobnail hemangioendothelioma|9136/1
C1304512|T191|SY|CDR0000779857|PDQ|retiform hemangioendothelioma|9136/1
C1304508|T191|AB|CDR0000779851|PDQ|SCH|9136/1
C1304508|T191|SY|CDR0000779851|PDQ|spindle cell hemangioendothelioma|9136/1
C1304508|T191|SY|CDR0000779851|PDQ|Spindle Cell Hemangioma|9136/1
C1304508|T191|SY|CDR0000779851|PDQ|spindle-cell hemangioma|9136/1
C1304508|T191|AB|Xa0Za|RCD|Spindle cell haemangendothelom|9136/1
C1304508|T191|PT|Xa0Za|RCD|Spindle cell haemangioendothelioma|9136/1
C1304508|T191|PT|Xa0Za|RCDAE|Spindle cell hemangioendothelioma|9136/1
C1304513|T191|PTGB|703660008|SNOMEDCT_US|Composite haemangioendothelioma|9136/1
C1304513|T191|PTGB|403984006|SNOMEDCT_US|Composite haemangioendothelioma|9136/1
C1304513|T191|PT|703660008|SNOMEDCT_US|Composite hemangioendothelioma|9136/1
C1304513|T191|PT|403984006|SNOMEDCT_US|Composite hemangioendothelioma|9136/1
C1304512|T191|PTGB|703659003|SNOMEDCT_US|Retiform haemangioendothelioma|9136/1
C1304512|T191|PTGB|403982005|SNOMEDCT_US|Retiform haemangioendothelioma|9136/1
C1304512|T191|PT|703659003|SNOMEDCT_US|Retiform hemangioendothelioma|9136/1
C1304512|T191|PT|403982005|SNOMEDCT_US|Retiform hemangioendothelioma|9136/1
C1304508|T191|SY|128769003|SNOMEDCT_US|Spindle cell angioendothelioma|9136/1
C1304508|T191|OAP|134304005|SNOMEDCT_US|Spindle cell haemangioendothelioma|9136/1
C1304508|T191|PTGB|128769003|SNOMEDCT_US|Spindle cell haemangioendothelioma|9136/1
C1304508|T191|PTGB|403967000|SNOMEDCT_US|Spindle cell haemangioma|9136/1
C1304508|T191|SYGB|128769003|SNOMEDCT_US|Spindle cell haemangioma|9136/1
C1304508|T191|OAP|134304005|SNOMEDCT_US|Spindle cell hemangioendothelioma|9136/1
C1304508|T191|PT|128769003|SNOMEDCT_US|Spindle cell hemangioendothelioma|9136/1
C1304508|T191|SY|128769003|SNOMEDCT_US|Spindle cell hemangioma|9136/1
C1304508|T191|PT|403967000|SNOMEDCT_US|Spindle cell hemangioma|9136/1
C1708550|T191|PT|C53677|NCI|Intimal Sarcoma|9137/3
C1708550|T191|PT|703661007|SNOMEDCT_US|Intimal sarcoma|9137/3
C0036220|T191|ET|0000004562|AOD|Kaposi sarcoma|9140/3
C0036220|T191|PT|BI00726|BI|kaposi's sarcoma|9140/3
C0036220|T191|AB|BI00726|BI|ks|9140/3
C0036220|T191|PT|0043734|CCPSS|KAPOSI SARCOMA|9140/3
C0036220|T191|PT|0000011049|CHV|kaposi sarcoma|9140/3
C0036220|T191|PT|NOCODE|COSTAR|Kaposi's Sarcoma|9140/3
C0036220|T191|PT|U000396|COSTAR|KAPOSIS SARCOMA|9140/3
C0036220|T191|ET|2007-1936|CSP|HHV 8|9140/3
C0036220|T191|ET|2007-1936|CSP|HHV8|9140/3
C0036220|T191|PT|2007-1936|CSP|Kaposi's sarcoma|9140/3
C0036220|T191|SY|NOCODE|DXP|ENDOTHELIOSARCOMA|9140/3
C0036220|T191|SY|NOCODE|DXP|KAPOSI CANCER, SARCOMA|9140/3
C0036220|T191|DI|U000963|DXP|KAPOSI SARCOMA|9140/3
C0036220|T191|FI|U002235|DXP|KAPOSI SARCOMA|9140/3
C0036220|T191|SY|NOCODE|DXP|SARCOMA, MULTIPLE IDIOPATHIC HEMORRHAGIC|9140/3
C0036220|T191|PT|HP:0100726|HPO|Kaposi's sarcoma|9140/3
C0036220|T191|HT|C46|ICD10|Kaposi's sarcoma|9140/3
C0036220|T191|PT|C46.9|ICD10|Kaposi's sarcoma, unspecified|9140/3
C0036220|T191|HT|C46|ICD10CM|Kaposi's sarcoma|9140/3
C0036220|T191|AB|C46|ICD10CM|Kaposi's sarcoma|9140/3
C0036220|T191|ET|C46.9|ICD10CM|Kaposi's sarcoma of unspecified site|9140/3
C0036220|T191|PT|C46.9|ICD10CM|Kaposi's sarcoma, unspecified|9140/3
C0036220|T191|AB|C46.9|ICD10CM|Kaposi's sarcoma, unspecified|9140/3
C0036220|T191|HT|176|ICD9CM|Kaposi's sarcoma|9140/3
C0036220|T191|AB|176.9|ICD9CM|Kaposi's sarcoma NOS|9140/3
C0036220|T191|PT|176.9|ICD9CM|Kaposi's sarcoma, unspecified site|9140/3
C0036220|T191|PT|MTHU040818|ICPC2ICD10ENG|Kaposi; sarcoma|9140/3
C0036220|T191|PT|MTHU040828|ICPC2ICD10ENG|Kaposi; sarcoma, unspecified site|9140/3
C0036220|T191|PT|MTHU065905|ICPC2ICD10ENG|sarcoma; Kaposi|9140/3
C0036220|T191|PT|MTHU065915|ICPC2ICD10ENG|sarcoma; Kaposi, unspecified site|9140/3
C0036220|T191|PTN|A79010|ICPC2P|Kaposis sarcoma|9140/3
C0036220|T191|PT|A79010|ICPC2P|Sarcoma;Kaposis|9140/3
C0036220|T191|PT|sh85071562|LCH_NW|Kaposi's sarcoma|9140/3
C0036220|T191|LA|LA26517-5|LNC|Kaposi sarcoma|9140/3
C0036220|T191|LLT|10023284|MDR|Kaposi's sarcoma|9140/3
C0036220|T191|PT|10023284|MDR|Kaposi's sarcoma|9140/3
C0036220|T191|LLT|10023290|MDR|Kaposi's sarcoma NOS|9140/3
C0036220|T191|LLT|10023298|MDR|Kaposi's sarcoma, unspecified|9140/3
C0036220|T191|HT|10023285|MDR|Kaposi's sarcomas|9140/3
C0036220|T191|LLT|10028220|MDR|Multiple haemorrhagic sarcoma|9140/3
C0036220|T191|LLT|10028221|MDR|Multiple hemorrhagic sarcoma|9140/3
C0036220|T191|LLT|10055863|MDR|Multiple idiopathic haemorrhagic sarcoma|9140/3
C0036220|T191|LLT|10028222|MDR|Multiple idiopathic hemorrhagic sarcoma|9140/3
C0036220|T191|PT|99697|MEDCIN|Kaposi's sarcoma|9140/3
C0036220|T191|SY|99697|MEDCIN|malignant neoplasm sarcoma Kaposi's|9140/3
C0036220|T191|PT|481|MEDLINEPLUS|Kaposi Sarcoma|9140/3
C0036220|T191|SY|481|MEDLINEPLUS|KS|9140/3
C0036220|T191|ET|D012514|MSH|Kaposi Sarcoma|9140/3
C0036220|T191|ET|D012514|MSH|Kaposi's Sarcoma|9140/3
C0036220|T191|PM|D012514|MSH|Kaposis Sarcoma|9140/3
C0036220|T191|ET|D012514|MSH|Multiple Idiopathic Pigmented Hemangiosarcoma|9140/3
C0036220|T191|MH|D012514|MSH|Sarcoma, Kaposi|9140/3
C0036220|T191|PM|D012514|MSH|Sarcoma, Kaposi's|9140/3
C0036220|T191|PN|NOCODE|MTH|Kaposi Sarcoma|9140/3
C0036220|T191|ET|176.9|MTHICD9|Kaposi's sarcoma, unspecified|9140/3
C0036220|T191|PT|C9087|NCI|Kaposi Sarcoma|9140/3
C0036220|T191|SY|C9087|NCI|Kaposi's Sarcoma|9140/3
C0036220|T191|AB|C9087|NCI|KS|9140/3
C0036220|T191|SY|C9087|NCI|Multiple Hemorrhagic Sarcoma|9140/3
C0036220|T191|PT|C9087|NCI_CPTAC|Kaposi Sarcoma|9140/3
C0036220|T191|DN|C9087|NCI_CTRP|Kaposi Sarcoma|9140/3
C0036220|T191|PT|C9087|NCI_CTRP|Kaposi Sarcoma|9140/3
C0036220|T191|PT|CDR0000045134|NCI_NCI-GLOSS|Kaposi's sarcoma|9140/3
C0036220|T191|PSC|CDR0000038811|PDQ|Kaposi sarcoma|9140/3
C0036220|T191|SY|CDR0000038811|PDQ|multiple hemorrhagic sarcoma|9140/3
C0036220|T191|SY|CDR0000038811|PDQ|sarcoma, Kaposi's|9140/3
C0036220|T191|SY|CDR0000038811|PDQ|sarcoma, multiple hemorrhagic|9140/3
C0036220|T191|ET|CDR0000038811|PDQ|Skin cancer, Kaposi sarcoma|9140/3
C0036220|T191|PT|XaBBF|RCD|Kaposi's sarcoma|9140/3
C0036220|T191|SY|XaBBF|RCD|KS - Kaposi's sarcoma|9140/3
C0036220|T191|SY|XaBBF|RCD|Multiple haemorrhagic sarcoma|9140/3
C0036220|T191|SY|XaBBF|RCDAE|Multiple hemorrhagic sarcoma|9140/3
C0036220|T191|PT|BBTA.|RCDSY|Kaposi's sarcoma|9140/3
C0036220|T191|OP|Byu53|RCDSY|Kaposi's sarcoma, unspecified|9140/3
C0036220|T191|OA|Byu53|RCDSY|Kaposi's sarcoma,unspecifd|9140/3
C0036220|T191|SY|109385007|SNOMEDCT_US|Kaposi sarcoma|9140/3
C0036220|T191|SY|49937004|SNOMEDCT_US|Kaposi sarcoma, morphology|9140/3
C0036220|T191|SY|109385007|SNOMEDCT_US|Kaposi's sarcoma|9140/3
C0036220|T191|OAP|154604006|SNOMEDCT_US|Kaposi's sarcoma|9140/3
C0036220|T191|OF|154604006|SNOMEDCT_US|Kaposi's sarcoma|9140/3
C0036220|T191|PT|49937004|SNOMEDCT_US|Kaposi's sarcoma|9140/3
C0036220|T191|SY|49937004|SNOMEDCT_US|Kaposi's sarcoma, morphology|9140/3
C0036220|T191|SY|109385007|SNOMEDCT_US|KS - Kaposi's sarcoma|9140/3
C0036220|T191|SYGB|49937004|SNOMEDCT_US|Multiple haemorrhagic sarcoma|9140/3
C0036220|T191|SY|49937004|SNOMEDCT_US|Multiple hemorrhagic sarcoma|9140/3
C1299260|T191|PT|C156475|NCI|Metastatic Kaposi Sarcoma|9140/6
C1299260|T191|SY|372149006|SNOMEDCT_US|Kaposi sarcoma, metastatic|9140/6
C1299260|T191|PT|372149006|SNOMEDCT_US|Kaposi's sarcoma, metastatic|9140/6
C0002985|T191|PT|0000001172|CHV|angiokeratoma|9141/0
C0002985|T191|SY|0000001172|CHV|angiokeratomas|9141/0
C0002985|T191|ET|2007-0683|CSP|angiokeratoma|9141/0
C0002985|T191|PT|HP:0001014|HPO|Angiokeratoma|9141/0
C0002985|T191|SY|HP:0001014|HPO|Angiokeratomas|9141/0
C0002985|T191|LLT|10061639|MDR|Angiokeratoma|9141/0
C0002985|T191|PT|10061639|MDR|Angiokeratoma|9141/0
C0002985|T191|LLT|10052166|MDR|Angiokeratoma NOS|9141/0
C0002985|T191|MH|D000794|MSH|Angiokeratoma|9141/0
C0002985|T191|PM|D000794|MSH|Angiokeratomas|9141/0
C0002985|T191|PT|C2874|NCI|Angiokeratoma|9141/0
C0002985|T191|PT|BBTB.|RCD|Angiokeratoma|9141/0
C0002985|T191|PT|26810009|SNOMEDCT_US|Angiokeratoma|9141/0
C0334540|T191|PT|MTHU033777|ICPC2ICD10ENG|hemangioma; verrucous keratotic|9142/0
C0334540|T191|PT|MTHU080320|ICPC2ICD10ENG|verrucous; hemangioma, keratotic|9142/0
C0334540|T191|PT|MTHU080321|ICPC2ICD10ENG|verrucous; keratotic hemangioma|9142/0
C0334540|T191|SY|10398|MEDCIN|hemangioma verrucous|9142/0
C0334540|T191|PT|10398|MEDCIN|verrucous hemangioma|9142/0
C0334540|T191|PT|C4299|NCI|Verrucous Hemangioma|9142/0
C0334540|T191|SY|C4299|NCI|Verrucous Keratotic Hemangioma|9142/0
C0334540|T191|AB|BBTC.|RCD|Verrucous keratot haemangioma|9142/0
C0334540|T191|PT|BBTC.|RCD|Verrucous keratotic haemangioma|9142/0
C0334540|T191|AB|BBTC.|RCDAE|Verrucous keratot hemangioma|9142/0
C0334540|T191|PT|BBTC.|RCDAE|Verrucous keratotic hemangioma|9142/0
C0334540|T191|PTGB|20985003|SNOMEDCT_US|Verrucous keratotic haemangioma|9142/0
C0334540|T191|PT|20985003|SNOMEDCT_US|Verrucous keratotic hemangioma|9142/0
C0334541|T191|PT|0000030003|CHV|benign hemangiopericytoma|9150/0
C0334541|T191|SY|0000030003|CHV|hemangiopericytoma benign|9150/0
C0334541|T191|OP|C4300|NCI|Benign Hemangiopericytoma|9150/0
C0334541|T191|PT|C4300|NCI|Benign Hemangiopericytoma|9150/0
C0334541|T191|PT|C4300|NCI_CDISC|HEMANGIOPERICYTOMA, BENIGN|9150/0
C0334541|T191|PT|BBTD0|RCD|Benign haemangiopericytoma|9150/0
C0334541|T191|PT|BBTD0|RCDAE|Benign hemangiopericytoma|9150/0
C0334541|T191|SYGB|53880006|SNOMEDCT_US|Benign haemangiopericytoma|9150/0
C0334541|T191|SY|53880006|SNOMEDCT_US|Benign hemangiopericytoma|9150/0
C0334541|T191|PTGB|53880006|SNOMEDCT_US|Haemangiopericytoma, benign|9150/0
C0334541|T191|PT|53880006|SNOMEDCT_US|Hemangiopericytoma, benign|9150/0
C0018922|T191|SY|0000005939|CHV|haemangiopericytoma|9150/1
C0018922|T191|PT|0000005939|CHV|hemangiopericytoma|9150/1
C0018922|T191|SY|0000005939|CHV|perithelioma|9150/1
C0018922|T191|ET|2007-1041|CSP|hemangiopericytoma|9150/1
C4761161|T191|LLT|10082347|MDR|Glomangiopericytoma|9150/1
C4761161|T191|PT|10082347|MDR|Glomangiopericytoma|9150/1
C0018922|T191|PT|10018825|MDR|Haemangiopericytoma|9150/1
C0018922|T191|LLT|10018825|MDR|Haemangiopericytoma|9150/1
C0018922|T191|LLT|10060541|MDR|Hemangiopericytoma|9150/1
C0018922|T191|MTH_PT|10018825|MDR|Hemangiopericytoma|9150/1
C0018922|T191|PT|357931|MEDCIN|hemangiopericytoma|9150/1
C0018922|T191|SY|357931|MEDCIN|neoplasm - soft tissue uncertain behavior blood vessel hemangiopericytoma|9150/1
C0018922|T191|MH|D006393|MSH|Hemangiopericytoma|9150/1
C0018922|T191|PM|D006393|MSH|Hemangiopericytomas|9150/1
C0018922|T191|PN|NOCODE|MTH|hemangiopericytoma|9150/1
C0018922|T191|PT|C3087|NCI|Hemangiopericytoma|9150/1
C0018922|T191|OP|C3087|NCI|Hemangiopericytoma|9150/1
C0018922|T191|PT|CDR0000045707|NCI_NCI-GLOSS|hemangiopericytoma|9150/1
C0018922|T191|PT|Xa9AR|RCD|Haemangiopericytoma|9150/1
C0018922|T191|SY|Xa9AR|RCD|HPA - Haemangiopericytoma|9150/1
C0018922|T191|PT|Xa9AR|RCDAE|Hemangiopericytoma|9150/1
C0018922|T191|SY|Xa9AR|RCDAE|HPA - Hemangiopericytoma|9150/1
C0018922|T191|OP|BBTD1|RCDSA|Hemangiopericytoma NOS|9150/1
C0018922|T191|OP|BBTD1|RCDSY|Haemangiopericytoma NOS|9150/1
C4761161|T191|PT|822965001|SNOMEDCT_US|Glomangiopericytoma|9150/1
C0018922|T191|PTGB|36060005|SNOMEDCT_US|Haemangiopericytoma|9150/1
C0018922|T191|PTGB|134335004|SNOMEDCT_US|Haemangiopericytoma|9150/1
C0018922|T191|IS|36060005|SNOMEDCT_US|Haemangiopericytoma, NOS|9150/1
C0018922|T191|PT|36060005|SNOMEDCT_US|Hemangiopericytoma|9150/1
C0018922|T191|PT|134335004|SNOMEDCT_US|Hemangiopericytoma|9150/1
C0018922|T191|IS|36060005|SNOMEDCT_US|Hemangiopericytoma, NOS|9150/1
C0018922|T191|IS|134335004|SNOMEDCT_US|HPA - Haemangiopericytoma|9150/1
C0018922|T191|SYGB|134335004|SNOMEDCT_US|HPA - haemangiopericytoma|9150/1
C0018922|T191|IS|134335004|SNOMEDCT_US|HPA - Hemangiopericytoma|9150/1
C0018922|T191|SY|134335004|SNOMEDCT_US|HPA - hemangiopericytoma|9150/1
C0018922|T191|SY|36060005|SNOMEDCT_US|Perithelioma|9150/1
C0334542|T191|LLT|10025566|MDR|Malignant haemangiopericytoma|9150/3
C0334542|T191|PT|10025566|MDR|Malignant haemangiopericytoma|9150/3
C0334542|T191|LLT|10025569|MDR|Malignant haemangiopericytoma NOS|9150/3
C0334542|T191|LLT|10025571|MDR|Malignant haemangiopericytoma stage unspecified|9150/3
C0334542|T191|LLT|10060650|MDR|Malignant hemangiopericytoma|9150/3
C0334542|T191|MTH_PT|10025566|MDR|Malignant hemangiopericytoma|9150/3
C0334542|T191|MTH_LLT|10025569|MDR|Malignant hemangiopericytoma NOS|9150/3
C0334542|T191|LLT|10060654|MDR|Malignant hemangiopericytoma stage unspecified|9150/3
C0334542|T191|PT|271557|MEDCIN|malignant hemangiopericytoma|9150/3
C0334542|T191|NM|C562740|MSH|Hemangiopericytoma, Malignant|9150/3
C0334542|T191|PN|NOCODE|MTH|Hemangiopericytoma, Malignant|9150/3
C0334542|T191|OP|C4301|NCI|Malignant Hemangiopericytoma|9150/3
C0334542|T191|PT|C4301|NCI|Malignant Hemangiopericytoma|9150/3
C0334542|T191|OP|C4301|NCI|Malignant Hemangiopericytoma NOS|9150/3
C0334542|T191|PT|C4301|NCI_CDISC|HEMANGIOPERICYTOMA, MALIGNANT|9150/3
C0334542|T191|SY|C4301|NCI_CDISC|Malignant Hemangiopericytoma NOS|9150/3
C0334542|T191|PT|BBTD2|RCD|Malignant haemangiopericytoma|9150/3
C0334542|T191|PT|BBTD2|RCDAE|Malignant hemangiopericytoma|9150/3
C0334542|T191|PTGB|84664004|SNOMEDCT_US|Haemangiopericytoma, malignant|9150/3
C0334542|T191|PT|84664004|SNOMEDCT_US|Hemangiopericytoma, malignant|9150/3
C0334542|T191|SYGB|84664004|SNOMEDCT_US|Malignant haemangiopericytoma|9150/3
C0334542|T191|SY|84664004|SNOMEDCT_US|Malignant hemangiopericytoma|9150/3
C0206731|T191|PT|HP:0010615|HPO|Angiofibromas|9160/0
C0206731|T191|PT|MTHU028117|ICPC2ICD10ENG|fibrous; papule|9160/0
C0206731|T191|PT|MTHU057268|ICPC2ICD10ENG|papule; fibrous|9160/0
C0206731|T191|LLT|10002429|MDR|Angiofibroma|9160/0
C0206731|T191|PT|10002429|MDR|Angiofibroma|9160/0
C0206731|T191|LLT|10002430|MDR|Angiofibromatous hyperplasia|9160/0
C0206731|T191|MH|D018322|MSH|Angiofibroma|9160/0
C0206731|T191|PM|D018322|MSH|Angiofibromas|9160/0
C0206731|T191|PN|NOCODE|MTH|Angiofibroma|9160/0
C0206731|T191|PT|C3799|NCI|Angiofibroma|9160/0
C0206731|T191|SY|C3799|NCI|Angiofibromatous Hyperplasia|9160/0
C0206731|T191|SY|C3799|NCI|Fibrous Papule|9160/0
C0206731|T191|SY|C3799|NCI|Telangiectatic Fibroma|9160/0
C0206731|T191|PT|C3799|NCI_CDISC|ANGIOFIBROMA, BENIGN|9160/0
C0206731|T191|SY|C3799|NCI_CDISC|Angiofibromatous Hyperplasia|9160/0
C0206731|T191|SY|C3799|NCI_CDISC|Fibroangioma, Benign|9160/0
C0206731|T191|SY|C3799|NCI_CDISC|Fibrous Papule|9160/0
C0206731|T191|SY|C3799|NCI_CDISC|Telangiectatic Fibroma|9160/0
C0206731|T191|SY|CDR0000779848|PDQ|Angiofibroma|9160/0
C0206731|T191|SY|CDR0000779848|PDQ|angiofibromatous hyperplasia|9160/0
C0206731|T191|SY|CDR0000779848|PDQ|fibrous papule|9160/0
C0206731|T191|SY|CDR0000779848|PDQ|telangiectatic fibroma|9160/0
C0206731|T191|PT|Xa9AS|RCD|Angiofibroma|9160/0
C0206731|T191|OP|BBTE.|RCDSY|Angiofibroma NOS|9160/0
C0206731|T191|PT|302857002|SNOMEDCT_US|Angiofibroma|9160/0
C0206731|T191|PT|60392001|SNOMEDCT_US|Angiofibroma|9160/0
C0206731|T191|SY|60392001|SNOMEDCT_US|Angiofibroma, no ICD-O subtype|9160/0
C0206731|T191|SY|60392001|SNOMEDCT_US|Angiofibroma, no International Classification of Diseases for Oncology subtype|9160/0
C0206731|T191|IS|60392001|SNOMEDCT_US|Angiofibroma, NOS|9160/0
C0206731|T191|PT|1778|WHO|ANGIOFIBROMA|9160/0
C0206731|T191|IT|1778|WHO|ANGIOFIBROMATOUS HYPERPLASIA|9160/0
C0346073|T191|SY|HP:0012329|HPO|Angioblastoma|9161/0
C0346073|T191|SY|HP:0012329|HPO|Angioblastoma of Nakagawa|9161/0
C0346073|T191|SY|HP:0012329|HPO|Hypertrophic hemangioma|9161/0
C0346073|T191|SY|HP:0012329|HPO|Progressive capillary hemangioma|9161/0
C0346073|T191|PT|HP:0012329|HPO|Tufted angioma|9161/0
C0346073|T191|SY|HP:0012329|HPO|Tufted hemangioma|9161/0
C0346073|T191|CE|C536924|MSH|Angioma, tufted|9161/0
C0346073|T191|NM|C536924|MSH|Tufted angioma|9161/0
C0346073|T191|PN|NOCODE|MTH|Tufted angioma of skin|9161/0
C1266161|T191|PN|NOCODE|MTH|Tufted hemangioma|9161/0
C0346073|T191|SY|C4487|NCI|Angioblastoma of Nakagawa|9161/0
C0346073|T191|SY|C4487|NCI|Tufted Angioma|9161/0
C0346073|T191|SY|C4487|NCI|Tufted Angioma of Skin|9161/0
C0346073|T191|SY|C4487|NCI|Tufted Angioma of the Skin|9161/0
C0346073|T191|PT|C4487|NCI|Tufted Hemangioma|9161/0
C0346073|T191|SY|C4487|NCI|Tufted Hemangioma of Skin|9161/0
C0346073|T191|SY|C4487|NCI|Tufted Hemangioma of the Skin|9161/0
C0346073|T191|SY|C4487|NCI|Tufted Skin Angioma|9161/0
C0346073|T191|PT|CDR0000779850|PDQ|adult tufted hemangioma|9161/0
C0346073|T191|SY|CDR0000779850|PDQ|angioblastoma of Nakagawa|9161/0
C0346073|T191|SY|CDR0000779850|PDQ|tufted angioma|9161/0
C0346073|T191|SY|CDR0000779850|PDQ|tufted angioma of skin|9161/0
C0346073|T191|SY|CDR0000779850|PDQ|tufted angioma of the skin|9161/0
C0346073|T191|SY|CDR0000779850|PDQ|tufted hemangioma|9161/0
C0346073|T191|SY|CDR0000779850|PDQ|tufted hemangioma of skin|9161/0
C0346073|T191|SY|CDR0000779850|PDQ|tufted hemangioma of the skin|9161/0
C0346073|T191|SY|CDR0000779850|PDQ|tufted skin angioma|9161/0
C0346073|T191|PT|X78Uc|RCD|Tufted angioma of skin|9161/0
C1266161|T191|OP|128903007|SNOMEDCT_US|Acquired tufted haemangioma|9161/0
C1266161|T191|OP|128903007|SNOMEDCT_US|Acquired tufted hemangioma|9161/0
C0346073|T191|PT|705155008|SNOMEDCT_US|Tufted angioma|9161/0
C0346073|T191|PT|254786000|SNOMEDCT_US|Tufted angioma of skin|9161/0
C1266161|T191|PTGB|128903007|SNOMEDCT_US|Tufted haemangioma|9161/0
C1266161|T191|PT|128903007|SNOMEDCT_US|Tufted hemangioma|9161/0
C0206734|T191|ET|0000004548|AOD|hemangioblastoma|9161/1
C0206734|T191|PT|0053527|CCPSS|HEMANGIOBLASTOMA|9161/1
C0206734|T191|SY|0000021058|CHV|angioblastoma|9161/1
C0206734|T191|SY|0000021058|CHV|haemangioblastoma|9161/1
C0206734|T191|PT|0000021058|CHV|hemangioblastoma|9161/1
C0206734|T191|SY|0000021058|CHV|hemangioblastomas|9161/1
C0206734|T191|SY|HP:0010797|HPO|Haemangioblastoma|9161/1
C0206734|T191|PT|HP:0010797|HPO|Hemangioblastoma|9161/1
C0206734|T191|LLT|10018813|MDR|Haemangioblastoma|9161/1
C0206734|T191|PT|10018813|MDR|Haemangioblastoma|9161/1
C0206734|T191|LLT|10019385|MDR|Hemangioblastoma|9161/1
C0206734|T191|MTH_PT|10018813|MDR|Hemangioblastoma|9161/1
C0206734|T191|MH|D018325|MSH|Hemangioblastoma|9161/1
C0206734|T191|PM|D018325|MSH|Hemangioblastomas|9161/1
C0206734|T191|PN|NOCODE|MTH|Hemangioblastoma|9161/1
C0206734|T191|SY|C3801|NCI|Angioblastoma|9161/1
C0206734|T191|SY|C3801|NCI|Capillary Hemangioblastoma|9161/1
C0206734|T191|PT|C3801|NCI|Hemangioblastoma|9161/1
C0206734|T191|SY|TCGA|NCI|Hemangioblastoma|9161/1
C0206734|T191|SY|BBTF.|RCD|Angioblastoma|9161/1
C0206734|T191|PT|BBTF.|RCD|Haemangioblastoma|9161/1
C0206734|T191|PT|BBTF.|RCDAE|Hemangioblastoma|9161/1
C0206734|T191|SY|81201000|SNOMEDCT_US|Angioblastoma|9161/1
C0206734|T191|PTGB|81201000|SNOMEDCT_US|Haemangioblastoma|9161/1
C0206734|T191|PT|81201000|SNOMEDCT_US|Hemangioblastoma|9161/1
C0024221|T191|PT|1006008|CCPSS|LYMPHANGIOMA|9170/0
C0024221|T191|SY|0000007598|CHV|congenital lymphangioma|9170/0
C0024221|T191|PT|0000007598|CHV|lymphangioma|9170/0
C0024221|T191|SY|0000007598|CHV|lymphangiomas|9170/0
C0024221|T191|PT|NOCODE|COSTAR|Lymphangioma|9170/0
C0024221|T191|ET|2004-0139|CSP|lymphangioma|9170/0
C0024221|T191|PT|HP:0100764|HPO|Lymphangioma|9170/0
C0024221|T191|PT|D18.1|ICD10|Lymphangioma, any site|9170/0
C0024221|T191|AB|D18.1|ICD10CM|Lymphangioma, any site|9170/0
C0024221|T191|PT|D18.1|ICD10CM|Lymphangioma, any site|9170/0
C0024221|T191|PT|228.1|ICD9CM|Lymphangioma, any site|9170/0
C0024221|T191|AB|228.1|ICD9CM|Lymphangioma, any site|9170/0
C0024221|T191|PT|MTHU046582|ICPC2ICD10ENG|lymphangioma|9170/0
C0024221|T191|PTN|K72007|ICPC2P|lymphangioma|9170/0
C0024221|T191|OP|K99046|ICPC2P|Lymphangioma|9170/0
C0024221|T191|PT|K72007|ICPC2P|Lymphangioma|9170/0
C0024221|T191|OPN|K99046|ICPC2P|lymphangioma|9170/0
C0024221|T191|PT|10025219|MDR|Lymphangioma|9170/0
C0024221|T191|LLT|10025219|MDR|Lymphangioma|9170/0
C0024221|T191|LLT|10025220|MDR|Lymphangioma, any site|9170/0
C0024221|T191|PT|30773|MEDCIN|benign lymphangioma|9170/0
C0024221|T191|MH|D008202|MSH|Lymphangioma|9170/0
C0024221|T191|PM|D008202|MSH|Lymphangiomas|9170/0
C0024221|T191|ET|228.1|MTHICD9|Congenital lymphangioma|9170/0
C0024221|T191|PT|C8965|NCI|Lymphangioma|9170/0
C0024221|T191|PT|C8965|NCI_CDISC|LYMPHANGIOMA, BENIGN|9170/0
C0024221|T191|PT|C8965|NCI_NICHD|Lymphangioma|9170/0
C0024221|T191|PT|X77p7|RCD|Benign lymphangioma|9170/0
C0024221|T191|PT|X78WK|RCD|Congenital lymphangioma|9170/0
C0024221|T191|SY|X78WK|RCD|Lymphangioma|9170/0
C0024221|T191|PT|Xa9AT|RCD|Lymphangioma morphology|9170/0
C0024221|T191|OP|BBU0.|RCDSY|Lymphangioma NOS|9170/0
C0024221|T191|PT|253057002|SNOMEDCT_US|Benign lymphangioma|9170/0
C0024221|T191|OAP|189200000|SNOMEDCT_US|Congenital lymphangioma|9170/0
C0024221|T191|OF|189200000|SNOMEDCT_US|Congenital lymphangioma|9170/0
C0024221|T191|PT|254836000|SNOMEDCT_US|Congenital lymphangioma|9170/0
C0024221|T191|IS|254836000|SNOMEDCT_US|Lymphangioma|9170/0
C0024221|T191|OAS|154625006|SNOMEDCT_US|Lymphangioma|9170/0
C0024221|T191|PT|69044001|SNOMEDCT_US|Lymphangioma|9170/0
C0024221|T191|OAS|269646001|SNOMEDCT_US|Lymphangioma|9170/0
C0024221|T191|PT|400178008|SNOMEDCT_US|Lymphangioma|9170/0
C0024221|T191|SY|69044001|SNOMEDCT_US|Lymphangioma morphology|9170/0
C0024221|T191|OAP|93168006|SNOMEDCT_US|Lymphangioma of unspecified site|9170/0
C0024221|T191|SY|69044001|SNOMEDCT_US|Lymphangioma, no ICD-O subtype|9170/0
C0024221|T191|SY|69044001|SNOMEDCT_US|Lymphangioma, no International Classification of Diseases for Oncology subtype|9170/0
C0024221|T191|IS|69044001|SNOMEDCT_US|Lymphangioma, NOS|9170/0
C0024221|T191|SY|69044001|SNOMEDCT_US|Lymphangioma, site unspecified|9170/0
C0024221|T191|PT|1495|WHO|LYMPHANGIOMA|9170/0
C0024224|T191|ET|0000004535|AOD|lymphangiosarcoma|9170/3
C0024224|T191|PT|0000007599|CHV|lymphangiosarcoma|9170/3
C0024224|T191|ET|2007-1041|CSP|lymphangiosarcoma|9170/3
C0024224|T191|PT|MTHU046578|ICPC2ICD10ENG|lymphangioendothelial; sarcoma|9170/3
C0024224|T191|PT|MTHU065918|ICPC2ICD10ENG|sarcoma; lymphangioendothelial|9170/3
C0024224|T191|PT|10025223|MDR|Lymphangiosarcoma|9170/3
C0024224|T191|LLT|10025223|MDR|Lymphangiosarcoma|9170/3
C0024224|T191|LLT|10025225|MDR|Lymphangiosarcoma NOS|9170/3
C0024224|T191|HT|10025224|MDR|Lymphangiosarcomas|9170/3
C0024224|T191|PT|271558|MEDCIN|lymphangiosarcoma|9170/3
C0024224|T191|ET|D008204|MSH|Lymphangioendothelioma, Malignant|9170/3
C0024224|T191|PM|D008204|MSH|Lymphangioendotheliomas, Malignant|9170/3
C0024224|T191|MH|D008204|MSH|Lymphangiosarcoma|9170/3
C0024224|T191|PM|D008204|MSH|Lymphangiosarcomas|9170/3
C0024224|T191|PM|D008204|MSH|Malignant Lymphangioendothelioma|9170/3
C0024224|T191|PM|D008204|MSH|Malignant Lymphangioendotheliomas|9170/3
C0024224|T191|PN|NOCODE|MTH|lymphangiosarcoma|9170/3
C0024224|T191|SY|C3205|NCI|Lymphangioendothelial Sarcoma|9170/3
C0024224|T191|PT|C3205|NCI|Lymphangiosarcoma|9170/3
C0024224|T191|SY|C3205|NCI|Malignant Lymphangioendothelioma|9170/3
C0024224|T191|SY|C3205|NCI_CDISC|Lymphangioendothelial Sarcoma|9170/3
C0024224|T191|PT|C3205|NCI_CDISC|LYMPHANGIOSARCOMA, MALIGNANT|9170/3
C0024224|T191|SY|C3205|NCI_CDISC|Malignant Lymphangioendothelioma|9170/3
C0024224|T191|PT|CDR0000335070|NCI_NCI-GLOSS|lymphangiosarcoma|9170/3
C0024224|T191|SY|BBU1.|RCD|Lymphangioendothelial sarcoma|9170/3
C0024224|T191|PT|BBU1.|RCD|Lymphangiosarcoma|9170/3
C0024224|T191|AB|BBU1.|RCD|Malign lymphangioendothelioma|9170/3
C0024224|T191|SY|BBU1.|RCD|Malignant lymphangioendothelioma|9170/3
C0024224|T191|SY|63373002|SNOMEDCT_US|Lymphangioendothelial sarcoma|9170/3
C0024224|T191|SY|63373002|SNOMEDCT_US|Lymphangioendothelioma, malignant|9170/3
C0024224|T191|PT|403986008|SNOMEDCT_US|Lymphangiosarcoma|9170/3
C0024224|T191|PT|63373002|SNOMEDCT_US|Lymphangiosarcoma|9170/3
C0024224|T191|SY|63373002|SNOMEDCT_US|Malignant lymphangioendothelioma|9170/3
C0343089|T191|PT|0000030832|CHV|lymphangioma circumscriptum|9171/0
C0334543|T191|PT|MTHU014661|ICPC2ICD10ENG|capillary; lymphangioma|9171/0
C0334543|T191|PT|MTHU046583|ICPC2ICD10ENG|lymphangioma; capillary|9171/0
C0343089|T191|PT|C45485|NCI|Lymphangioma Circumscriptum|9171/0
C0334543|T191|PT|BBU2.|RCD|Capillary lymphangioma|9171/0
C0343089|T191|PT|X50Bo|RCD|Lymphangioma circumscriptum|9171/0
C0334543|T191|PT|11467009|SNOMEDCT_US|Capillary lymphangioma|9171/0
C0343089|T191|PT|238799002|SNOMEDCT_US|Lymphangioma circumscriptum|9171/0
C0205828|T191|DI|U001114|DXP|LYMPHANGIOMA, CAVERNOUS|9172/0
C0205828|T191|PT|MTHU015300|ICPC2ICD10ENG|cavernous; lymphangioma|9172/0
C0205828|T191|PT|MTHU046584|ICPC2ICD10ENG|lymphangioma; cavernous|9172/0
C0205828|T191|PM|D008202|MSH|Cavernous Lymphangioma|9172/0
C0205828|T191|PM|D008202|MSH|Cavernous Lymphangiomas|9172/0
C0205828|T191|PEP|D008202|MSH|Lymphangioma, Cavernous|9172/0
C0205828|T191|PM|D008202|MSH|Lymphangiomas, Cavernous|9172/0
C0205828|T191|PN|NOCODE|MTH|Cavernous lymphangioma|9172/0
C0205828|T191|PT|C53316|NCI|Cavernous Lymphangioma|9172/0
C0205828|T191|PT|BBU3.|RCD|Cavernous lymphangioma|9172/0
C0205828|T191|PT|89056007|SNOMEDCT_US|Cavernous lymphangioma|9172/0
C0206620|T191|PT|0059029|CCPSS|CYSTIC HYGROMA|9173/0
C0206620|T191|SY|0000020973|CHV|cystic hygroma|9173/0
C0206620|T191|SY|0000020973|CHV|cystic hygromas|9173/0
C0206620|T191|PT|0000020973|CHV|cystic lymphangioma|9173/0
C0206620|T191|SY|0000020973|CHV|cystic lymphangiomas|9173/0
C0206620|T191|SY|0000020973|CHV|hygroma|9173/0
C0206620|T191|SY|0000020973|CHV|hygromas|9173/0
C0206620|T191|PT|HP:0000476|HPO|Cystic hygroma|9173/0
C0206620|T191|SY|HP:0000476|HPO|Cystic hygroma of the neck|9173/0
C0206620|T191|PT|MTHU020765|ICPC2ICD10ENG|cystic; lymphangioma|9173/0
C0206620|T191|PT|MTHU036019|ICPC2ICD10ENG|hygroma|9173/0
C0206620|T191|PT|MTHU046585|ICPC2ICD10ENG|lymphangioma; cystic|9173/0
C0206620|T191|PTN|K72008|ICPC2P|cystic lymphangioma|9173/0
C0206620|T191|OPN|K99048|ICPC2P|cystic lymphangioma|9173/0
C0206620|T191|OP|K99048|ICPC2P|Lymphangioma;cystic|9173/0
C0206620|T191|PT|K72008|ICPC2P|Lymphangioma;cystic|9173/0
C0206620|T191|LLT|10011769|MDR|Cystic hygroma|9173/0
C0206620|T191|LLT|10058949|MDR|Cystic lymphangioma|9173/0
C0206620|T191|PT|10058949|MDR|Cystic lymphangioma|9173/0
C0206620|T191|LLT|10020543|MDR|Hygroma cystic|9173/0
C0206620|T191|PT|362060|MEDCIN|Cystic hygroma|9173/0
C0206620|T191|PM|D018191|MSH|Colli, Cystic Hygroma|9173/0
C0206620|T191|PM|D018191|MSH|Cystic Hygroma|9173/0
C0206620|T191|ET|D018191|MSH|Cystic Hygroma Colli|9173/0
C0206620|T191|PM|D018191|MSH|Cystic Hygromas|9173/0
C0206620|T191|PM|D018191|MSH|Cystic Lymphangioma|9173/0
C0206620|T191|PM|D018191|MSH|Cystic Lymphangiomas|9173/0
C0206620|T191|ET|D018191|MSH|Hygroma|9173/0
C0206620|T191|PM|D018191|MSH|Hygroma Colli, Cystic|9173/0
C0206620|T191|ET|D018191|MSH|Hygroma, Cystic|9173/0
C0206620|T191|PM|D018191|MSH|Hygromas|9173/0
C0206620|T191|PM|D018191|MSH|Hygromas, Cystic|9173/0
C0206620|T191|MH|D018191|MSH|Lymphangioma, Cystic|9173/0
C0206620|T191|PM|D018191|MSH|Lymphangiomas, Cystic|9173/0
C0206620|T191|PT|C3724|NCI|Cystic Hygroma|9173/0
C0206620|T191|SY|C3724|NCI|Cystic Lymphangioma|9173/0
C0206620|T191|SY|C3724|NCI|Hygroma|9173/0
C0206620|T191|PT|C3724|NCI_NICHD|Cystic Hygroma|9173/0
C0206620|T191|SY|C3724|NCI_NICHD|Cystic Lymphangioma|9173/0
C0206620|T191|SY|BBU4.|RCD|Cystic hygroma|9173/0
C0206620|T191|PT|BBU4.|RCD|Cystic lymphangioma|9173/0
C0206620|T191|SY|BBU4.|RCD|Hygroma|9173/0
C0206620|T191|SY|40225001|SNOMEDCT_US|Cystic hygroma|9173/0
C0206620|T191|PT|399882002|SNOMEDCT_US|Cystic hygroma|9173/0
C0206620|T191|PT|40225001|SNOMEDCT_US|Cystic lymphangioma|9173/0
C0206620|T191|PT|423984004|SNOMEDCT_US|Hygroma|9173/0
C0206620|T191|SY|40225001|SNOMEDCT_US|Hygroma|9173/0
C0206620|T191|IS|40225001|SNOMEDCT_US|Hygroma, NOS|9173/0
C0206620|T191|SY|423984004|SNOMEDCT_US|Non-neoplastic hygroma|9173/0
C0206620|T191|PT|1582|WHO|HYGROMA CYSTIC|9173/0
C0024223|T191|PT|MTHU046581|ICPC2ICD10ENG|lymphangiomyoma|9174/0
C0024223|T191|ET|D008203|MSH|Lymphangioleiomyoma|9174/0
C0024223|T191|PM|D008203|MSH|Lymphangioleiomyomas|9174/0
C0024223|T191|MH|D008203|MSH|Lymphangiomyoma|9174/0
C0024223|T191|PM|D008203|MSH|Lymphangiomyomas|9174/0
C0024223|T191|PT|C3204|NCI|Lymphangioleiomyoma|9174/0
C0024223|T191|SY|C3204|NCI|Lymphangiomyoma|9174/0
C0024223|T191|PT|BBU5.|RCD|Lymphangiomyoma|9174/0
C0024223|T191|PT|25239006|SNOMEDCT_US|Lymphangiomyoma|9174/0
C0751674|T191|PT|0000048475|CHV|lymphangioleiomyomatosis|9174/1
C0751674|T191|SY|0000048475|CHV|lymphangiomyomatosis|9174/1
C0751674|T191|AB|4009-0064|CSP|LAM|9174/1
C0751674|T191|PT|4009-0064|CSP|lymphangioleiomyomatosis|9174/1
C0751674|T191|ET|4009-0064|CSP|lymphangiomyomatosis|9174/1
C0751674|T191|ET|HP:0012798|HPO|Lymphangioleiomyomatosis|9174/1
C0751674|T191|AB|J84.81|ICD10CM|Lymphangioleiomyomatosis|9174/1
C0751674|T191|PT|J84.81|ICD10CM|Lymphangioleiomyomatosis|9174/1
C0751674|T191|ET|J84.81|ICD10CM|Lymphangiomyomatosis|9174/1
C0751674|T191|AB|516.4|ICD9CM|Lymphangioleiomyomatosis|9174/1
C0751674|T191|PT|516.4|ICD9CM|Lymphangioleiomyomatosis|9174/1
C0751674|T191|PT|sh99000736|LCH_NW|Lymphangiomyomatosis|9174/1
C0751674|T191|LLT|10049459|MDR|Lymphangioleiomyomatosis|9174/1
C0751674|T191|PT|10049459|MDR|Lymphangioleiomyomatosis|9174/1
C0751674|T191|LLT|10049462|MDR|Lymphangiomyomatosis|9174/1
C0751674|T191|PT|367668|MEDCIN|Lymphangioleiomyomatosis|9174/1
C0751674|T191|PT|31177|MEDCIN|lymphangiomyomatosis|9174/1
C0751674|T191|PM|D018192|MSH|Lymphangioleiomyomatoses|9174/1
C0751674|T191|MH|D018192|MSH|Lymphangioleiomyomatosis|9174/1
C0751674|T191|PM|D018192|MSH|Lymphangiomyomatoses|9174/1
C0751674|T191|ET|D018192|MSH|Lymphangiomyomatosis|9174/1
C0751674|T191|PN|NOCODE|MTH|Lymphangioleiomyomatosis|9174/1
C0751674|T191|ET|516.4|MTHICD9|Lymphangiomyomatosis|9174/1
C0751674|T191|AB|C3725|NCI|LAM|9174/1
C0751674|T191|PT|C3725|NCI|Lymphangioleiomyomatosis|9174/1
C0751674|T191|SY|C3725|NCI|Lymphangiomyomatosis|9174/1
C0751674|T191|DN|C3725|NCI_CTRP|Lymphangioleiomyomatosis|9174/1
C0751674|T191|AB|CDR0000532373|PDQ|LAM|9174/1
C0751674|T191|PT|CDR0000532373|PDQ|lymphangioleiomyomatosis|9174/1
C0751674|T191|LV|CDR0000532373|PDQ|Lymphangiomyomatosis|9174/1
C0751674|T191|PT|BBU6.|RCD|Lymphangiomyomatosis|9174/1
C0751674|T191|SY|73017001|SNOMEDCT_US|Lymphangioleiomyomatosis|9174/1
C0751674|T191|PT|73017001|SNOMEDCT_US|Lymphangiomyomatosis|9174/1
C0334544|T191|PT|MTHU034084|ICPC2ICD10ENG|hemolymphangioma|9175/0
C0334544|T191|PT|C66792|NCI|Hemolymphangioma|9175/0
C0334544|T191|SY|C66792|NCI|Lymphangioma with Hemorrhage|9175/0
C0334544|T191|PT|BBU7.|RCD|Haemolymphangioma|9175/0
C0334544|T191|PT|BBU7.|RCDAE|Hemolymphangioma|9175/0
C0334544|T191|PTGB|8241005|SNOMEDCT_US|Haemolymphangioma|9175/0
C0334544|T191|PT|8241005|SNOMEDCT_US|Hemolymphangioma|9175/0
C0029440|T191|ET|0000004554|AOD|osteoma|9180/0
C0029440|T191|PT|0014185|CCPSS|OSTEOMA|9180/0
C0029440|T191|PT|0000009085|CHV|osteoma|9180/0
C0029440|T191|SY|0000009085|CHV|osteomas|9180/0
C0029440|T191|PT|NOCODE|COSTAR|Osteoma|9180/0
C0029440|T191|DI|U001350|DXP|OSTEOMA|9180/0
C0029440|T191|PT|HP:0100246|HPO|Osteoma|9180/0
C0029440|T191|PT|L71010|ICPC2P|Osteoma|9180/0
C0029440|T191|PTN|L71010|ICPC2P|osteoma|9180/0
C0029440|T191|LLT|10031249|MDR|Osteoma|9180/0
C0029440|T191|PT|10031249|MDR|Osteoma|9180/0
C0029440|T191|PT|31714|MEDCIN|benign osteoma of bone|9180/0
C0029440|T191|MH|D010016|MSH|Osteoma|9180/0
C0029440|T191|PM|D010016|MSH|Osteomas|9180/0
C1332523|T191|PN|NOCODE|MTH|Benign Osteogenic Neoplasm|9180/0
C1332523|T191|SY|C6602|NCI|Benign Osseous Neoplasm|9180/0
C1332523|T191|SY|C6602|NCI|Benign Osseous Tumor|9180/0
C1332523|T191|PT|C6602|NCI|Benign Osteogenic Neoplasm|9180/0
C1332523|T191|SY|C6602|NCI|Benign Osteogenic Tumor|9180/0
C0029440|T191|PT|C3296|NCI|Osteoma|9180/0
C0029440|T191|PT|C3296|NCI_CDISC|OSTEOMA, BENIGN|9180/0
C0029440|T191|PT|Xa9AU|RCD|Osteoma|9180/0
C0029440|T191|OP|BBV0.|RCDSY|Osteoma NOS|9180/0
C1332523|T191|PT|726115006|SNOMEDCT_US|Benign osteogenic neoplasm|9180/0
C1332523|T191|SY|726115006|SNOMEDCT_US|Benign osteogenic tumor|9180/0
C1332523|T191|SYGB|726115006|SNOMEDCT_US|Benign osteogenic tumour|9180/0
C0029440|T191|OAS|154611005|SNOMEDCT_US|Osteoma|9180/0
C0029440|T191|OAS|187899007|SNOMEDCT_US|Osteoma|9180/0
C0029440|T191|PT|83612000|SNOMEDCT_US|Osteoma|9180/0
C0029440|T191|OAS|188904008|SNOMEDCT_US|Osteoma|9180/0
C0029440|T191|OAP|302858007|SNOMEDCT_US|Osteoma|9180/0
C0029440|T191|OAS|269638002|SNOMEDCT_US|Osteoma|9180/0
C0029440|T191|SY|83612000|SNOMEDCT_US|Osteoma, no ICD-O subtype|9180/0
C0029440|T191|SY|83612000|SNOMEDCT_US|Osteoma, no International Classification of Diseases for Oncology subtype|9180/0
C0029440|T191|IS|83612000|SNOMEDCT_US|Osteoma, NOS|9180/0
C0029440|T191|PT|1412|WHO|OSTEOMA|9180/0
C0029463|T191|ET|0000004536|AOD|osteosarcoma|9180/3
C0029463|T191|PT|1001695|CCPSS|OSTEOSARCOMA|9180/3
C0029463|T191|PT|0000009099|CHV|bone sarcoma|9180/3
C0029463|T191|SY|0000009099|CHV|bone sarcomas|9180/3
C0029463|T191|SY|0000009099|CHV|osteochondrosarcoma|9180/3
C0029463|T191|SY|0000009099|CHV|osteogenic sarcoma|9180/3
C0029463|T191|SY|0000009099|CHV|osteosarcoma|9180/3
C0029463|T191|SY|0000009099|CHV|osteosarcomas|9180/3
C0029463|T191|PT|NOCODE|COSTAR|Osteogenic Sarcoma|9180/3
C0029463|T191|PT|U000495|COSTAR|OSTEOSARCOMA|9180/3
C0029463|T191|ET|2019-1578|CSP|osteochondrosarcoma|9180/3
C0029463|T191|ET|2019-1578|CSP|osteogenic sarcoma|9180/3
C0029463|T191|ET|2019-1578|CSP|osteoid sarcoma|9180/3
C0029463|T191|PT|2019-1578|CSP|osteosarcoma|9180/3
C0029463|T191|GT|SARCOMA BONE|CST|SARCOMA OSTEOGENIC|9180/3
C0029463|T191|SY|NOCODE|DXP|BONE CANCER, OSTEOGENIC SARCOMA|9180/3
C0029463|T191|DI|U001349|DXP|OSTEOGENIC SARCOMA|9180/3
C0029463|T191|SY|NOCODE|DXP|OSTEOSARCOMA|9180/3
C0029463|T191|SY|HP:0002669|HPO|Bone cell cancer|9180/3
C0029463|T191|SY|HP:0002669|HPO|Osteogenic sarcoma|9180/3
C0029463|T191|PT|HP:0002669|HPO|Osteosarcoma|9180/3
C0029463|T191|PTN|L71018|ICPC2P|osteosarcoma|9180/3
C0029463|T191|PT|L71018|ICPC2P|Osteosarcoma|9180/3
C0029463|T191|PT|sh85095987|LCH_NW|Osteosarcoma|9180/3
C0029463|T191|LLT|10031244|MDR|Osteogenic sarcoma|9180/3
C0029463|T191|LLT|10031291|MDR|Osteosarcoma|9180/3
C0029463|T191|PT|10031291|MDR|Osteosarcoma|9180/3
C0029463|T191|LLT|10031295|MDR|Osteosarcoma NOS|9180/3
C0029463|T191|LLT|10039496|MDR|Sarcoma osteogenic|9180/3
C0029463|T191|ET|169|MEDLINEPLUS|Osteosarcoma|9180/3
C0029463|T191|ET|D012516|MSH|Osteogenic Sarcoma|9180/3
C0029463|T191|PM|D012516|MSH|Osteogenic Sarcomas|9180/3
C0029463|T191|MH|D012516|MSH|Osteosarcoma|9180/3
C0029463|T191|ET|D012516|MSH|Osteosarcoma Tumor|9180/3
C0029463|T191|PM|D012516|MSH|Osteosarcoma Tumors|9180/3
C0029463|T191|PM|D012516|MSH|Osteosarcomas|9180/3
C0029463|T191|ET|D012516|MSH|Sarcoma, Osteogenic|9180/3
C0029463|T191|PM|D012516|MSH|Sarcomas, Osteogenic|9180/3
C0029463|T191|PM|D012516|MSH|Tumor, Osteosarcoma|9180/3
C0029463|T191|PM|D012516|MSH|Tumors, Osteosarcoma|9180/3
C0029463|T191|PN|NOCODE|MTH|Osteosarcoma|9180/3
C0029463|T191|SY|C9145|NCI|Osteogenic Sarcoma|9180/3
C0029463|T191|PT|C9145|NCI|Osteosarcoma|9180/3
C0029463|T191|SY|C9145|NCI_CDISC|Osteogenic Sarcoma|9180/3
C0029463|T191|PT|C9145|NCI_CDISC|OSTEOSARCOMA, MALIGNANT|9180/3
C0029463|T191|PT|C9145|NCI_CPTAC|Osteosarcoma|9180/3
C0029463|T191|PT|10031291|NCI_CTEP-SDC|Osteosarcoma|9180/3
C0029463|T191|DN|C9145|NCI_CTRP|Osteosarcoma|9180/3
C0029463|T191|PT|C9145|NCI_CTRP|Osteosarcoma|9180/3
C0029463|T191|PT|CDR0000044069|NCI_NCI-GLOSS|osteogenic sarcoma|9180/3
C0029463|T191|PT|CDR0000045395|NCI_NCI-GLOSS|osteosarcoma|9180/3
C0029463|T191|PT|C9145|NCI_NICHD|Osteosarcoma|9180/3
C0029463|T191|SY|CDR0000041729|PDQ|osteogenic sarcoma|9180/3
C0029463|T191|ET|CDR0000041729|PDQ|Osteosarcoma|9180/3
C0029463|T191|PSC|CDR0000041729|PDQ|osteosarcoma|9180/3
C0029463|T191|SY|CDR0000041729|PDQ|sarcoma, osteogenic|9180/3
C0029463|T191|SY|Xa9AV|RCD|Osteochondrosarcoma|9180/3
C0029463|T191|SY|Xa9AV|RCD|Osteogenic sarcoma|9180/3
C0029463|T191|PT|Xa9AV|RCD|Osteosarcoma|9180/3
C0029463|T191|SY|Xa9AV|RCDSY|Osteosarcoma NOS|9180/3
C0029463|T191|SY|21708004|SNOMEDCT_US|Osteochondrosarcoma|9180/3
C0029463|T191|SY|21708004|SNOMEDCT_US|Osteogenic sarcoma|9180/3
C0029463|T191|IS|21708004|SNOMEDCT_US|Osteogenic sarcoma, NOS|9180/3
C0029463|T191|OAP|189878003|SNOMEDCT_US|Osteosarcoma|9180/3
C0029463|T191|OAS|408387006|SNOMEDCT_US|Osteosarcoma|9180/3
C0029463|T191|OF|189878003|SNOMEDCT_US|Osteosarcoma|9180/3
C0029463|T191|PT|21708004|SNOMEDCT_US|Osteosarcoma|9180/3
C0029463|T191|SY|307576001|SNOMEDCT_US|Osteosarcoma|9180/3
C0029463|T191|OAP|408387006|SNOMEDCT_US|Osteosarcoma - disorder|9180/3
C0029463|T191|SY|307576001|SNOMEDCT_US|Osteosarcoma - disorder|9180/3
C0029463|T191|SY|21708004|SNOMEDCT_US|Osteosarcoma, no ICD-O subtype|9180/3
C0029463|T191|SY|21708004|SNOMEDCT_US|Osteosarcoma, no International Classification of Diseases for Oncology subtype|9180/3
C0029463|T191|IS|21708004|SNOMEDCT_US|Osteosarcoma, NOS|9180/3
C3838970|T191|PT|703693004|SNOMEDCT_US|Post-radiation osteosarcoma|9180/3
C0279603|T191|PT|MTHU016328|ICPC2ICD10ENG|chondroblastic; osteosarcoma|9181/3
C0279603|T191|PT|MTHU056360|ICPC2ICD10ENG|osteosarcoma; chondroblastic|9181/3
C0279603|T191|LLT|10008740|MDR|Chondrosarcomatous osteosarcoma|9181/3
C0279603|T191|SY|C4021|NCI|Chondroblastic Osteogenic Sarcoma|9181/3
C0279603|T191|PT|C4021|NCI|Chondroblastic Osteosarcoma|9181/3
C0279603|T191|DN|C4021|NCI_CTRP|Chondroblastic Osteosarcoma|9181/3
C0279603|T191|SY|CDR0000039885|PDQ|chondroblastic osteogenic sarcoma|9181/3
C0279603|T191|SY|CDR0000039885|PDQ|chondroblastic osteosarcoma|9181/3
C0279603|T191|SY|CDR0000039885|PDQ|chondrosarcomatous osteogenic sarcoma|9181/3
C0279603|T191|PT|CDR0000039885|PDQ|chondrosarcomatous osteosarcoma|9181/3
C0279603|T191|SY|CDR0000039885|PDQ|osteogenic sarcoma, chondroblastic|9181/3
C0279603|T191|SY|CDR0000039885|PDQ|osteogenic sarcoma, chondrosarcomatous|9181/3
C0279603|T191|SY|CDR0000039885|PDQ|osteosarcoma, chondroblastic|9181/3
C0279603|T191|SY|CDR0000039885|PDQ|osteosarcoma, chondrosarcomatous|9181/3
C0279603|T191|SY|CDR0000039885|PDQ|sarcoma, osteogenic, chondrosarcomatous|9181/3
C0279603|T191|PT|BBV2.|RCD|Chondroblastic osteosarcoma|9181/3
C0279603|T191|PT|76312009|SNOMEDCT_US|Chondroblastic osteosarcoma|9181/3
C0279602|T191|PT|MTHU028174|ICPC2ICD10ENG|fibroblastic; osteosarcoma|9182/3
C0279602|T191|PT|MTHU056361|ICPC2ICD10ENG|osteosarcoma; fibroblastic|9182/3
C0279602|T191|SY|C4020|NCI|Fibroblastic Osteogenic Sarcoma|9182/3
C0279602|T191|PT|C4020|NCI|Fibroblastic Osteosarcoma|9182/3
C0279602|T191|SY|C4020|NCI|Fibrosarcomatous Osteogenic Sarcoma|9182/3
C0279602|T191|SY|C4020|NCI|Fibrosarcomatous Osteosarcoma|9182/3
C0279602|T191|PT|C4020|NCI_CDISC|FIBROSARCOMA, OSTEOGENIC, MALIGNANT|9182/3
C0279602|T191|SY|C4020|NCI_CDISC|Osteogenic Fibrosarcoma|9182/3
C0279602|T191|DN|C4020|NCI_CTRP|Fibroblastic Osteosarcoma|9182/3
C0279602|T191|SY|CDR0000039884|PDQ|fibroblastic osteogenic sarcoma|9182/3
C0279602|T191|SY|CDR0000039884|PDQ|fibroblastic osteosarcoma|9182/3
C0279602|T191|SY|CDR0000039884|PDQ|fibrosarcomatous osteogenic sarcoma|9182/3
C0279602|T191|PT|CDR0000039884|PDQ|fibrosarcomatous osteosarcoma|9182/3
C0279602|T191|SY|CDR0000039884|PDQ|osteogenic sarcoma, fibroblastic|9182/3
C0279602|T191|SY|CDR0000039884|PDQ|osteogenic sarcoma, fibrosarcomatous|9182/3
C0279602|T191|SY|CDR0000039884|PDQ|osteosarcoma, fibroblastic|9182/3
C0279602|T191|SY|CDR0000039884|PDQ|osteosarcoma, fibrosarcomatous|9182/3
C0279602|T191|SY|CDR0000039884|PDQ|sarcoma, osteogenic fibroblastic|9182/3
C0279602|T191|PT|BBV3.|RCD|Fibroblastic osteosarcoma|9182/3
C0279602|T191|SY|BBV3.|RCD|Osteofibrosarcoma|9182/3
C0279602|T191|PT|12690005|SNOMEDCT_US|Fibroblastic osteosarcoma|9182/3
C0279602|T191|SY|12690005|SNOMEDCT_US|Osteofibrosarcoma|9182/3
C0259782|T191|PT|MTHU056365|ICPC2ICD10ENG|osteosarcoma; telangiectatic|9183/3
C0259782|T191|PT|MTHU073642|ICPC2ICD10ENG|telangiectatic; osteosarcoma|9183/3
C0259782|T191|LLT|10043195|MDR|Telangiectatic osteosarcoma|9183/3
C0259782|T191|SY|C3902|NCI|Malignant Bone Aneurysm|9183/3
C0259782|T191|SY|C3902|NCI|Telangiectatic Osteogenic Sarcoma|9183/3
C0259782|T191|PT|C3902|NCI|Telangiectatic Osteosarcoma|9183/3
C0259782|T191|DN|C3902|NCI_CTRP|Telangiectatic Osteosarcoma|9183/3
C0259782|T191|SY|CDR0000039888|PDQ|Malignant Bone Aneurysm|9183/3
C0259782|T191|SY|CDR0000039888|PDQ|osteogenic sarcoma, telangiectatic|9183/3
C0259782|T191|SY|CDR0000039888|PDQ|osteosarcoma, telangiectatic|9183/3
C0259782|T191|SY|CDR0000039888|PDQ|sarcoma, osteogenic telangiectatic|9183/3
C0259782|T191|SY|CDR0000039888|PDQ|telangiectatic osteogenic sarcoma|9183/3
C0259782|T191|PT|CDR0000039888|PDQ|telangiectatic osteosarcoma|9183/3
C0259782|T191|PT|BBV4.|RCD|Telangiectatic osteosarcoma|9183/3
C0259782|T191|PT|78453009|SNOMEDCT_US|Telangiectatic osteosarcoma|9183/3
C0334546|T191|PT|MTHU056359|ICPC2ICD10ENG|osteosarcoma; in Paget's disease of bone|9184/3
C1335148|T191|PT|MTHU057031|ICPC2ICD10ENG|Paget; osteosarcoma|9184/3
C0334546|T191|PT|230792|MEDCIN|osteosarcoma in Paget disease of bone|9184/3
C1335148|T191|SY|C6469|NCI|Osteosarcoma Arising in Bone Paget's Disease|9184/3
C1335148|T191|SY|C6469|NCI|Osteosarcoma Arising in Osseous Paget's Disease|9184/3
C1335148|T191|SY|C6469|NCI|Osteosarcoma Arising in Osteitis Deformans|9184/3
C1335148|T191|PT|C6469|NCI|Osteosarcoma Arising in Paget Disease of Bone|9184/3
C1335148|T191|SY|C6469|NCI|Osteosarcoma Arising in Paget's Disease of Bone|9184/3
C1335148|T191|SY|C6469|NCI|Paget Osteosarcoma|9184/3
C1335148|T191|SY|C6469|NCI|Paget's Osteosarcoma|9184/3
C1710042|T191|SY|C53704|NCI|Secondary Bone Osteosarcoma|9184/3
C1710042|T191|PT|C53704|NCI|Secondary Osteosarcoma|9184/3
C0334546|T191|AB|BBV5.|RCD|Osteosarc in Paget's dis bone|9184/3
C0334546|T191|PT|BBV5.|RCD|Osteosarcoma in Paget's disease of bone|9184/3
C0334546|T191|SY|33681003|SNOMEDCT_US|Osteosarcoma in Paget disease of bone|9184/3
C0334546|T191|PT|33681003|SNOMEDCT_US|Osteosarcoma in Paget's disease of bone|9184/3
C1710042|T191|PT|703692009|SNOMEDCT_US|Secondary osteosarcoma|9184/3
C0279622|T191|PT|MTHU056363|ICPC2ICD10ENG|osteosarcoma; small cell|9185/3
C0279622|T191|PT|MTHU041513|ICPC2ICD10ENG|small cell; osteosarcoma|9185/3
C0279622|T191|PT|230756|MEDCIN|small cell sarcoma of bone|9185/3
C0279622|T191|SY|C4023|NCI|Small Cell Osteogenic Sarcoma|9185/3
C0279622|T191|PT|C4023|NCI|Small Cell Osteosarcoma|9185/3
C0279622|T191|OP|CDR0000039907|PDQ|small cell bone sarcoma|9185/3
C0279622|T191|SY|CDR0000039907|PDQ|small cell osteogenic sarcoma|9185/3
C0279622|T191|SY|CDR0000039907|PDQ|small cell osteosarcoma|9185/3
C0279622|T191|PT|X77pA|RCD|Small cell osteosarcoma|9185/3
C0279622|T191|OP|BBVA.|RCDSY|Small cell osteosarcoma|9185/3
C0279622|T191|SY|12302002|SNOMEDCT_US|Round cell osteosarcoma|9185/3
C0279622|T191|PT|12302002|SNOMEDCT_US|Small cell osteosarcoma|9185/3
C1266166|T191|LLT|10002236|MDR|Anaplastic osteosarcoma|9186/3
C1266166|T191|PT|90258|MEDCIN|undifferentiated sarcoma of bone|9186/3
C1266166|T191|SY|C35870|NCI|Central Osteosarcoma|9186/3
C1266166|T191|SY|C35870|NCI|Conventional Central Osteosarcoma|9186/3
C1266166|T191|PT|C35870|NCI|Conventional Osteosarcoma|9186/3
C1266166|T191|SY|C35870|NCI|Intracortical Osteogenic Sarcoma|9186/3
C1266166|T191|SY|C35870|NCI|Intracortical Osteosarcoma|9186/3
C1266166|T191|SY|C35870|NCI|Medullary Osteosarcoma|9186/3
C1266166|T191|DN|C35870|NCI_CTRP|Conventional Osteosarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|anaplastic osteogenic sarcoma|9186/3
C1266166|T191|PT|CDR0000039890|PDQ|anaplastic osteosarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|Central Osteosarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|Conventional Central Osteosarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|Conventional Osteosarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|Intracortical Osteogenic Sarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|Intracortical Osteosarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|Medullary Osteosarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|osteogenic sarcoma, anaplastic|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|osteogenic sarcoma, undifferentiated|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|osteosarcoma, anaplastic|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|osteosarcoma, undifferentiated|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|sarcoma, osteogenic anaplastic|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|sarcoma, osteogenic undifferentiated|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|undifferentiated osteogenic sarcoma|9186/3
C1266166|T191|SY|CDR0000039890|PDQ|undifferentiated osteosarcoma|9186/3
C1266166|T191|PT|128770002|SNOMEDCT_US|Central osteosarcoma|9186/3
C1266166|T191|SY|128770002|SNOMEDCT_US|Conventional central osteosarcoma|9186/3
C1266166|T191|PT|128774006|SNOMEDCT_US|Intracortical osteosarcoma|9186/3
C1266166|T191|SY|128770002|SNOMEDCT_US|Medullary osteosarcoma|9186/3
C1266163|T191|PN|NOCODE|MTH|Intraosseous well differentiated osteosarcoma|9187/3
C3814534|T191|PN|NOCODE|MTH|Low grade central osteosarcoma|9187/3
C1266163|T191|SY|C6474|NCI|Intraosseous Well-Differentiated Osteogenic Sarcoma|9187/3
C1266163|T191|SY|C6474|NCI|Intraosseous Well-Differentiated Osteosarcoma|9187/3
C1266163|T191|PT|C6474|NCI|Low Grade Central Osteosarcoma|9187/3
C1266163|T191|SY|C6474|NCI|Low Grade Intramedullary Osteosarcoma|9187/3
C1266163|T191|SY|C6474|NCI|Low-Grade Intramedullary Osteosarcoma|9187/3
C1266163|T191|SY|128771003|SNOMEDCT_US|Intraosseous low grade osteosarcoma|9187/3
C1266163|T191|PT|128771003|SNOMEDCT_US|Intraosseous well differentiated osteosarcoma|9187/3
C3814534|T191|PT|703694005|SNOMEDCT_US|Low grade central osteosarcoma|9187/3
C0029441|T191|PT|0000009086|CHV|osteoid osteoma|9191/0
C0029441|T191|SY|0000009086|CHV|osteoid osteomas|9191/0
C0029441|T191|SY|0000009086|CHV|osteoma osteoid|9191/0
C0029441|T191|PT|NOCODE|COSTAR|Osteoid Osteoma|9191/0
C0029441|T191|PT|HP:0030433|HPO|Osteoid osteoma|9191/0
C0029441|T191|PT|31494|MEDCIN|benign osteoid osteoma of bone|9191/0
C0029441|T191|ET|D010017|MSH|Osteoid Osteoma|9191/0
C0029441|T191|PM|D010017|MSH|Osteoid Osteomas|9191/0
C0029441|T191|MH|D010017|MSH|Osteoma, Osteoid|9191/0
C0029441|T191|PM|D010017|MSH|Osteomas, Osteoid|9191/0
C0029441|T191|PN|NOCODE|MTH|Osteoid osteoma|9191/0
C0029441|T191|PT|C3297|NCI|Osteoid Osteoma|9191/0
C0029441|T191|PT|Xa9AW|RCD|Osteoid osteoma|9191/0
C0029441|T191|OP|BBV7.|RCDSY|Osteoid osteoma NOS|9191/0
C0029441|T191|PT|71666005|SNOMEDCT_US|Osteoid osteoma|9191/0
C0029441|T191|OAP|302859004|SNOMEDCT_US|Osteoid osteoma|9191/0
C0029441|T191|IS|71666005|SNOMEDCT_US|Osteoid osteoma, NOS|9191/0
C0206642|T191|SY|0000020990|CHV|osteosarcomas periosteal|9192/3
C0206642|T191|PT|0000020990|CHV|parosteal osteosarcoma|9192/3
C0206642|T191|SY|0000020990|CHV|periosteal osteosarcoma|9192/3
C0206642|T191|PT|MTHU040708|ICPC2ICD10ENG|juxtacortical; osteosarcoma|9192/3
C0206642|T191|PT|MTHU056362|ICPC2ICD10ENG|osteosarcoma; juxtacortical|9192/3
C0206642|T191|PT|MTHU056364|ICPC2ICD10ENG|osteosarcoma; parosteal|9192/3
C0206642|T191|PT|MTHU057942|ICPC2ICD10ENG|parosteal; osteosarcoma|9192/3
C0206642|T191|PT|39717|MEDCIN|juxtacortical osteosarcoma|9192/3
C0206642|T191|PM|D018217|MSH|Juxtacortical Osteosarcoma|9192/3
C0206642|T191|PM|D018217|MSH|Juxtacortical Osteosarcomas|9192/3
C0206642|T191|MH|D018217|MSH|Osteosarcoma, Juxtacortical|9192/3
C0206642|T191|PM|D018217|MSH|Osteosarcomas, Juxtacortical|9192/3
C0206642|T191|PN|NOCODE|MTH|Parosteal Osteosarcoma|9192/3
C0206642|T191|SY|C8969|NCI|Juxtacortical Osteogenic Sarcoma|9192/3
C0206642|T191|SY|C8969|NCI|Juxtacortical Osteosarcoma|9192/3
C0206642|T191|SY|C8969|NCI|Parosteal Osteogenic Sarcoma|9192/3
C0206642|T191|PT|C8969|NCI|Parosteal Osteosarcoma|9192/3
C0206642|T191|AB|BBV6.|RCD|Juxtacortical osteogenic sarc|9192/3
C0206642|T191|SY|BBV6.|RCD|Juxtacortical osteogenic sarcoma|9192/3
C0206642|T191|PT|BBV6.|RCD|Juxtacortical osteosarcoma|9192/3
C0206642|T191|SY|BBV6.|RCD|Parosteal osteosarcoma|9192/3
C0206642|T191|IS|91242000|SNOMEDCT_US|Juxtacortical osteogenic sarcoma|9192/3
C0206642|T191|OAP|189879006|SNOMEDCT_US|Juxtacortical osteosarcoma|9192/3
C0206642|T191|OAP|91242000|SNOMEDCT_US|Juxtacortical osteosarcoma|9192/3
C0206642|T191|SY|128918008|SNOMEDCT_US|Juxtacortical osteosarcoma|9192/3
C0206642|T191|IS|91242000|SNOMEDCT_US|Juxtacortical osteosarcoma -RETIRED-|9192/3
C0206642|T191|OF|91242000|SNOMEDCT_US|Juxtacortical osteosarcoma -RETIRED-|9192/3
C0206642|T191|PT|128918008|SNOMEDCT_US|Parosteal osteosarcoma|9192/3
C0206642|T191|IS|91242000|SNOMEDCT_US|Parosteal osteosarcoma|9192/3
C1377843|T191|PN|NOCODE|MTH|Periosteal Osteosarcoma|9193/3
C1377843|T191|SY|C8970|NCI|Juxtacortical Chondroblastic Osteosarcoma|9193/3
C1377843|T191|PT|C8970|NCI|Periosteal Osteosarcoma|9193/3
C1377843|T191|SY|BBV6.|RCD|Periosteal osteogenic sarcoma|9193/3
C1377843|T191|IS|91242000|SNOMEDCT_US|Periosteal osteogenic sarcoma|9193/3
C1377843|T191|IS|91242000|SNOMEDCT_US|Periosteal osteosarcoma|9193/3
C1377843|T191|PT|128772005|SNOMEDCT_US|Periosteal osteosarcoma|9193/3
C1266165|T191|PT|C53958|NCI|High Grade Surface Osteosarcoma|9194/3
C1266165|T191|PT|128773000|SNOMEDCT_US|High grade surface osteosarcoma|9194/3
C1266166|T191|LLT|10002236|MDR|Anaplastic osteosarcoma|9195/3
C1266166|T191|PT|90258|MEDCIN|undifferentiated sarcoma of bone|9195/3
C1266166|T191|SY|C35870|NCI|Central Osteosarcoma|9195/3
C1266166|T191|SY|C35870|NCI|Conventional Central Osteosarcoma|9195/3
C1266166|T191|PT|C35870|NCI|Conventional Osteosarcoma|9195/3
C1266166|T191|SY|C35870|NCI|Intracortical Osteogenic Sarcoma|9195/3
C1266166|T191|SY|C35870|NCI|Intracortical Osteosarcoma|9195/3
C1266166|T191|SY|C35870|NCI|Medullary Osteosarcoma|9195/3
C1266166|T191|DN|C35870|NCI_CTRP|Conventional Osteosarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|anaplastic osteogenic sarcoma|9195/3
C1266166|T191|PT|CDR0000039890|PDQ|anaplastic osteosarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|Central Osteosarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|Conventional Central Osteosarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|Conventional Osteosarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|Intracortical Osteogenic Sarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|Intracortical Osteosarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|Medullary Osteosarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|osteogenic sarcoma, anaplastic|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|osteogenic sarcoma, undifferentiated|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|osteosarcoma, anaplastic|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|osteosarcoma, undifferentiated|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|sarcoma, osteogenic anaplastic|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|sarcoma, osteogenic undifferentiated|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|undifferentiated osteogenic sarcoma|9195/3
C1266166|T191|SY|CDR0000039890|PDQ|undifferentiated osteosarcoma|9195/3
C1266166|T191|PT|128770002|SNOMEDCT_US|Central osteosarcoma|9195/3
C1266166|T191|SY|128770002|SNOMEDCT_US|Conventional central osteosarcoma|9195/3
C1266166|T191|PT|128774006|SNOMEDCT_US|Intracortical osteosarcoma|9195/3
C1266166|T191|SY|128770002|SNOMEDCT_US|Medullary osteosarcoma|9195/3
C0029417|T191|PT|0000009071|CHV|osteoblastoma|9200/0
C0029417|T191|SY|NOCODE|DXP|FIBROMA, OSTEOGENIC, OF BONE|9200/0
C0029417|T191|DI|U001345|DXP|OSTEOBLASTOMA, BENIGN|9200/0
C0029417|T191|SY|NOCODE|DXP|OSTEOID OSTEOMA, GIANT|9200/0
C0029417|T191|PT|HP:0011846|HPO|Osteoblastoma|9200/0
C0029417|T191|LLT|10004430|MDR|Benign osteoblastoma|9200/0
C0029417|T191|ET|D018215|MSH|Giant Osteoid Osteoma|9200/0
C0029417|T191|PM|D018215|MSH|Giant Osteoid Osteomas|9200/0
C0029417|T191|MH|D018215|MSH|Osteoblastoma|9200/0
C0029417|T191|PM|D018215|MSH|Osteoblastomas|9200/0
C0029417|T191|PM|D018215|MSH|Osteoid Osteoma, Giant|9200/0
C0029417|T191|PM|D018215|MSH|Osteoid Osteomas, Giant|9200/0
C0029417|T191|ET|D018215|MSH|Osteoma, Giant Osteoid|9200/0
C0029417|T191|PM|D018215|MSH|Osteomas, Giant Osteoid|9200/0
C0029417|T191|PN|NOCODE|MTH|Osteoblastoma|9200/0
C0029417|T191|SY|C3294|NCI|Giant Osteoid Osteoma|9200/0
C0029417|T191|SY|C3294|NCI|Ossifying Giant Cell Tumor|9200/0
C0029417|T191|PT|C3294|NCI|Osteoblastoma|9200/0
C0029417|T191|SY|C3294|NCI_CDISC|Giant Osteoid Osteoma|9200/0
C0029417|T191|SY|C3294|NCI_CDISC|Ossifying Giant Cell Tumor|9200/0
C0029417|T191|PT|C3294|NCI_CDISC|OSTEOBLASTOMA, BENIGN|9200/0
C0029417|T191|SY|BBV8.|RCD|Giant osteoid osteoma|9200/0
C0029417|T191|SY|BBV8.|RCD|Osteoblastoma|9200/0
C0029417|T191|SY|55333008|SNOMEDCT_US|Giant osteoid osteoma|9200/0
C0029417|T191|PT|55333008|SNOMEDCT_US|Osteoblastoma|9200/0
C0029417|T191|IS|55333008|SNOMEDCT_US|Osteoblastoma, NOS|9200/0
C0334547|T191|PT|C66796|NCI|Aggressive Osteoblastoma|9200/1
C0334547|T191|PT|X77pD|RCD|Aggressive osteoblastoma|9200/1
C0334547|T191|PT|70511009|SNOMEDCT_US|Aggressive osteoblastoma|9200/1
C0029423|T191|PT|0000009076|CHV|cartilaginous exostosis|9210/0
C0029423|T191|SY|0000009076|CHV|ecchondroma|9210/0
C0029423|T191|SY|0000009076|CHV|exostosis|9210/0
C0029423|T191|SY|0000009076|CHV|osteochondroma|9210/0
C0029423|T191|SY|0000009076|CHV|osteochondromas|9210/0
C0029423|T191|PT|NOCODE|COSTAR|Osteochondroma|9210/0
C0029423|T191|SY|HP:0030431|HPO|Osteocartilaginous exostoses|9210/0
C0029423|T191|PT|HP:0030431|HPO|Osteochondroma|9210/0
C0029423|T191|SY|HP:0030431|HPO|Osteochondromas|9210/0
C0029423|T191|PT|L97016|ICPC2P|Osteochondroma|9210/0
C0029423|T191|PTN|L97016|ICPC2P|osteochondroma|9210/0
C0029423|T191|OP|L71019|ICPC2P|Osteochondroma|9210/0
C0029423|T191|PT|U005373|LCH|Osteochondroma|9210/0
C0029423|T191|PT|sh85095962|LCH_NW|Osteochondroma|9210/0
C0029423|T191|PT|10059587|MDR|Osteochondroma|9210/0
C0029423|T191|LLT|10059587|MDR|Osteochondroma|9210/0
C0029423|T191|PT|31490|MEDCIN|benign chondroma of bone|9210/0
C0029423|T191|PM|D015831|MSH|Cartilaginous Exostoses|9210/0
C0029423|T191|PM|D015831|MSH|Cartilaginous Exostosis|9210/0
C0029423|T191|ET|D015831|MSH|Chondrosteoma|9210/0
C0029423|T191|PM|D015831|MSH|Chondrosteomas|9210/0
C0029423|T191|PM|D015831|MSH|Exostoses, Cartilaginous|9210/0
C0029423|T191|PM|D015831|MSH|Exostoses, Osteocartilaginous|9210/0
C0029423|T191|ET|D015831|MSH|Exostosis, Cartilaginous|9210/0
C0029423|T191|ET|D015831|MSH|Exostosis, Osteocartilaginous|9210/0
C0029423|T191|PM|D015831|MSH|Osteocartilaginous Exostoses|9210/0
C0029423|T191|PM|D015831|MSH|Osteocartilaginous Exostosis|9210/0
C0029423|T191|MH|D015831|MSH|Osteochondroma|9210/0
C0029423|T191|PM|D015831|MSH|Osteochondromas|9210/0
C0029423|T191|PN|NOCODE|MTH|Cartilaginous exostosis|9210/0
C0029423|T191|SY|C3295|NCI|Osteocartilaginous Exostosis|9210/0
C0029423|T191|PT|C3295|NCI|Osteochondroma|9210/0
C0029423|T191|PT|C3295|NCI_CDISC|OSTEOCHONDROMA, BENIGN|9210/0
C0029423|T191|PT|XaB9w|RCD|Chondroma of bone|9210/0
C0029423|T191|SY|BBW0.|RCD|Ecchondroma|9210/0
C0029423|T191|SY|BBW0.|RCD|Osteocartilaginous exostosis|9210/0
C0029423|T191|PT|BBW0.|RCD|Osteochondroma|9210/0
C0029423|T191|SY|52299001|SNOMEDCT_US|Cartilaginous exostosis|9210/0
C0029423|T191|PT|307573009|SNOMEDCT_US|Chondroma of bone|9210/0
C0029423|T191|SY|52299001|SNOMEDCT_US|Ecchondroma|9210/0
C0029423|T191|SY|52299001|SNOMEDCT_US|Osteocartilaginous exostosis|9210/0
C0029423|T191|PT|52299001|SNOMEDCT_US|Osteochondroma|9210/0
C0029423|T191|PT|443093007|SNOMEDCT_US|Osteochondroma|9210/0
C0206641|T191|PT|0000020989|CHV|osteochondromatosis|9210/1
C0206641|T191|PT|NOCODE|COSTAR|Osteochondromatosis|9210/1
C0206641|T191|PT|MTHU024639|ICPC2ICD10ENG|ecchondrosis|9210/1
C0206641|T191|PT|MTHU056140|ICPC2ICD10ENG|osteochondromatosis|9210/1
C0206641|T191|PM|D018216|MSH|Osteochondromatoses|9210/1
C0206641|T191|MH|D018216|MSH|Osteochondromatosis|9210/1
C0206641|T191|PN|NOCODE|MTH|Osteochondromatosis|9210/1
C0206641|T191|PT|C53457|NCI|Multiple Osteochondromas|9210/1
C0206641|T191|SY|C53457|NCI|Osteochondromatosis|9210/1
C0206641|T191|SY|CDR0000654671|PDQ|Multiple Osteochondromas|9210/1
C0206641|T191|PT|CDR0000654671|PDQ|osteochondromatosis|9210/1
C0206641|T191|SY|Xa9AX|RCD|Ecchondrosis|9210/1
C0206641|T191|PT|Xa9AX|RCD|Osteochondromatosis|9210/1
C0206641|T191|OP|BBW1.|RCDSY|Osteochondromatosis NOS|9210/1
C0206641|T191|OAS|302860009|SNOMEDCT_US|Ecchondrosis|9210/1
C0206641|T191|SY|66467005|SNOMEDCT_US|Ecchondrosis|9210/1
C0206641|T191|OAP|302860009|SNOMEDCT_US|Osteochondromatosis|9210/1
C0206641|T191|PT|66467005|SNOMEDCT_US|Osteochondromatosis|9210/1
C0206641|T191|IS|66467005|SNOMEDCT_US|Osteochondromatosis, NOS|9210/1
C3839106|T191|PT|C121842|NCI|Osteochondromyxoma|9211/0
C3839106|T191|PT|703695006|SNOMEDCT_US|Osteochondromyxoma|9211/0
C2960319|T191|PT|355233|MEDCIN|Bizarre parosteal osteochondromatous proliferation|9212/0
C2960319|T191|PT|C121845|NCI|Bizarre Parosteal Osteochondromatous Proliferation|9212/0
C2960319|T191|AB|C121845|NCI|BPOP|9212/0
C2960319|T191|SY|C121845|NCI|Nora's Lesion|9212/0
C2960319|T191|PT|703696007|SNOMEDCT_US|Bizarre parosteal osteochondromatous proliferation|9212/0
C2960319|T191|PT|446593006|SNOMEDCT_US|Bizarre parosteal osteochondromatous proliferation|9212/0
C2960319|T191|SY|446593006|SNOMEDCT_US|Nora lesion|9212/0
C0038604|T191|NM|C535723|MSH|Subungual exostoses|9213/0
C0038604|T191|SY|C121844|NCI|Dupuytren Exostosis|9213/0
C0038604|T191|PT|C121844|NCI|Subungual Exostosis|9213/0
C0038604|T191|PT|X50Fw|RCD|Subungual exostosis|9213/0
C0038604|T191|OAP|202895008|SNOMEDCT_US|Subungual exostosis|9213/0
C0038604|T191|OF|202895008|SNOMEDCT_US|Subungual exostosis|9213/0
C0038604|T191|PT|703697003|SNOMEDCT_US|Subungual exostosis|9213/0
C0038604|T191|PT|26904005|SNOMEDCT_US|Subungual exostosis|9213/0
C0936248|T191|ET|0000004539|AOD|chondroma|9220/0
C0936248|T191|SY|0000052862|CHV|chondroma|9220/0
C0936248|T191|SY|0000052862|CHV|chondromas|9220/0
C1704356|T191|PT|0000004432|CHV|enchondroma|9220/0
C1704356|T191|PT|0000052862|CHV|enchondroma|9220/0
C1704356|T191|SY|0000004432|CHV|enchondromas|9220/0
C0936248|T191|PT|NOCODE|COSTAR|Chondroma|9220/0
C1704356|T191|PT|NOCODE|COSTAR|Enchondroma|9220/0
C1704356|T191|PT|HP:0030038|HPO|Enchondroma|9220/0
C1704356|T191|PT|U005372|LCH|Enchondroma|9220/0
C1704356|T191|PT|sh85042985|LCH_NW|Enchondroma|9220/0
C0936248|T191|LLT|10008725|MDR|Chondroma|9220/0
C0936248|T191|PT|10008725|MDR|Chondroma|9220/0
C1704356|T191|LLT|10069069|MDR|Enchondroma|9220/0
C0936248|T191|MH|D002812|MSH|Chondroma|9220/0
C0936248|T191|PM|D002812|MSH|Chondromas|9220/0
C1704356|T191|PEP|D002812|MSH|Enchondroma|9220/0
C1704356|T191|PM|D002812|MSH|Enchondromas|9220/0
C0936248|T191|PN|NOCODE|MTH|Chondroma|9220/0
C1704356|T191|PN|NOCODE|MTH|Enchondroma|9220/0
C1704356|T191|SY|C3007|NCI|Central Chondroma|9220/0
C0936248|T191|PT|C53459|NCI|Chondroma|9220/0
C1704356|T191|PT|C3007|NCI|Enchondroma|9220/0
C0936248|T191|PT|C53459|NCI_CDISC|CHONDROMA, BENIGN|9220/0
C1704356|T191|PT|CDR0000044252|NCI_NCI-GLOSS|enchondroma|9220/0
C0936248|T191|PT|Xa9AY|RCD|Chondroma|9220/0
C1704356|T191|SY|Xa9AY|RCD|Enchondroma|9220/0
C0936248|T191|OP|BBW2.|RCDSY|Chondroma NOS|9220/0
C0936248|T191|OAS|269638002|SNOMEDCT_US|Chondroma|9220/0
C0936248|T191|OAS|188980001|SNOMEDCT_US|Chondroma|9220/0
C0936248|T191|PT|31186001|SNOMEDCT_US|Chondroma|9220/0
C0936248|T191|OAS|187899007|SNOMEDCT_US|Chondroma|9220/0
C0936248|T191|OAS|154611005|SNOMEDCT_US|Chondroma|9220/0
C0936248|T191|IS|31186001|SNOMEDCT_US|Chondroma, NOS|9220/0
C1704356|T191|PT|423699002|SNOMEDCT_US|Enchondroma|9220/0
C1704356|T191|SY|31186001|SNOMEDCT_US|Enchondroma|9220/0
C1704356|T191|SY|423699002|SNOMEDCT_US|True chondroma|9220/0
C0206636|T191|PT|0000020985|CHV|chondromatosis|9220/1
C0008476|T191|PT|0000002903|CHV|synovial chondromatosis|9220/1
C0008476|T191|SY|0000002903|CHV|synovial chondrometaplasia|9220/1
C0206636|T191|PTN|L71016|ICPC2P|chondromatosis|9220/1
C0206636|T191|PT|L71016|ICPC2P|Chondromatosis|9220/1
C0206636|T191|LLT|10051503|MDR|Chondromatosis|9220/1
C0206636|T191|PT|10051503|MDR|Chondromatosis|9220/1
C0008476|T191|LLT|10051522|MDR|Synovial chondromatosis|9220/1
C0008476|T191|SY|31579|MEDCIN|synovial chondromatosis|9220/1
C0008476|T191|PT|31579|MEDCIN|synovial chondromatosis of joint|9220/1
C0206636|T191|PM|D018210|MSH|Chondromatoses|9220/1
C0008476|T191|PM|D015838|MSH|Chondromatoses, Synovial|9220/1
C0206636|T191|MH|D018210|MSH|Chondromatosis|9220/1
C0008476|T191|MH|D015838|MSH|Chondromatosis, Synovial|9220/1
C0008476|T191|PM|D015838|MSH|Chondrometaplasia, Synovial|9220/1
C0008476|T191|PM|D015838|MSH|Chondrometaplasias, Synovial|9220/1
C0008476|T191|PM|D015838|MSH|Henderson Jones Syndrome|9220/1
C0008476|T191|ET|D015838|MSH|Henderson-Jones Syndrome|9220/1
C0008476|T191|PM|D015838|MSH|Reichel Syndrome|9220/1
C0008476|T191|ET|D015838|MSH|Reichel's Syndrome|9220/1
C0008476|T191|PM|D015838|MSH|Reichels Syndrome|9220/1
C0008476|T191|PM|D015838|MSH|Syndrome, Henderson-Jones|9220/1
C0008476|T191|PM|D015838|MSH|Syndrome, Reichel's|9220/1
C0008476|T191|PM|D015838|MSH|Synovial Chondromatoses|9220/1
C0008476|T191|ET|D015838|MSH|Synovial Chondromatosis|9220/1
C0008476|T191|ET|D015838|MSH|Synovial Chondrometaplasia|9220/1
C0008476|T191|PM|D015838|MSH|Synovial Chondrometaplasias|9220/1
C0008476|T191|PN|NOCODE|MTH|Chondromatosis, Synovial|9220/1
C0206636|T191|PT|C35259|NCI|Chondromatosis|9220/1
C0008476|T191|SY|C34467|NCI|Henderson-Jones Syndrome|9220/1
C0008476|T191|SY|C34467|NCI|Reichel's Syndrome|9220/1
C0008476|T191|PT|C34467|NCI|Synovial Chondromatosis|9220/1
C0206636|T191|PT|Xa9AZ|RCD|Chondromatosis|9220/1
C0008476|T191|PT|X70CY|RCD|Synovial chondromatosis|9220/1
C0206636|T191|OP|BBW3.|RCDSY|Chondromatosis NOS|9220/1
C0206636|T191|SY|83944004|SNOMEDCT_US|Cartilage analog of fibromatosis|9220/1
C0206636|T191|SYGB|83944004|SNOMEDCT_US|Cartilage analogue of fibromatosis|9220/1
C0206636|T191|PT|302861008|SNOMEDCT_US|Chondromatosis|9220/1
C0206636|T191|PT|83944004|SNOMEDCT_US|Chondromatosis|9220/1
C0206636|T191|IS|83944004|SNOMEDCT_US|Chondromatosis, NOS|9220/1
C0008476|T191|PT|133850008|SNOMEDCT_US|Primary synovial chondromatosis|9220/1
C0008476|T191|SY|133850008|SNOMEDCT_US|Synovial chondromatosis|9220/1
C0008476|T191|SY|66467005|SNOMEDCT_US|Synovial chondromatosis|9220/1
C0008476|T191|PT|240207006|SNOMEDCT_US|Synovial chondromatosis|9220/1
C0008479|T191|PT|0000002904|CHV|chondrosarcoma|9220/3
C0008479|T191|SY|0000002904|CHV|chondrosarcomas|9220/3
C0008479|T191|DI|U000341|DXP|CHONDROSARCOMA|9220/3
C0008479|T191|PT|HP:0006765|HPO|Chondrosarcoma|9220/3
C0008479|T191|LLT|10008726|MDR|Chondroma sarcomatosum|9220/3
C0008479|T191|LLT|10008734|MDR|Chondrosarcoma|9220/3
C0008479|T191|PT|10008734|MDR|Chondrosarcoma|9220/3
C0008479|T191|LLT|10008737|MDR|Chondrosarcoma NOS|9220/3
C0008479|T191|PT|355170|MEDCIN|chondrosarcoma|9220/3
C0008479|T191|SY|355170|MEDCIN|malignant neoplasm chondrosarcoma|9220/3
C0008479|T191|MH|D002813|MSH|Chondrosarcoma|9220/3
C0008479|T191|PM|D002813|MSH|Chondrosarcomas|9220/3
C0008479|T191|PN|NOCODE|MTH|Chondrosarcoma|9220/3
C0008479|T191|PT|C2946|NCI|Chondrosarcoma|9220/3
C0008479|T191|PT|C2946|NCI_CDISC|CHONDROSARCOMA, MALIGNANT|9220/3
C0008479|T191|PT|C2946|NCI_CPTAC|Chondrosarcoma|9220/3
C0008479|T191|PT|10008737|NCI_CTEP-SDC|Chondrosarcoma|9220/3
C0008479|T191|PT|C2946|NCI_CTRP|Chondrosarcoma|9220/3
C0008479|T191|DN|C2946|NCI_CTRP|Chondrosarcoma|9220/3
C0008479|T191|PT|CDR0000045221|NCI_NCI-GLOSS|chondrosarcoma|9220/3
C0008479|T191|PSC|CDR0000039486|PDQ|chondrosarcoma|9220/3
C0008479|T191|ET|CDR0000039486|PDQ|Chondrosarcoma|9220/3
C0008479|T191|PT|XaB9x|RCD|Chondrosarcoma morphology|9220/3
C0008479|T191|OP|BBW4.|RCDSY|Chondrosarcoma NOS|9220/3
C0008479|T191|PT|443520009|SNOMEDCT_US|Chondrosarcoma|9220/3
C0008479|T191|SY|14990007|SNOMEDCT_US|Chondrosarcoma|9220/3
C0008479|T191|SY|14990007|SNOMEDCT_US|Chondrosarcoma morphology|9220/3
C3838951|T191|PT|703699000|SNOMEDCT_US|Chondrosarcoma, grade 2|9220/3
C3838808|T191|PT|703700004|SNOMEDCT_US|Chondrosarcoma, grade 3|9220/3
C0008479|T191|PT|14990007|SNOMEDCT_US|Chondrosarcoma, no ICD-O subtype|9220/3
C0008479|T191|SY|14990007|SNOMEDCT_US|Chondrosarcoma, no International Classification of Diseases for Oncology subtype|9220/3
C0008479|T191|IS|14990007|SNOMEDCT_US|Chondrosarcoma, NOS|9220/3
C0008479|T191|SY|443520009|SNOMEDCT_US|Fibrochondrosarcoma|9220/3
C0334548|T191|SY|0000030004|CHV|juxtacortical chondroma|9221/0
C0334548|T191|PT|0000030004|CHV|periosteal chondroma|9221/0
C0334548|T191|SY|C4302|NCI|Juxtacortical Chondroma|9221/0
C0334548|T191|PT|C4302|NCI|Periosteal Chondroma|9221/0
C0334548|T191|PT|BBW5.|RCD|Juxtacortical chondroma|9221/0
C0334548|T191|SY|BBW5.|RCD|Periosteal chondroma|9221/0
C0334548|T191|PT|9266000|SNOMEDCT_US|Juxtacortical chondroma|9221/0
C0334548|T191|SY|9266000|SNOMEDCT_US|Periosteal chondroma|9221/0
C0334549|T191|SY|C7357|NCI|Juxtacortical Chondrosarcoma|9221/3
C0334549|T191|PT|C7357|NCI|Periosteal Chondrosarcoma|9221/3
C0334549|T191|PT|BBW6.|RCD|Juxtacortical chondrosarcoma|9221/3
C0334549|T191|PT|26211003|SNOMEDCT_US|Juxtacortical chondrosarcoma|9221/3
C0334549|T191|SY|26211003|SNOMEDCT_US|Periosteal chondrosarcoma|9221/3
C3838825|T191|PT|703701000|SNOMEDCT_US|Atypical cartilaginous tumor|9222/1
C3838825|T191|PTGB|703701000|SNOMEDCT_US|Atypical cartilaginous tumour|9222/1
C3838825|T191|SY|703701000|SNOMEDCT_US|Chondrosarcoma, grade 1|9222/1
C0008441|T191|ET|0000004546|AOD|chondroblastoma|9230/0
C0008441|T191|PT|0000002897|CHV|chondroblastoma|9230/0
C0008441|T191|SY|0000002897|CHV|chondroblastomas|9230/0
C0008441|T191|ET|2019-1220|CSP|chondroblastoma|9230/0
C0008441|T191|PT|HP:0030432|HPO|Chondroblastoma|9230/0
C0008441|T191|PT|U000994|LCH|Chondroblastoma|9230/0
C0008441|T191|PT|sh85024676|LCH_NW|Chondroblastoma|9230/0
C0008441|T191|LLT|10008686|MDR|Chondroblastoma|9230/0
C0008441|T191|PT|10008686|MDR|Chondroblastoma|9230/0
C0008441|T191|MH|D002804|MSH|Chondroblastoma|9230/0
C0008441|T191|PM|D002804|MSH|Chondroblastomas|9230/0
C0008441|T191|PT|C2945|NCI|Chondroblastoma|9230/0
C0008441|T191|SY|Xa9Ab|RCD|Chondroblastoma|9230/0
C0008441|T191|PT|XaB9y|RCD|Chondroblastoma morphology|9230/0
C0008441|T191|PT|Xa9Ab|RCD|Chondroblastoma of bone|9230/0
C0008441|T191|AB|Xa9Ab|RCD|Chondromatous giant cell tum|9230/0
C0008441|T191|SY|Xa9Ab|RCD|Chondromatous giant cell tumour|9230/0
C0008441|T191|SY|Xa9Ab|RCD|Codman's tumour|9230/0
C0008441|T191|SY|Xa9Ab|RCDAE|Chondromatous giant cell tumor|9230/0
C0008441|T191|SY|Xa9Ab|RCDAE|Codman's tumor|9230/0
C0008441|T191|OP|BBW7.|RCDSY|Chondroblastoma NOS|9230/0
C0008441|T191|PT|9001003|SNOMEDCT_US|Chondroblastoma|9230/0
C0008441|T191|SY|9001003|SNOMEDCT_US|Chondroblastoma morphology|9230/0
C0008441|T191|OAP|134337007|SNOMEDCT_US|Chondroblastoma of bone|9230/0
C0008441|T191|OF|134337007|SNOMEDCT_US|Chondroblastoma of bone|9230/0
C0008441|T191|IS|9001003|SNOMEDCT_US|Chondroblastoma, NOS|9230/0
C0008441|T191|SY|9001003|SNOMEDCT_US|Chondromatous giant cell tumor|9230/0
C0008441|T191|SYGB|9001003|SNOMEDCT_US|Chondromatous giant cell tumour|9230/0
C0008441|T191|SY|9001003|SNOMEDCT_US|Codman's tumor|9230/0
C0008441|T191|SYGB|9001003|SNOMEDCT_US|Codman's tumour|9230/0
C0008441|T191|ET|0000004546|AOD|chondroblastoma|9230/1
C0008441|T191|PT|0000002897|CHV|chondroblastoma|9230/1
C0008441|T191|SY|0000002897|CHV|chondroblastomas|9230/1
C0008441|T191|ET|2019-1220|CSP|chondroblastoma|9230/1
C0008441|T191|PT|HP:0030432|HPO|Chondroblastoma|9230/1
C0008441|T191|PT|U000994|LCH|Chondroblastoma|9230/1
C0008441|T191|PT|sh85024676|LCH_NW|Chondroblastoma|9230/1
C0008441|T191|LLT|10008686|MDR|Chondroblastoma|9230/1
C0008441|T191|PT|10008686|MDR|Chondroblastoma|9230/1
C0008441|T191|MH|D002804|MSH|Chondroblastoma|9230/1
C0008441|T191|PM|D002804|MSH|Chondroblastomas|9230/1
C0008441|T191|PT|C2945|NCI|Chondroblastoma|9230/1
C0008441|T191|SY|Xa9Ab|RCD|Chondroblastoma|9230/1
C0008441|T191|PT|XaB9y|RCD|Chondroblastoma morphology|9230/1
C0008441|T191|PT|Xa9Ab|RCD|Chondroblastoma of bone|9230/1
C0008441|T191|AB|Xa9Ab|RCD|Chondromatous giant cell tum|9230/1
C0008441|T191|SY|Xa9Ab|RCD|Chondromatous giant cell tumour|9230/1
C0008441|T191|SY|Xa9Ab|RCD|Codman's tumour|9230/1
C0008441|T191|SY|Xa9Ab|RCDAE|Chondromatous giant cell tumor|9230/1
C0008441|T191|SY|Xa9Ab|RCDAE|Codman's tumor|9230/1
C0008441|T191|OP|BBW7.|RCDSY|Chondroblastoma NOS|9230/1
C0008441|T191|PT|9001003|SNOMEDCT_US|Chondroblastoma|9230/1
C0008441|T191|SY|9001003|SNOMEDCT_US|Chondroblastoma morphology|9230/1
C0008441|T191|OAP|134337007|SNOMEDCT_US|Chondroblastoma of bone|9230/1
C0008441|T191|OF|134337007|SNOMEDCT_US|Chondroblastoma of bone|9230/1
C0008441|T191|IS|9001003|SNOMEDCT_US|Chondroblastoma, NOS|9230/1
C0008441|T191|SY|9001003|SNOMEDCT_US|Chondromatous giant cell tumor|9230/1
C0008441|T191|SYGB|9001003|SNOMEDCT_US|Chondromatous giant cell tumour|9230/1
C0008441|T191|SY|9001003|SNOMEDCT_US|Codman's tumor|9230/1
C0008441|T191|SYGB|9001003|SNOMEDCT_US|Codman's tumour|9230/1
C4054527|T191|PT|C66799|NCI|Metastasizing Chondroblastoma|9230/3
C0334550|T191|PT|BBW8.|RCD|Malignant chondroblastoma|9230/3
C0334550|T191|PT|74279005|SNOMEDCT_US|Chondroblastoma, malignant|9230/3
C0334550|T191|SY|74279005|SNOMEDCT_US|Malignant chondroblastoma|9230/3
C0334551|T191|PT|0000030005|CHV|myxoid chondrosarcoma|9231/3
C0334551|T191|PT|C4303|NCI|Myxoid Chondrosarcoma|9231/3
C0334551|T191|PT|X77pB|RCD|Myxoid chondrosarcoma|9231/3
C0334551|T191|OP|BBV9.|RCDSY|Myxoid chondrosarcoma|9231/3
C0334551|T191|PT|75622000|SNOMEDCT_US|Myxoid chondrosarcoma|9231/3
C0206637|T191|PT|0014549|CCPSS|CHONDROSARCOMA MESENCHYMAL|9240/3
C0206637|T191|SY|0000020986|CHV|chondrosarcoma mesenchymal|9240/3
C0206637|T191|PT|0000020986|CHV|mesenchymal chondrosarcoma|9240/3
C0206637|T191|LLT|10027389|MDR|Mesenchymal chondrosarcoma|9240/3
C0206637|T191|MH|D018211|MSH|Chondrosarcoma, Mesenchymal|9240/3
C0206637|T191|PM|D018211|MSH|Chondrosarcomas, Mesenchymal|9240/3
C0206637|T191|PM|D018211|MSH|Mesenchymal Chondrosarcoma|9240/3
C0206637|T191|PM|D018211|MSH|Mesenchymal Chondrosarcomas|9240/3
C0206637|T191|PN|NOCODE|MTH|Mesenchymal Chondrosarcoma|9240/3
C0206637|T191|PT|C3737|NCI|Mesenchymal Chondrosarcoma|9240/3
C0206637|T191|PT|BBW9.|RCD|Mesenchymal chondrosarcoma|9240/3
C0206637|T191|PT|56565002|SNOMEDCT_US|Mesenchymal chondrosarcoma|9240/3
C0221290|T191|DI|U000647|DXP|FIBROMA, CHONDROMYXOID|9241/0
C0221290|T191|LLT|10008733|MDR|Chondromyxoid fibroma|9241/0
C0221290|T191|PT|C3830|NCI|Chondromyxoid Fibroma|9241/0
C0221290|T191|PT|BBWA.|RCD|Chondromyxoid fibroma|9241/0
C0221290|T191|SY|BBWA.|RCD|CMF - Chondromyxoid fibroma|9241/0
C0221290|T191|PT|39553005|SNOMEDCT_US|Chondromyxoid fibroma|9241/0
C0221290|T191|SY|39553005|SNOMEDCT_US|CMF - Chondromyxoid fibroma|9241/0
C1266167|T191|MH|D000077207|MSH|Chondrosarcoma, Clear Cell|9242/3
C1266167|T191|PM|D000077207|MSH|Chondrosarcomas, Clear Cell|9242/3
C1266167|T191|ET|D000077207|MSH|Clear Cell Chondrosarcoma|9242/3
C1266167|T191|PM|D000077207|MSH|Clear Cell Chondrosarcomas|9242/3
C1266167|T191|PT|C6475|NCI|Clear Cell Chondrosarcoma|9242/3
C1266167|T191|PT|128775007|SNOMEDCT_US|Clear cell chondrosarcoma|9242/3
C0862878|T191|LLT|10011986|MDR|Dedifferentiated chondrosarcoma|9243/3
C0862878|T191|PT|C6476|NCI|Dedifferentiated Chondrosarcoma|9243/3
C0862878|T191|PT|128776008|SNOMEDCT_US|Dedifferentiated chondrosarcoma|9243/3
C0206638|T191|SY|0000020987|CHV|bone cell giant tumor|9250/1
C0206638|T191|SY|0000020987|CHV|bone cell giant tumours|9250/1
C0206638|T191|SY|0000020987|CHV|giant cell bone tumor|9250/1
C0206638|T191|SY|0000020987|CHV|giant cell tumor bone|9250/1
C0206638|T191|SY|0000020987|CHV|giant cell tumor of bone|9250/1
C0206638|T191|PT|0000020987|CHV|osteoclastoma|9250/1
C0206638|T191|SY|0000020987|CHV|osteoclastomas|9250/1
C0206638|T191|PT|U000027|COSTAR|GIANT CELL TUMOR OF BONE|9250/1
C0206638|T191|DI|U000228|DXP|BONE, GIANT CELL TUMOR|9250/1
C0206638|T191|SY|NOCODE|DXP|OSTEOCLASTOMA|9250/1
C0206638|T191|PT|HP:0011847|HPO|Giant cell tumor of bone|9250/1
C0206638|T191|PT|MTHU064709|ICPC2ICD10ENG|giant cell; tumor, bone|9250/1
C0206638|T191|PT|MTHU056233|ICPC2ICD10ENG|osteoclastoma|9250/1
C0206638|T191|PT|MTHU077146|ICPC2ICD10ENG|tumor; giant cell, bone|9250/1
C0206638|T191|LLT|10062381|MDR|Benign bone giant cell tumor|9250/1
C0206638|T191|LLT|10004239|MDR|Benign bone giant cell tumour|9250/1
C0206638|T191|LLT|10005968|MDR|Bone giant cell tumor|9250/1
C0206638|T191|MTH_PT|10005969|MDR|Bone giant cell tumor|9250/1
C0206638|T191|LLT|10062385|MDR|Bone giant cell tumor benign|9250/1
C0206638|T191|MTH_PT|10005970|MDR|Bone giant cell tumor benign|9250/1
C0206638|T191|LLT|10005969|MDR|Bone giant cell tumour|9250/1
C0206638|T191|PT|10005969|MDR|Bone giant cell tumour|9250/1
C0206638|T191|LLT|10005970|MDR|Bone giant cell tumour benign|9250/1
C0206638|T191|PT|10005970|MDR|Bone giant cell tumour benign|9250/1
C0206638|T191|PT|31492|MEDCIN|benign giant cell tumor of bone|9250/1
C0206638|T191|SY|31492|MEDCIN|benign giant-cell tumor in the bone|9250/1
C0206638|T191|MH|D018212|MSH|Giant Cell Tumor of Bone|9250/1
C0206638|T191|PN|NOCODE|MTH|Giant Cell Tumor of Bone|9250/1
C0206638|T191|PT|C121932|NCI|Giant Cell Tumor of Bone|9250/1
C0206638|T191|SY|C121932|NCI|Giant Cell Tumor of the Bone|9250/1
C4048303|T191|PT|C3738|NCI|Osteoclastic Giant Cell-Rich Tumor of Bone|9250/1
C4048303|T191|SY|C3738|NCI|Osteoclastic Giant Cell-Rich Tumor of the Bone|9250/1
C0206638|T191|SY|C121932|NCI|Osteoclastoma|9250/1
C0206638|T191|SY|C121932|NCI_CDISC|Benign Bone Giant Cell Tumor|9250/1
C0206638|T191|PT|C121932|NCI_CDISC|GIANT CELL TUMOR, BENIGN|9250/1
C0206638|T191|SY|C121932|NCI_CDISC|Osteoclastoma, Benign|9250/1
C0206638|T191|PT|CDR0000530111|PDQ|benign giant cell tumor of bone|9250/1
C0206638|T191|PT|Xa9Ac|RCD|Giant cell tumour of bone|9250/1
C0206638|T191|SY|Xa9Ac|RCD|Osteoclastoma|9250/1
C0206638|T191|PT|Xa9Ac|RCDAE|Giant cell tumor of bone|9250/1
C0206638|T191|OA|BBX0.|RCDSA|Giant cell bone tumor NOS|9250/1
C0206638|T191|OP|BBX0.|RCDSA|Giant cell tumor of bone NOS|9250/1
C0206638|T191|OA|BBX0.|RCDSY|Giant cell bone tumour NOS|9250/1
C0206638|T191|OP|BBX0.|RCDSY|Giant cell tumour of bone NOS|9250/1
C0206638|T191|PT|57500000|SNOMEDCT_US|Giant cell tumor of bone|9250/1
C0206638|T191|PT|697970009|SNOMEDCT_US|Giant cell tumor of bone|9250/1
C0206638|T191|IS|57500000|SNOMEDCT_US|Giant cell tumor of bone, NOS|9250/1
C0206638|T191|PTGB|697970009|SNOMEDCT_US|Giant cell tumour of bone|9250/1
C0206638|T191|PTGB|57500000|SNOMEDCT_US|Giant cell tumour of bone|9250/1
C0206638|T191|SY|697970009|SNOMEDCT_US|GTCT - Giant cell tumor of bone|9250/1
C0206638|T191|SY|57500000|SNOMEDCT_US|Osteoclastoma|9250/1
C0206638|T191|IS|57500000|SNOMEDCT_US|Osteoclastoma, NOS|9250/1
C0334552|T191|LLT|10073108|MDR|Bone giant cell tumor malignant|9250/3
C0334552|T191|MTH_PT|10073106|MDR|Bone giant cell tumor malignant|9250/3
C0334552|T191|LLT|10073106|MDR|Bone giant cell tumour malignant|9250/3
C0334552|T191|PT|10073106|MDR|Bone giant cell tumour malignant|9250/3
C0334552|T191|PT|230755|MEDCIN|giant cell sarcoma of bone|9250/3
C0334552|T191|PN|NOCODE|MTH|Malignant Giant Cell Tumor of Bone|9250/3
C0334552|T191|SY|C4304|NCI|Dedifferentiated Giant Cell Tumor|9250/3
C0334552|T191|SY|C4304|NCI|Giant Cell Bone Sarcoma|9250/3
C0334552|T191|SY|C4304|NCI|Giant Cell Sarcoma of Bone|9250/3
C0334552|T191|SY|C4304|NCI|Giant Cell Sarcoma of the Bone|9250/3
C0334552|T191|PT|C4304|NCI|Malignancy in Giant Cell Tumor of Bone|9250/3
C0334552|T191|SY|C4304|NCI|Malignancy in Giant Cell Tumor of the Bone|9250/3
C0334552|T191|SY|C4304|NCI|Malignant Giant Cell Tumor of Bone|9250/3
C0334552|T191|SY|C4304|NCI_CDISC|Dedifferentiated Giant Cell Tumor|9250/3
C0334552|T191|SY|C4304|NCI_CDISC|Giant Cell Bone Sarcoma|9250/3
C0334552|T191|SY|C4304|NCI_CDISC|Giant Cell Sarcoma of Bone|9250/3
C0334552|T191|SY|C4304|NCI_CDISC|Giant Cell Sarcoma of the Bone|9250/3
C0334552|T191|PT|C4304|NCI_CDISC|OSTEOCLASTOMA, MALIGNANT|9250/3
C0334552|T191|DN|C4304|NCI_CTRP|Malignancy in Giant Cell Tumor of Bone|9250/3
C0334552|T191|PT|CDR0000530113|PDQ|malignant giant cell tumor of bone|9250/3
C0334552|T191|SY|BBX1.|RCD|Giant cell sarcoma of bone|9250/3
C0334552|T191|AB|BBX1.|RCD|Malig giant cell tum of bone|9250/3
C0334552|T191|PT|BBX1.|RCD|Malignant giant cell tumour of bone|9250/3
C0334552|T191|SY|BBX1.|RCD|Malignant osteoclastoma|9250/3
C0334552|T191|PT|BBX1.|RCDAE|Malignant giant cell tumor of bone|9250/3
C0334552|T191|SY|10069009|SNOMEDCT_US|Giant cell sarcoma of bone|9250/3
C0334552|T191|PT|10069009|SNOMEDCT_US|Giant cell tumor of bone, malignant|9250/3
C0334552|T191|PTGB|10069009|SNOMEDCT_US|Giant cell tumour of bone, malignant|9250/3
C0334552|T191|SY|10069009|SNOMEDCT_US|Malignant giant cell tumor of bone|9250/3
C0334552|T191|SYGB|10069009|SNOMEDCT_US|Malignant giant cell tumour of bone|9250/3
C0334552|T191|SY|10069009|SNOMEDCT_US|Malignant osteoclastoma|9250/3
C0334552|T191|SY|10069009|SNOMEDCT_US|Osteoclastoma, malignant|9250/3
C0039106|T191|SY|0000057940|CHV|pigmented synovitis villonodular|9251/0
C0039106|T191|SY|0000011984|CHV|pigmented synovitis villonodular|9251/0
C0039106|T191|PT|0000057940|CHV|pigmented villonodular synovitis|9251/0
C0039106|T191|PT|0000011984|CHV|pigmented villonodular synovitis|9251/0
C0039106|T191|SY|0000057940|CHV|villonodular synovitis|9251/0
C0039106|T191|DI|U001802|DXP|SYNOVITIS, VILLONODULAR, PIGMENTED|9251/0
C0039106|T191|PT|MTHU073148|ICPC2ICD10ENG|synovitis; villonodular|9251/0
C0039106|T191|PT|MTHU080787|ICPC2ICD10ENG|villonodular; synovitis|9251/0
C0039106|T191|PT|32592|MEDCIN|pigmented villonodular synovitis|9251/0
C0039106|T191|ET|D013586|MSH|Diffuse Tenosynovial Giant Cell Tumor|9251/0
C0039106|T191|PM|D013586|MSH|Pigmented Villonodular Synovitides|9251/0
C0039106|T191|PM|D013586|MSH|Pigmented Villonodular Synovitis|9251/0
C0039106|T191|PM|D013586|MSH|Synovitides, Pigmented Villonodular|9251/0
C0039106|T191|MH|D013586|MSH|Synovitis, Pigmented Villonodular|9251/0
C0039106|T191|PM|D013586|MSH|Villonodular Synovitides, Pigmented|9251/0
C0039106|T191|PM|D013586|MSH|Villonodular Synovitis, Pigmented|9251/0
C0039106|T191|PN|NOCODE|MTH|Pigmented villonodular synovitis|9251/0
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Neoplasm of Tendon Sheath|9251/0
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Neoplasm of Tenosynovium|9251/0
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Neoplasm of the Tenosynovium|9251/0
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Tumor of Tendon Sheath|9251/0
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Tumor of Tenosynovium|9251/0
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Tumor of the Tenosynovium|9251/0
C0039106|T191|SY|C3401|NCI|Diffuse Tenosynovial Giant Cell Neoplasm|9251/0
C0039106|T191|SY|C3401|NCI|Diffuse Tenosynovial Giant Cell Tumor|9251/0
C0039106|T191|SY|C3401|NCI|Pigmented Villonodular Synovitis|9251/0
C0039106|T191|PT|C3401|NCI|Tenosynovial Giant Cell Tumor, Diffuse Type|9251/0
C0039106|T191|AB|N092.|RCD|Pigmented villonod synovitis|9251/0
C0039106|T191|PT|N092.|RCD|Pigmented villonodular synovitis|9251/0
C0039106|T191|SY|N092.|RCD|PVNS - Pigmented villonodular synovitis|9251/0
C0039106|T191|AB|N092.|RCD|PVNS-Pigmen villonod synovitis|9251/0
C0039106|T191|SYGB|95412009|SNOMEDCT_US|Chronic haemorrhagic villous synovitis|9251/0
C0039106|T191|SY|95412009|SNOMEDCT_US|Chronic hemorrhagic villous synovitis|9251/0
C0039106|T191|IS|71508003|SNOMEDCT_US|Pigmented villonodular synovitis|9251/0
C0039106|T191|OAP|202903009|SNOMEDCT_US|Pigmented villonodular synovitis|9251/0
C0039106|T191|OF|202903009|SNOMEDCT_US|Pigmented villonodular synovitis|9251/0
C0039106|T191|SY|703703002|SNOMEDCT_US|Pigmented villonodular synovitis|9251/0
C0039106|T191|PT|95412009|SNOMEDCT_US|Pigmented villonodular synovitis|9251/0
C0039106|T191|SY|95412009|SNOMEDCT_US|PVNS - Pigmented villonodular synovitis|9251/0
C0039106|T191|PT|703703002|SNOMEDCT_US|Tenosynovial giant cell tumor, diffuse|9251/0
C0039106|T191|PTGB|703703002|SNOMEDCT_US|Tenosynovial giant cell tumour, diffuse|9251/0
C0039106|T191|IS|95412009|SNOMEDCT_US|Villonodular synovitis|9251/0
C0039106|T191|IS|95412009|SNOMEDCT_US|Villous tenosynovitis|9251/0
C0039106|T191|IS|71508003|SNOMEDCT_US|Villous tenosynovitis|9251/0
C0334553|T191|PT|231999|MEDCIN|giant cell tumor of soft tissue|9251/1
C0334553|T191|PN|NOCODE|MTH|Giant Cell Tumor of Soft Tissue|9251/1
C0334553|T191|AB|C49107|NCI|GCT-ST|9251/1
C0334553|T191|PT|C49107|NCI|Giant Cell Tumor of Soft Tissue|9251/1
C0334553|T191|SY|C49107|NCI|Osteoclastoma of Soft Tissue|9251/1
C0334553|T191|AB|Xa9Ad|RCD|Giant cell tum of soft tissue|9251/1
C0334553|T191|PT|Xa9Ad|RCD|Giant cell tumour of soft tissue|9251/1
C0334553|T191|PT|Xa9Ad|RCDAE|Giant cell tumor of soft tissue|9251/1
C0334553|T191|OP|BBX2.|RCDSA|Giant cell tumor of soft parts NOS|9251/1
C0334553|T191|OA|BBX2.|RCDSY|Giant cell tum/soft prt NOS|9251/1
C0334553|T191|OP|BBX2.|RCDSY|Giant cell tumour of soft parts NOS|9251/1
C0334553|T191|PT|82125002|SNOMEDCT_US|Giant cell tumor of soft parts|9251/1
C0334553|T191|IS|82125002|SNOMEDCT_US|Giant cell tumor of soft parts, NOS|9251/1
C0334553|T191|SY|82125002|SNOMEDCT_US|Giant cell tumor of soft tissue|9251/1
C0334553|T191|PTGB|82125002|SNOMEDCT_US|Giant cell tumour of soft parts|9251/1
C0334553|T191|SYGB|82125002|SNOMEDCT_US|Giant cell tumour of soft tissue|9251/1
C0334554|T191|LLT|10073141|MDR|Malignant giant cell fibrous histiocytoma|9251/3
C0334554|T191|PT|10073141|MDR|Malignant giant cell fibrous histiocytoma|9251/3
C0334554|T191|PN|NOCODE|MTH|Giant Cell Fibrous Histiocytoma|9251/3
C0334554|T191|OP|C8380|NCI|Giant Cell Fibrous Histiocytoma|9251/3
C0334554|T191|OP|C8380|NCI|Giant Cell Malignant Fibrous Histiocytoma|9251/3
C0334554|T191|OP|C8380|NCI|Malignant Giant Cell Neoplasm of Soft Parts|9251/3
C0334554|T191|OP|C8380|NCI|Malignant Giant Cell Tumor of Soft Parts|9251/3
C0334554|T191|OP|C8380|NCI|Malignant Osteoclastoma|9251/3
C0334554|T191|PT|C8380|NCI|Undifferentiated Pleomorphic Sarcoma with Osteoclast-Like Giant Cells|9251/3
C0334554|T191|AB|BBX3.|RCD|Malig giant cell tum soft tiss|9251/3
C0334554|T191|PT|BBX3.|RCD|Malignant giant cell tumour of soft tissue|9251/3
C0334554|T191|PT|BBX3.|RCDAE|Malignant giant cell tumor of soft tissue|9251/3
C0334554|T191|PT|48460009|SNOMEDCT_US|Malignant giant cell tumor of soft parts|9251/3
C0334554|T191|SY|48460009|SNOMEDCT_US|Malignant giant cell tumor of soft tissue|9251/3
C0334554|T191|PTGB|48460009|SNOMEDCT_US|Malignant giant cell tumour of soft parts|9251/3
C0334554|T191|SYGB|48460009|SNOMEDCT_US|Malignant giant cell tumour of soft tissue|9251/3
C0588125|T191|SY|0000040957|CHV|cell giant sheath tendon tumor|9252/0
C0588125|T191|SY|0000040957|CHV|cell giant sheath tendon tumour|9252/0
C0588125|T191|SY|0000040957|CHV|giant cell tendon sheath tumor|9252/0
C0588125|T191|SY|0000040957|CHV|giant cell tumor tendon sheath|9252/0
C0588125|T191|SY|0000040957|CHV|giant cell tumour tendon sheath|9252/0
C0588125|T191|PT|0000040957|CHV|nodular tenosynovitis|9252/0
C1318543|T191|DI|U001823|DXP|TENDON SHEATH, GIANT CELL TUMOR|9252/0
C1318543|T191|PT|727.02|ICD9CM|Giant cell tumor of tendon sheath|9252/0
C1318543|T191|AB|727.02|ICD9CM|Giant cell tumor tendon|9252/0
C1318543|T191|LLT|10018253|MDR|Giant cell tumor of tendon sheath|9252/0
C1318543|T191|MTH_PT|10018255|MDR|Giant cell tumor of tendon sheath|9252/0
C1318543|T191|LLT|10018255|MDR|Giant cell tumour of tendon sheath|9252/0
C1318543|T191|PT|10018255|MDR|Giant cell tumour of tendon sheath|9252/0
C0588125|T191|LLT|10082904|MDR|Nodular tenosynovitis|9252/0
C1318543|T191|PT|91479|MEDCIN|giant cell tumor of tendon sheath|9252/0
C1318543|T191|ET|D000070779|MSH|Fibrous Histiocytoma of Tendon Sheath|9252/0
C1318543|T191|MH|D000070779|MSH|Giant Cell Tumor of Tendon Sheath|9252/0
C0588125|T191|PEP|D000070779|MSH|Localized Giant Cell Tumor of the Tendon Sheath|9252/0
C0588125|T191|PM|D000070779|MSH|Localized Nodular Tenosynovitides|9252/0
C0588125|T191|ET|D000070779|MSH|Localized Nodular Tenosynovitis|9252/0
C0588125|T191|ET|D000070779|MSH|Localized Pigmented Villonodular Synovitis|9252/0
C0588125|T191|PM|D000070779|MSH|Nodular Tenosynovitides|9252/0
C0588125|T191|PM|D000070779|MSH|Nodular Tenosynovitides, Localized|9252/0
C0588125|T191|ET|D000070779|MSH|Nodular Tenosynovitis|9252/0
C0588125|T191|PM|D000070779|MSH|Nodular Tenosynovitis, Localized|9252/0
C1318543|T191|ET|D000070779|MSH|Tenosynovial Giant Cell Tumor|9252/0
C0588125|T191|PM|D000070779|MSH|Tenosynovitides, Localized Nodular|9252/0
C0588125|T191|PM|D000070779|MSH|Tenosynovitides, Nodular|9252/0
C0588125|T191|PM|D000070779|MSH|Tenosynovitis, Localized Nodular|9252/0
C0588125|T191|PM|D000070779|MSH|Tenosynovitis, Nodular|9252/0
C1318543|T191|PN|NOCODE|MTH|Fibrous histiocytoma of tendon sheath|9252/0
C0588125|T191|PN|NOCODE|MTH|Nodular tenosynovitis|9252/0
C1318543|T191|SY|C3402|NCI|Fibrous Histiocytoma of Tendon Sheath|9252/0
C1318543|T191|SY|C3402|NCI|Giant Cell Neoplasm of Tendon Sheath|9252/0
C1318543|T191|SY|C3402|NCI|Giant Cell Neoplasm of Tenosynovium|9252/0
C1318543|T191|SY|C3402|NCI|Giant Cell Neoplasm of the Tenosynovium|9252/0
C1318543|T191|SY|C3402|NCI|Giant Cell Tumor of Tendon Sheath|9252/0
C1318543|T191|SY|C3402|NCI|Giant Cell Tumor of Tenosynovium|9252/0
C1318543|T191|SY|C3402|NCI|Giant Cell Tumor of the Tenosynovium|9252/0
C0588125|T191|SY|C6532|NCI|Localized Giant Cell Neoplasm of Tendon Sheath|9252/0
C0588125|T191|SY|C6532|NCI|Localized Giant Cell Neoplasm of Tenosynovium|9252/0
C0588125|T191|SY|C6532|NCI|Localized Giant Cell Neoplasm of the Tenosynovium|9252/0
C0588125|T191|SY|C6532|NCI|Localized Giant Cell Tumor of Tendon Sheath|9252/0
C0588125|T191|SY|C6532|NCI|Localized Giant Cell Tumor of Tenosynovium|9252/0
C0588125|T191|SY|C6532|NCI|Localized Giant Cell Tumor of the Tenosynovium|9252/0
C0588125|T191|SY|C6532|NCI|Localized Tenosynovial Giant Cell Neoplasm|9252/0
C0588125|T191|SY|C6532|NCI|Localized Tenosynovial Giant Cell Tumor|9252/0
C0588125|T191|SY|C6532|NCI|Nodular Tenosynovitis|9252/0
C1318543|T191|SY|C3402|NCI|Tendon Sheath Giant Cell Neoplasm|9252/0
C1318543|T191|SY|C3402|NCI|Tendon Sheath Giant Cell Tumor|9252/0
C1318543|T191|SY|C3402|NCI|Tenosynovial Giant Cell Neoplasm|9252/0
C1318543|T191|PT|C3402|NCI|Tenosynovial Giant Cell Tumor|9252/0
C0588125|T191|PT|C6532|NCI|Tenosynovial Giant Cell Tumor, Localized Type|9252/0
C1318543|T191|AB|XaCL4|RCD|Fibr histiocytom tendon sheath|9252/0
C1318543|T191|PT|XaCL4|RCD|Fibrous histiocytoma of tendon sheath|9252/0
C1318543|T191|SY|N092.|RCD|Tendon sheath giant cell tumor|9252/0
C1318543|T191|PT|310605004|SNOMEDCT_US|Fibrous histiocytoma of tendon sheath|9252/0
C1318543|T191|SY|128777004|SNOMEDCT_US|Fibrous histiocytoma of tendon sheath|9252/0
C1318543|T191|SY|95413004|SNOMEDCT_US|Giant cell tumor of tendon sheath|9252/0
C1318543|T191|SY|128777004|SNOMEDCT_US|Giant cell tumor of tendon sheath|9252/0
C1318543|T191|IS|71508003|SNOMEDCT_US|Giant cell tumor of tendon sheath|9252/0
C1318543|T191|SYGB|95413004|SNOMEDCT_US|Giant cell tumour of tendon sheath|9252/0
C1318543|T191|SYGB|128777004|SNOMEDCT_US|Giant cell tumour of tendon sheath|9252/0
C0588125|T191|OAP|71508003|SNOMEDCT_US|Nodular tenosynovitis|9252/0
C0588125|T191|PT|95413004|SNOMEDCT_US|Nodular tenosynovitis|9252/0
C0588125|T191|IS|71508003|SNOMEDCT_US|Nodular tenosynovitis -RETIRED-|9252/0
C0588125|T191|OF|71508003|SNOMEDCT_US|Nodular tenosynovitis -RETIRED-|9252/0
C1318543|T191|IS|95412009|SNOMEDCT_US|Tendon sheath giant cell tumor|9252/0
C1318543|T191|IS|95412009|SNOMEDCT_US|Tendon sheath giant cell tumour|9252/0
C1318543|T191|PT|128777004|SNOMEDCT_US|Tenosynovial giant cell tumor|9252/0
C0588125|T191|PT|703702007|SNOMEDCT_US|Tenosynovial giant cell tumor, localized|9252/0
C1318543|T191|PTGB|128777004|SNOMEDCT_US|Tenosynovial giant cell tumour|9252/0
C0588125|T191|PTGB|703702007|SNOMEDCT_US|Tenosynovial giant cell tumour, localised|9252/0
C0039106|T191|SY|0000057940|CHV|pigmented synovitis villonodular|9252/1
C0039106|T191|SY|0000011984|CHV|pigmented synovitis villonodular|9252/1
C0039106|T191|PT|0000057940|CHV|pigmented villonodular synovitis|9252/1
C0039106|T191|PT|0000011984|CHV|pigmented villonodular synovitis|9252/1
C0039106|T191|SY|0000057940|CHV|villonodular synovitis|9252/1
C0039106|T191|DI|U001802|DXP|SYNOVITIS, VILLONODULAR, PIGMENTED|9252/1
C0039106|T191|PT|MTHU073148|ICPC2ICD10ENG|synovitis; villonodular|9252/1
C0039106|T191|PT|MTHU080787|ICPC2ICD10ENG|villonodular; synovitis|9252/1
C0039106|T191|PT|32592|MEDCIN|pigmented villonodular synovitis|9252/1
C0039106|T191|ET|D013586|MSH|Diffuse Tenosynovial Giant Cell Tumor|9252/1
C0039106|T191|PM|D013586|MSH|Pigmented Villonodular Synovitides|9252/1
C0039106|T191|PM|D013586|MSH|Pigmented Villonodular Synovitis|9252/1
C0039106|T191|PM|D013586|MSH|Synovitides, Pigmented Villonodular|9252/1
C0039106|T191|MH|D013586|MSH|Synovitis, Pigmented Villonodular|9252/1
C0039106|T191|PM|D013586|MSH|Villonodular Synovitides, Pigmented|9252/1
C0039106|T191|PM|D013586|MSH|Villonodular Synovitis, Pigmented|9252/1
C0039106|T191|PN|NOCODE|MTH|Pigmented villonodular synovitis|9252/1
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Neoplasm of Tendon Sheath|9252/1
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Neoplasm of Tenosynovium|9252/1
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Neoplasm of the Tenosynovium|9252/1
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Tumor of Tendon Sheath|9252/1
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Tumor of Tenosynovium|9252/1
C0039106|T191|SY|C3401|NCI|Diffuse Giant Cell Tumor of the Tenosynovium|9252/1
C0039106|T191|SY|C3401|NCI|Diffuse Tenosynovial Giant Cell Neoplasm|9252/1
C0039106|T191|SY|C3401|NCI|Diffuse Tenosynovial Giant Cell Tumor|9252/1
C0039106|T191|SY|C3401|NCI|Pigmented Villonodular Synovitis|9252/1
C0039106|T191|PT|C3401|NCI|Tenosynovial Giant Cell Tumor, Diffuse Type|9252/1
C0039106|T191|AB|N092.|RCD|Pigmented villonod synovitis|9252/1
C0039106|T191|PT|N092.|RCD|Pigmented villonodular synovitis|9252/1
C0039106|T191|SY|N092.|RCD|PVNS - Pigmented villonodular synovitis|9252/1
C0039106|T191|AB|N092.|RCD|PVNS-Pigmen villonod synovitis|9252/1
C0039106|T191|SYGB|95412009|SNOMEDCT_US|Chronic haemorrhagic villous synovitis|9252/1
C0039106|T191|SY|95412009|SNOMEDCT_US|Chronic hemorrhagic villous synovitis|9252/1
C0039106|T191|PT|95412009|SNOMEDCT_US|Pigmented villonodular synovitis|9252/1
C0039106|T191|IS|71508003|SNOMEDCT_US|Pigmented villonodular synovitis|9252/1
C0039106|T191|OAP|202903009|SNOMEDCT_US|Pigmented villonodular synovitis|9252/1
C0039106|T191|OF|202903009|SNOMEDCT_US|Pigmented villonodular synovitis|9252/1
C0039106|T191|SY|703703002|SNOMEDCT_US|Pigmented villonodular synovitis|9252/1
C0039106|T191|SY|95412009|SNOMEDCT_US|PVNS - Pigmented villonodular synovitis|9252/1
C0039106|T191|PT|703703002|SNOMEDCT_US|Tenosynovial giant cell tumor, diffuse|9252/1
C0039106|T191|PTGB|703703002|SNOMEDCT_US|Tenosynovial giant cell tumour, diffuse|9252/1
C0039106|T191|IS|95412009|SNOMEDCT_US|Villonodular synovitis|9252/1
C0039106|T191|IS|95412009|SNOMEDCT_US|Villous tenosynovitis|9252/1
C0039106|T191|IS|71508003|SNOMEDCT_US|Villous tenosynovitis|9252/1
C1266168|T191|SY|C6535|NCI|Malignant Giant Cell Neoplasm of Tendon Sheath|9252/3
C1266168|T191|SY|C6535|NCI|Malignant Giant Cell Neoplasm of the Tendon Sheath|9252/3
C1266168|T191|SY|C6535|NCI|Malignant Giant Cell Tumor of Tendon Sheath|9252/3
C1266168|T191|SY|C6535|NCI|Malignant Giant Cell Tumor of the Tendon Sheath|9252/3
C1266168|T191|SY|C6535|NCI|Malignant Tendon Sheath Giant Cell Neoplasm|9252/3
C1266168|T191|SY|C6535|NCI|Malignant Tendon Sheath Giant Cell Tumor|9252/3
C1266168|T191|PT|C6535|NCI|Malignant Tenosynovial Giant Cell Tumor|9252/3
C1266168|T191|SY|128778009|SNOMEDCT_US|Giant cell tumor of tendon sheath, malignant|9252/3
C1266168|T191|SYGB|128778009|SNOMEDCT_US|Giant cell tumour of tendon sheath, malignant|9252/3
C1266168|T191|PT|128778009|SNOMEDCT_US|Malignant tenosynovial giant cell tumor|9252/3
C1266168|T191|PTGB|128778009|SNOMEDCT_US|Malignant tenosynovial giant cell tumour|9252/3
C0152244|T047|PT|0000017232|CHV|aneurysmal bone cyst|9260/0
C0152244|T047|SY|0000017232|CHV|aneurysmal bone cysts|9260/0
C0152244|T047|SY|0000017232|CHV|bone cyst aneurysmal|9260/0
C0152244|T047|PT|HP:0012063|HPO|Aneurysmal bone cyst|9260/0
C0152244|T047|PT|M85.5|ICD10|Aneurysmal bone cyst|9260/0
C0152244|T047|AB|M85.5|ICD10CM|Aneurysmal bone cyst|9260/0
C0152244|T047|HT|M85.5|ICD10CM|Aneurysmal bone cyst|9260/0
C0152244|T047|AB|M85.50|ICD10CM|Aneurysmal bone cyst, unspecified site|9260/0
C0152244|T047|PT|M85.50|ICD10CM|Aneurysmal bone cyst, unspecified site|9260/0
C0152244|T047|AB|733.22|ICD9CM|Aneurysmal bone cyst|9260/0
C0152244|T047|PT|733.22|ICD9CM|Aneurysmal bone cyst|9260/0
C0152244|T047|PT|MTHU020367|ICPC2ICD10ENG|cyst; bone, aneurysmal|9260/0
C0152244|T047|LLT|10002362|MDR|Aneurysmal bone cyst|9260/0
C0152244|T047|PT|10002362|MDR|Aneurysmal bone cyst|9260/0
C0152244|T047|PT|91784|MEDCIN|aneurysmal bone cyst|9260/0
C0152244|T047|PT|31489|MEDCIN|aneurysmal cyst in bone|9260/0
C0152244|T047|ET|D017824|MSH|Aneurysmal Bone Cysts|9260/0
C0152244|T047|PM|D017824|MSH|Bone Cyst, Aneurysmal|9260/0
C0152244|T047|MH|D017824|MSH|Bone Cysts, Aneurysmal|9260/0
C0152244|T047|PM|D017824|MSH|Cyst, Aneurysmal Bone|9260/0
C0152244|T047|PM|D017824|MSH|Cysts, Aneurysmal Bone|9260/0
C0152244|T047|PN|NOCODE|MTH|Bone Cysts, Aneurysmal|9260/0
C0152244|T047|AB|C3516|NCI|ABC|9260/0
C0152244|T047|PT|C3516|NCI|Aneurysmal Bone Cyst|9260/0
C0152244|T047|SY|C3516|NCI|Aneurysmal Cyst of Bone|9260/0
C0152244|T047|SY|C3516|NCI|Aneurysmal Cyst of the Bone|9260/0
C0152244|T047|SY|N3322|RCD|ABC - Aneurysmal bone cyst|9260/0
C0152244|T047|PT|N3322|RCD|Aneurysmal bone cyst|9260/0
C0152244|T047|SY|203468000|SNOMEDCT_US|ABC - Aneurysmal bone cyst|9260/0
C0152244|T047|PT|203468000|SNOMEDCT_US|Aneurysmal bone cyst|9260/0
C0152244|T047|PT|76000001|SNOMEDCT_US|Aneurysmal bone cyst|9260/0
C0553580|T191|SY|0000039089|CHV|ewing sarcoma|9260/3
C0553580|T191|SY|0000039089|CHV|ewing tumor|9260/3
C0553580|T191|PT|0000039089|CHV|ewing's sarcoma|9260/3
C0553580|T191|SY|0000039089|CHV|ewing's tumor|9260/3
C0553580|T191|SY|0000039089|CHV|ewing's tumors|9260/3
C0553580|T191|SY|0000039089|CHV|ewings sarcoma|9260/3
C0553580|T191|SY|0000039089|CHV|ewings tumor|9260/3
C0553580|T191|SY|0000039089|CHV|ewings tumors|9260/3
C0553580|T191|SY|0000039089|CHV|ewings's sarcoma|9260/3
C0553580|T191|SY|0000039089|CHV|sarcoma ewing|9260/3
C0553580|T191|SY|0000039089|CHV|sarcoma ewing's|9260/3
C0553580|T191|SY|0000039089|CHV|sarcoma ewings|9260/3
C0553580|T191|PT|NOCODE|COSTAR|Ewing's Sarcoma|9260/3
C0553580|T191|ET|2008-4746|CSP|Ewing's sarcoma|9260/3
C0553580|T191|PT|2008-4746|CSP|Ewing's tumor|9260/3
C0553580|T191|SY|NOCODE|DXP|EWING TUMOR|9260/3
C0553580|T191|DI|U001700|DXP|SARCOMA, EWING|9260/3
C0553580|T191|PT|HP:0012254|HPO|Ewing sarcoma|9260/3
C0553580|T191|SY|HP:0012254|HPO|Ewing sarcoma|9260/3
C0553580|T191|SY|HP:0012254|HPO|Ewing's sarcoma|9260/3
C0553580|T191|PT|sh85046050|LCH_NW|Ewing's sarcoma|9260/3
C0553580|T191|PT|10015560|MDR|Ewing's sarcoma|9260/3
C0553580|T191|LLT|10015560|MDR|Ewing's sarcoma|9260/3
C0553580|T191|LLT|10015563|MDR|Ewing's sarcoma NOS|9260/3
C0553580|T191|LLT|10015565|MDR|Ewing's sarcoma stage unspecified|9260/3
C0553580|T191|LLT|10015566|MDR|Ewing's tumor|9260/3
C0553580|T191|LLT|10015570|MDR|Ewing's tumour|9260/3
C0553580|T191|ET|169|MEDLINEPLUS|Ewing's Sarcoma|9260/3
C0553580|T191|ET|169|MEDLINEPLUS|Sarcoma, Ewing's|9260/3
C0553580|T191|ET|D012512|MSH|Ewing Sarcoma|9260/3
C0553580|T191|ET|D012512|MSH|Ewing Tumor|9260/3
C0553580|T191|ET|D012512|MSH|Ewing's Sarcoma|9260/3
C0553580|T191|ET|D012512|MSH|Ewing's Tumor|9260/3
C0553580|T191|PM|D012512|MSH|Ewings Sarcoma|9260/3
C0553580|T191|PM|D012512|MSH|Ewings Tumor|9260/3
C0553580|T191|MH|D012512|MSH|Sarcoma, Ewing|9260/3
C0553580|T191|ET|D012512|MSH|Sarcoma, Ewing's|9260/3
C0553580|T191|PM|D012512|MSH|Sarcoma, Ewings|9260/3
C0553580|T191|PM|D012512|MSH|Tumor, Ewing|9260/3
C0553580|T191|PM|D012512|MSH|Tumor, Ewing's|9260/3
C0553580|T191|PN|NOCODE|MTH|Ewings sarcoma|9260/3
C0553580|T191|SY|C4817|NCI|ES|9260/3
C0553580|T191|PT|C4817|NCI|Ewing Sarcoma|9260/3
C0553580|T191|SY|C4817|NCI|Ewing's Sarcoma|9260/3
C0553580|T191|SY|C4817|NCI|Ewing's Tumor|9260/3
C0553580|T191|PT|C4817|NCI_CPTAC|Ewing Sarcoma|9260/3
C0553580|T191|PT|C4817|NCI_CTRP|Ewing Sarcoma|9260/3
C0553580|T191|DN|C4817|NCI_CTRP|Ewing Sarcoma|9260/3
C0553580|T191|PT|CDR0000046031|NCI_NCI-GLOSS|Ewing sarcoma|9260/3
C0553580|T191|PT|C4817|NCI_NICHD|Ewing Sarcoma|9260/3
C0553580|T191|PT|CDR0000546979|PDQ|Ewing sarcoma|9260/3
C0553580|T191|SY|CDR0000546979|PDQ|Ewing's Sarcoma|9260/3
C0553580|T191|SY|CDR0000546979|PDQ|Ewing's Tumor|9260/3
C0553580|T191|PT|BBY0.|RCD|Ewing's sarcoma|9260/3
C0553580|T191|SY|BBY0.|RCD|Ewing's tumour|9260/3
C0553580|T191|SY|BBY0.|RCDAE|Ewing's tumor|9260/3
C0553580|T191|SY|76909002|SNOMEDCT_US|Ewing sarcoma|9260/3
C0553580|T191|PT|76909002|SNOMEDCT_US|Ewing's sarcoma|9260/3
C0553580|T191|SY|76909002|SNOMEDCT_US|Ewing's tumor|9260/3
C0553580|T191|SYGB|76909002|SNOMEDCT_US|Ewing's tumour|9260/3
C0334556|T191|PT|MTHU003260|ICPC2ICD10ENG|adamantinoma; long bones|9261/3
C1273017|T191|PT|MTHU003265|ICPC2ICD10ENG|adamantinoma; tibia|9261/3
C0334556|T191|PT|MTHU005183|ICPC2ICD10ENG|ameloblastoma; long bones|9261/3
C1273017|T191|PT|MTHU005188|ICPC2ICD10ENG|ameloblastoma; tibia|9261/3
C0334556|T191|PT|MTHU042858|ICPC2ICD10ENG|long bones; adamantinoma|9261/3
C0334556|T191|PT|MTHU042859|ICPC2ICD10ENG|long bones; ameloblastoma|9261/3
C1273017|T191|PT|MTHU074214|ICPC2ICD10ENG|tibia; adamantinoma|9261/3
C1273017|T191|PT|MTHU074216|ICPC2ICD10ENG|tibia; ameloblastoma|9261/3
C0334556|T191|SY|356678|MEDCIN|bone neoplasm malignant adamantinoma of long bone|9261/3
C1273017|T191|SY|356694|MEDCIN|bone neoplasm, malignant - long bones of lower limb tibial adamantinoma|9261/3
C0334556|T191|PT|356678|MEDCIN|malignant adamantinoma of long bone|9261/3
C1273017|T191|PT|356694|MEDCIN|Tibial adamantinoma|9261/3
C1367554|T191|MH|D050398|MSH|Adamantinoma|9261/3
C0334556|T191|NM|C562741|MSH|Adamantinoma Of Long Bones|9261/3
C1367554|T191|PM|D050398|MSH|Adamantinomas|9261/3
C1367554|T191|PN|NOCODE|MTH|Adamantinoma|9261/3
C0334556|T191|PN|NOCODE|MTH|Adamantinoma of Long Bones|9261/3
C1273017|T191|PN|NOCODE|MTH|Tibial adamantinoma|9261/3
C1367554|T191|PT|C7644|NCI|Adamantinoma|9261/3
C1367554|T191|SY|C7644|NCI|Adamantinoma of Long Bones|9261/3
C1367554|T191|SY|C7644|NCI|Extragnathic Adamantinoma|9261/3
C1273017|T191|PT|C8461|NCI|Tibial Adamantinoma|9261/3
C1367554|T191|SY|C7644|NCI_CDISC|Adamantinoma|9261/3
C1367554|T191|PT|C7644|NCI_CDISC|ADAMANTINOMA, MALIGNANT|9261/3
C0334556|T191|PT|XaBB2|RCD|Adamantinoma of long bone|9261/3
C0334556|T191|SY|XE1wZ|RCD|Adamantinoma of long bones|9261/3
C1273017|T191|OP|Xa1qs|RCD|Tibial adamantinoma|9261/3
C0334556|T191|PT|307609003|SNOMEDCT_US|Adamantinoma of long bone|9261/3
C0334556|T191|PT|56763007|SNOMEDCT_US|Adamantinoma of long bones|9261/3
C1273017|T191|PT|281702006|SNOMEDCT_US|Tibial adamantinoma|9261/3
C1273017|T191|SY|210233007|SNOMEDCT_US|Tibial adamantinoma|9261/3
C1273017|T191|IS|56763007|SNOMEDCT_US|Tibial adamantinoma|9261/3
C1273017|T191|PT|210233007|SNOMEDCT_US|Tibial adamantinoma morphology|9261/3
C0206640|T191|SY|0000020988|CHV|fibro osteoma|9262/0
C0206640|T191|SY|0000020988|CHV|fibro-osteoma|9262/0
C0206640|T191|SY|0000020988|CHV|fibroma ossified|9262/0
C0206640|T191|PT|0000020988|CHV|ossifying fibroma|9262/0
C0206640|T191|SY|0000020988|CHV|ossifying fibromas|9262/0
C0206640|T191|PT|HP:0030426|HPO|Ossifying fibroma|9262/0
C0206640|T191|MH|D018214|MSH|Fibroma, Ossifying|9262/0
C0206640|T191|PM|D018214|MSH|Fibromas, Ossifying|9262/0
C0206640|T191|PM|D018214|MSH|Ossifying Fibroma|9262/0
C0206640|T191|PM|D018214|MSH|Ossifying Fibromas|9262/0
C0206640|T191|PN|NOCODE|MTH|Ossifying Fibroma|9262/0
C0206640|T191|SY|C8422|NCI|Cementifying Fibroma|9262/0
C0206640|T191|SY|C8422|NCI|Cemento-Ossifying Fibroma|9262/0
C0206640|T191|PT|C8422|NCI|Ossifying Fibroma|9262/0
C0206640|T191|SY|C8422|NCI_CDISC|Cementifying Fibroma|9262/0
C0206640|T191|SY|C8422|NCI_CDISC|Cemento-Ossifying Fibroma|9262/0
C0206640|T191|PT|C8422|NCI_CDISC|FIBROMA, OSSIFYING, BENIGN|9262/0
C0206640|T191|SY|C8422|NCI_CDISC|Ossifying Fibroma|9262/0
C0206640|T191|OP|BBZ6.|RCD|Cementifying fibroma|9262/0
C0206640|T191|PT|Xa9Ag|RCD|Cemento-ossifying fibroma|9262/0
C0206640|T191|PT|Xa9Ae|RCD|Fibro-osteoma|9262/0
C0206640|T191|OP|BBY2.|RCD|Ossifying fibroma|9262/0
C0206640|T191|PT|80699009|SNOMEDCT_US|Cementifying fibroma|9262/0
C0206640|T191|SY|80699009|SNOMEDCT_US|Cementifying fibroma, calcified structure|9262/0
C0206640|T191|PT|302863006|SNOMEDCT_US|Cemento-ossifying fibroma|9262/0
C0206640|T191|SY|80699009|SNOMEDCT_US|Cemento-ossifying fibroma|9262/0
C0206640|T191|SY|25603007|SNOMEDCT_US|Fibro-osteoma|9262/0
C0206640|T191|PT|302862001|SNOMEDCT_US|Fibro-osteoma|9262/0
C0206640|T191|SY|302862001|SNOMEDCT_US|Ossifying fibroma|9262/0
C0206640|T191|PT|25603007|SNOMEDCT_US|Ossifying fibroma|9262/0
C0206640|T191|OAP|189896007|SNOMEDCT_US|Ossifying fibroma|9262/0
C0206640|T191|SY|25603007|SNOMEDCT_US|Ossifying fibroma, calcified structure|9262/0
C0206640|T191|SY|0000020988|CHV|fibro osteoma|9270/0
C0206640|T191|SY|0000020988|CHV|fibro-osteoma|9270/0
C0206640|T191|SY|0000020988|CHV|fibroma ossified|9270/0
C0206640|T191|PT|0000020988|CHV|ossifying fibroma|9270/0
C0206640|T191|SY|0000020988|CHV|ossifying fibromas|9270/0
C0206640|T191|PT|HP:0030426|HPO|Ossifying fibroma|9270/0
C0334557|T191|PT|MTHU053955|ICPC2ICD10ENG|odontogenic; tumor, benign|9270/0
C0334557|T191|PT|MTHU077111|ICPC2ICD10ENG|tumor; odontogenic, benign|9270/0
C0206640|T191|MH|D018214|MSH|Fibroma, Ossifying|9270/0
C0206640|T191|PM|D018214|MSH|Fibromas, Ossifying|9270/0
C0206640|T191|PM|D018214|MSH|Ossifying Fibroma|9270/0
C0206640|T191|PM|D018214|MSH|Ossifying Fibromas|9270/0
C0206640|T191|PN|NOCODE|MTH|Ossifying Fibroma|9270/0
C0334557|T191|PT|C4306|NCI|Benign Odontogenic Neoplasm|9270/0
C0334557|T191|SY|C4306|NCI|Benign Odontogenic Tumor|9270/0
C0206640|T191|SY|C8422|NCI|Cementifying Fibroma|9270/0
C0206640|T191|SY|C8422|NCI|Cemento-Ossifying Fibroma|9270/0
C0206640|T191|PT|C8422|NCI|Ossifying Fibroma|9270/0
C0334557|T191|SY|C4306|NCI_CDISC|Benign Odontogenic Tumor|9270/0
C0206640|T191|SY|C8422|NCI_CDISC|Cementifying Fibroma|9270/0
C0206640|T191|SY|C8422|NCI_CDISC|Cemento-Ossifying Fibroma|9270/0
C0206640|T191|PT|C8422|NCI_CDISC|FIBROMA, OSSIFYING, BENIGN|9270/0
C0334557|T191|PT|C4306|NCI_CDISC|ODONTOGENIC TUMOR, BENIGN|9270/0
C0206640|T191|SY|C8422|NCI_CDISC|Ossifying Fibroma|9270/0
C0334557|T191|DN|C4306|NCI_CTRP|Benign Odontogenic Tumor|9270/0
C0334557|T191|PT|BBZ0.|RCD|Benign odontogenic tumour|9270/0
C0206640|T191|OP|BBZ6.|RCD|Cementifying fibroma|9270/0
C0206640|T191|PT|Xa9Ag|RCD|Cemento-ossifying fibroma|9270/0
C0206640|T191|PT|Xa9Ae|RCD|Fibro-osteoma|9270/0
C0206640|T191|OP|BBY2.|RCD|Ossifying fibroma|9270/0
C0334557|T191|PT|BBZ0.|RCDAE|Benign odontogenic tumor|9270/0
C0334557|T191|SY|74839008|SNOMEDCT_US|Benign odontogenic tumor|9270/0
C0334557|T191|SYGB|74839008|SNOMEDCT_US|Benign odontogenic tumour|9270/0
C0206640|T191|PT|80699009|SNOMEDCT_US|Cementifying fibroma|9270/0
C0206640|T191|SY|80699009|SNOMEDCT_US|Cementifying fibroma, calcified structure|9270/0
C0206640|T191|PT|302863006|SNOMEDCT_US|Cemento-ossifying fibroma|9270/0
C0206640|T191|SY|80699009|SNOMEDCT_US|Cemento-ossifying fibroma|9270/0
C0206640|T191|PT|302862001|SNOMEDCT_US|Fibro-osteoma|9270/0
C0206640|T191|SY|25603007|SNOMEDCT_US|Fibro-osteoma|9270/0
C3698372|T191|PT|699228001|SNOMEDCT_US|Focal cemento-osseous dysplasia|9270/0
C3698372|T191|SY|715634002|SNOMEDCT_US|Focal cemento-osseous dysplasia|9270/0
C0334557|T191|PT|74839008|SNOMEDCT_US|Odontogenic tumor, benign|9270/0
C0334557|T191|PTGB|74839008|SNOMEDCT_US|Odontogenic tumour, benign|9270/0
C0206640|T191|PT|25603007|SNOMEDCT_US|Ossifying fibroma|9270/0
C0206640|T191|OAP|189896007|SNOMEDCT_US|Ossifying fibroma|9270/0
C0206640|T191|SY|302862001|SNOMEDCT_US|Ossifying fibroma|9270/0
C0206640|T191|SY|25603007|SNOMEDCT_US|Ossifying fibroma, calcified structure|9270/0
C0457523|T191|PT|0000036730|CHV|cemento-osseous dysplasia|9270/1
C0028880|T191|SY|0000008908|CHV|odontogenic tumor|9270/1
C0028880|T191|PT|0000008908|CHV|odontogenic tumors|9270/1
C0028880|T191|SY|0000008908|CHV|odontogenic tumour|9270/1
C0028880|T191|ET|2013-2197|CSP|odontogenic tumor|9270/1
C0028880|T191|PT|HP:0100612|HPO|Odontogenic neoplasm|9270/1
C0028880|T191|SY|HP:0100612|HPO|Odontogenic tumor|9270/1
C0028880|T191|PT|MTHU053952|ICPC2ICD10ENG|odontogenic; tumor|9270/1
C0028880|T191|PT|MTHU077108|ICPC2ICD10ENG|tumor; odontogenic|9270/1
C0028880|T191|PT|U003325|LCH|Odontogenic tumors|9270/1
C0028880|T191|PT|sh85094100|LCH_NW|Odontogenic tumors|9270/1
C0457523|T191|LLT|10070313|MDR|Cemento osseous dysplasia|9270/1
C0457523|T191|PT|10070313|MDR|Cemento osseous dysplasia|9270/1
C0028880|T191|PT|219011|MEDCIN|odontogenic neoplasms|9270/1
C0028880|T191|PM|D009808|MSH|Odontogenic Tumor|9270/1
C0028880|T191|MH|D009808|MSH|Odontogenic Tumors|9270/1
C0028880|T191|PM|D009808|MSH|Tumor, Odontogenic|9270/1
C0028880|T191|PM|D009808|MSH|Tumors, Odontogenic|9270/1
C0028880|T191|PT|C3286|NCI|Odontogenic Neoplasm|9270/1
C0028880|T191|SY|C3286|NCI|Odontogenic Tumor|9270/1
C0028880|T191|DN|C3286|NCI_CTRP|Odontogenic Tumor|9270/1
C0457523|T191|PT|Xa0hn|RCD|Cemento-osseous dysplasia|9270/1
C0028880|T191|PT|BBZ..|RCD|Odontogenic tumour|9270/1
C0028880|T191|PT|BBZ..|RCDAE|Odontogenic tumor|9270/1
C0028880|T191|OP|BBZz.|RCDSA|Odontogenic tumor NOS|9270/1
C0028880|T191|OP|BBZz.|RCDSY|Odontogenic tumour NOS|9270/1
C0457523|T191|PT|278389000|SNOMEDCT_US|Cemento-osseous dysplasia|9270/1
C0028880|T191|SY|127578009|SNOMEDCT_US|Odontogenic neoplasm|9270/1
C0028880|T191|OAP|3833004|SNOMEDCT_US|Odontogenic tumor|9270/1
C0028880|T191|IS|3833004|SNOMEDCT_US|Odontogenic tumor, NOS|9270/1
C0028880|T191|OAP|3833004|SNOMEDCT_US|Odontogenic tumour|9270/1
C0334558|T191|PT|MTHU014805|ICPC2ICD10ENG|carcinoma; odontogenic|9270/3
C0334558|T191|PT|MTHU053936|ICPC2ICD10ENG|odontogenic; carcinoma|9270/3
C0334558|T191|PT|MTHU053957|ICPC2ICD10ENG|odontogenic; tumor, malignant|9270/3
C0334558|T191|PT|MTHU077114|ICPC2ICD10ENG|tumor; odontogenic, malignant|9270/3
C0334558|T191|PN|NOCODE|MTH|Malignant odontogenic tumor|9270/3
C1333260|T191|PT|C7493|NCI|Ameloblastic Carcinoma-Primary Type|9270/3
C1333260|T191|SY|C7493|NCI|De novo Ameloblastic Carcinoma|9270/3
C0334558|T191|PT|C4812|NCI|Malignant Odontogenic Neoplasm|9270/3
C0334558|T191|SY|C4812|NCI|Malignant Odontogenic Tumor|9270/3
C0334558|T191|SY|C4812|NCI|Odontogenic Carcinoma|9270/3
C0334558|T191|SY|C4812|NCI|Odontogenic Carcinosarcoma|9270/3
C1333260|T191|SY|C7493|NCI|Primary Ameloblastic Carcinoma|9270/3
C1335487|T191|SY|C7500|NCI|Primary Intraosseous Carcinoma Ex Odontogenic Cyst|9270/3
C1335486|T191|SY|C7491|NCI|Primary Intraosseous Squamous Cell Carcinoma Arising de novo|9270/3
C1335487|T191|PT|C7500|NCI|Primary Intraosseous Squamous Cell Carcinoma Derived From Odontogenic Cyst|9270/3
C1335486|T191|PT|C7491|NCI|Primary Intraosseous Squamous Cell Carcinoma-Solid Type|9270/3
C0334558|T191|SY|C4812|NCI_CDISC|Malignant Odontogenic Tumor|9270/3
C0334558|T191|SY|C4812|NCI_CDISC|Odontogenic Carcinoma|9270/3
C0334558|T191|SY|C4812|NCI_CDISC|Odontogenic Carcinosarcoma|9270/3
C0334558|T191|PT|C4812|NCI_CDISC|ODONTOMA, MALIGNANT|9270/3
C0334558|T191|DN|C4812|NCI_CTRP|Malignant Odontogenic Tumor|9270/3
C0334558|T191|PT|BBZ2.|RCD|Malignant odontogenic tumour|9270/3
C0334558|T191|PT|Xa0hk|RCD|Odontogenic carcinoma|9270/3
C0457542|T191|AB|Xa0iA|RCD|Primary intra-osseous carcinom|9270/3
C0457542|T191|PT|Xa0iA|RCD|Primary intra-osseous carcinoma|9270/3
C0334558|T191|PT|BBZ2.|RCDAE|Malignant odontogenic tumor|9270/3
C0334558|T191|SY|128780003|SNOMEDCT_US|Ameloblastic carcinosarcoma|9270/3
C0334558|T191|SY|26888009|SNOMEDCT_US|Carcinoma arising in an odontogenic cyst|9270/3
C0334558|T191|SY|26888009|SNOMEDCT_US|Malignant odontogenic tumor|9270/3
C0334558|T191|SYGB|26888009|SNOMEDCT_US|Malignant odontogenic tumour|9270/3
C0334558|T191|OAP|278386007|SNOMEDCT_US|Odontogenic carcinoma|9270/3
C0334558|T191|OF|278386007|SNOMEDCT_US|Odontogenic carcinoma|9270/3
C0334558|T191|SY|26888009|SNOMEDCT_US|Odontogenic carcinoma|9270/3
C0334558|T191|PT|128780003|SNOMEDCT_US|Odontogenic carcinosarcoma|9270/3
C0334558|T191|PT|26888009|SNOMEDCT_US|Odontogenic tumor, malignant|9270/3
C0334558|T191|PTGB|26888009|SNOMEDCT_US|Odontogenic tumour, malignant|9270/3
C1333260|T191|PT|773624006|SNOMEDCT_US|Primary ameloblastic carcinoma|9270/3
C1333260|T191|PT|733414001|SNOMEDCT_US|Primary ameloblastic carcinoma|9270/3
C0457542|T191|PT|278411006|SNOMEDCT_US|Primary intra-osseous carcinoma|9270/3
C0457542|T191|SY|26888009|SNOMEDCT_US|Primary intraosseous carcinoma|9270/3
C4518390|T191|PT|733913003|SNOMEDCT_US|Primary intraosseous squamous cell carcinoma derived from keratocystic odontogenic neoplasm|9270/3
C1335487|T191|PT|733912008|SNOMEDCT_US|Primary intraosseous squamous cell carcinoma derived from odontogenic cyst|9270/3
C1335486|T191|PT|734095001|SNOMEDCT_US|Primary solid type intraosseous squamous cell carcinoma|9270/3
C4518366|T191|PT|734064008|SNOMEDCT_US|Secondary dedifferentiated intraosseous ameloblastic carcinoma|9270/3
C4518365|T191|PT|734063002|SNOMEDCT_US|Secondary dedifferentiated peripheral ameloblastic carcinoma|9270/3
C0457520|T191|PT|MTHU022348|ICPC2ICD10ENG|dentinoma|9271/0
C0457520|T191|PN|NOCODE|MTH|Ameloblastic fibrodentinoma|9271/0
C0457520|T191|PT|C66800|NCI|Ameloblastic Fibrodentinoma|9271/0
C0457520|T191|PT|Xa0hi|RCD|Ameloblastic fibrodentinoma|9271/0
C0457520|T191|PT|BBZ3.|RCD|Dentinoma|9271/0
C0457520|T191|IS|6437002|SNOMEDCT_US|Ameloblastic fibrodentinoma|9271/0
C0457520|T191|OAP|134311009|SNOMEDCT_US|Ameloblastic fibrodentinoma|9271/0
C0457520|T191|OF|134311009|SNOMEDCT_US|Ameloblastic fibrodentinoma|9271/0
C0457520|T191|PT|6437002|SNOMEDCT_US|Ameloblastic fibrodentinoma|9271/0
C0457520|T191|SY|6437002|SNOMEDCT_US|Dentinoma|9271/0
C0007659|T191|PT|0000030006|CHV|cementoblastoma|9272/0
C0007659|T191|PT|0000002613|CHV|cementoma|9272/0
C0007659|T191|SY|0000002613|CHV|cementomas|9272/0
C0007659|T191|SY|0000002613|CHV|periapical cemental dysplasia|9272/0
C0007659|T191|PT|HP:0012328|HPO|Cementoma|9272/0
C0007659|T191|PT|MTHU015428|ICPC2ICD10ENG|cementoblastoma; benign|9272/0
C0007659|T191|PT|MTHU015430|ICPC2ICD10ENG|cementoma|9272/0
C0007659|T191|LLT|10062564|MDR|Cementoblastoma|9272/0
C0007659|T191|PT|10062564|MDR|Cementoblastoma|9272/0
C0007659|T191|PM|D002485|MSH|Cemento Ossifying Fibroma|9272/0
C0007659|T191|ET|D002485|MSH|Cemento-Ossifying Fibroma|9272/0
C0007659|T191|PM|D002485|MSH|Cemento-Ossifying Fibromas|9272/0
C0007659|T191|MH|D002485|MSH|Cementoma|9272/0
C0007659|T191|PM|D002485|MSH|Cementomas|9272/0
C0007659|T191|PM|D002485|MSH|Dysplasia, Periapical Fibrous|9272/0
C0007659|T191|PM|D002485|MSH|Fibroma, Cemento-Ossifying|9272/0
C0007659|T191|PM|D002485|MSH|Fibrous Dysplasia, Periapical|9272/0
C0007659|T191|PM|D002485|MSH|Fibrous Dysplasias, Periapical|9272/0
C0007659|T191|ET|D002485|MSH|Periapical Fibrous Dysplasia|9272/0
C0007659|T191|PM|D002485|MSH|Periapical Fibrous Dysplasias|9272/0
C0007659|T191|PN|NOCODE|MTH|Cementoma|9272/0
C0007659|T191|SY|C4308|NCI|Benign Cementoblastoma|9272/0
C0007659|T191|PT|C4308|NCI|Cementoblastoma|9272/0
C0007659|T191|SY|C4308|NCI|Cementoma|9272/0
C0007659|T191|PT|BBZ5.|RCD|Benign cementoblastoma|9272/0
C0007659|T191|SY|BBZ5.|RCD|Cementoblastoma|9272/0
C0007659|T191|PT|Xa9Af|RCD|Cementoma|9272/0
C0007659|T191|PT|Xa0ho|RCD|Periapical cemental dysplasia|9272/0
C0007659|T191|SY|Xa0ho|RCD|Periapical fibrous dysplasia|9272/0
C0007659|T191|SY|BBZ5.|RCD|True cementoma|9272/0
C0007659|T191|OP|BBZ4.|RCDSY|Cementoma NOS|9272/0
C0007659|T191|SY|23255001|SNOMEDCT_US|Benign cementoblastoma|9272/0
C0007659|T191|SY|23255001|SNOMEDCT_US|Cementoblastoma|9272/0
C0007659|T191|PT|23255001|SNOMEDCT_US|Cementoblastoma, benign|9272/0
C0007659|T191|PT|37258009|SNOMEDCT_US|Cementoma|9272/0
C0007659|T191|IS|37258009|SNOMEDCT_US|Cementoma, NOS|9272/0
C0007659|T191|SY|37258009|SNOMEDCT_US|Periapical cemental dysplasia|9272/0
C0007659|T191|OAP|278390009|SNOMEDCT_US|Periapical cemental dysplasia|9272/0
C0007659|T191|OF|278390009|SNOMEDCT_US|Periapical cemental dysplasia|9272/0
C0007659|T191|SY|37258009|SNOMEDCT_US|Periapical cemento-osseous dysplasia|9272/0
C0007659|T191|OAS|278390009|SNOMEDCT_US|Periapical fibrous dysplasia|9272/0
C0007659|T191|SY|37258009|SNOMEDCT_US|Periradicular cemental dysplasia|9272/0
C0007659|T191|SY|23255001|SNOMEDCT_US|True cementoma|9272/0
C0007659|T191|PT|0000030006|CHV|cementoblastoma|9273/0
C0007659|T191|PT|0000002613|CHV|cementoma|9273/0
C0007659|T191|SY|0000002613|CHV|cementomas|9273/0
C0007659|T191|SY|0000002613|CHV|periapical cemental dysplasia|9273/0
C0007659|T191|PT|HP:0012328|HPO|Cementoma|9273/0
C0007659|T191|PT|MTHU015428|ICPC2ICD10ENG|cementoblastoma; benign|9273/0
C0007659|T191|PT|MTHU015430|ICPC2ICD10ENG|cementoma|9273/0
C0007659|T191|LLT|10062564|MDR|Cementoblastoma|9273/0
C0007659|T191|PT|10062564|MDR|Cementoblastoma|9273/0
C0007659|T191|PM|D002485|MSH|Cemento Ossifying Fibroma|9273/0
C0007659|T191|ET|D002485|MSH|Cemento-Ossifying Fibroma|9273/0
C0007659|T191|PM|D002485|MSH|Cemento-Ossifying Fibromas|9273/0
C0007659|T191|MH|D002485|MSH|Cementoma|9273/0
C0007659|T191|PM|D002485|MSH|Cementomas|9273/0
C0007659|T191|PM|D002485|MSH|Dysplasia, Periapical Fibrous|9273/0
C0007659|T191|PM|D002485|MSH|Fibroma, Cemento-Ossifying|9273/0
C0007659|T191|PM|D002485|MSH|Fibrous Dysplasia, Periapical|9273/0
C0007659|T191|PM|D002485|MSH|Fibrous Dysplasias, Periapical|9273/0
C0007659|T191|ET|D002485|MSH|Periapical Fibrous Dysplasia|9273/0
C0007659|T191|PM|D002485|MSH|Periapical Fibrous Dysplasias|9273/0
C0007659|T191|PN|NOCODE|MTH|Cementoma|9273/0
C0007659|T191|SY|C4308|NCI|Benign Cementoblastoma|9273/0
C0007659|T191|PT|C4308|NCI|Cementoblastoma|9273/0
C0007659|T191|SY|C4308|NCI|Cementoma|9273/0
C0007659|T191|PT|BBZ5.|RCD|Benign cementoblastoma|9273/0
C0007659|T191|SY|BBZ5.|RCD|Cementoblastoma|9273/0
C0007659|T191|PT|Xa9Af|RCD|Cementoma|9273/0
C0007659|T191|PT|Xa0ho|RCD|Periapical cemental dysplasia|9273/0
C0007659|T191|SY|Xa0ho|RCD|Periapical fibrous dysplasia|9273/0
C0007659|T191|SY|BBZ5.|RCD|True cementoma|9273/0
C0007659|T191|OP|BBZ4.|RCDSY|Cementoma NOS|9273/0
C0007659|T191|SY|23255001|SNOMEDCT_US|Benign cementoblastoma|9273/0
C0007659|T191|SY|23255001|SNOMEDCT_US|Cementoblastoma|9273/0
C0007659|T191|PT|23255001|SNOMEDCT_US|Cementoblastoma, benign|9273/0
C0007659|T191|PT|37258009|SNOMEDCT_US|Cementoma|9273/0
C0007659|T191|IS|37258009|SNOMEDCT_US|Cementoma, NOS|9273/0
C0007659|T191|SY|37258009|SNOMEDCT_US|Periapical cemental dysplasia|9273/0
C0007659|T191|OAP|278390009|SNOMEDCT_US|Periapical cemental dysplasia|9273/0
C0007659|T191|OF|278390009|SNOMEDCT_US|Periapical cemental dysplasia|9273/0
C0007659|T191|SY|37258009|SNOMEDCT_US|Periapical cemento-osseous dysplasia|9273/0
C0007659|T191|OAS|278390009|SNOMEDCT_US|Periapical fibrous dysplasia|9273/0
C0007659|T191|SY|37258009|SNOMEDCT_US|Periradicular cemental dysplasia|9273/0
C0007659|T191|SY|23255001|SNOMEDCT_US|True cementoma|9273/0
C0206640|T191|SY|0000020988|CHV|fibro osteoma|9274/0
C0206640|T191|SY|0000020988|CHV|fibro-osteoma|9274/0
C0206640|T191|SY|0000020988|CHV|fibroma ossified|9274/0
C0206640|T191|PT|0000020988|CHV|ossifying fibroma|9274/0
C0206640|T191|SY|0000020988|CHV|ossifying fibromas|9274/0
C0206640|T191|PT|HP:0030426|HPO|Ossifying fibroma|9274/0
C0206640|T191|MH|D018214|MSH|Fibroma, Ossifying|9274/0
C0206640|T191|PM|D018214|MSH|Fibromas, Ossifying|9274/0
C0206640|T191|PM|D018214|MSH|Ossifying Fibroma|9274/0
C0206640|T191|PM|D018214|MSH|Ossifying Fibromas|9274/0
C0206640|T191|PN|NOCODE|MTH|Ossifying Fibroma|9274/0
C0206640|T191|SY|C8422|NCI|Cementifying Fibroma|9274/0
C0206640|T191|SY|C8422|NCI|Cemento-Ossifying Fibroma|9274/0
C0206640|T191|PT|C8422|NCI|Ossifying Fibroma|9274/0
C0206640|T191|SY|C8422|NCI_CDISC|Cementifying Fibroma|9274/0
C0206640|T191|SY|C8422|NCI_CDISC|Cemento-Ossifying Fibroma|9274/0
C0206640|T191|PT|C8422|NCI_CDISC|FIBROMA, OSSIFYING, BENIGN|9274/0
C0206640|T191|SY|C8422|NCI_CDISC|Ossifying Fibroma|9274/0
C0206640|T191|OP|BBZ6.|RCD|Cementifying fibroma|9274/0
C0206640|T191|PT|Xa9Ag|RCD|Cemento-ossifying fibroma|9274/0
C0206640|T191|PT|Xa9Ae|RCD|Fibro-osteoma|9274/0
C0206640|T191|OP|BBY2.|RCD|Ossifying fibroma|9274/0
C0206640|T191|PT|80699009|SNOMEDCT_US|Cementifying fibroma|9274/0
C0206640|T191|SY|80699009|SNOMEDCT_US|Cementifying fibroma, calcified structure|9274/0
C0206640|T191|SY|80699009|SNOMEDCT_US|Cemento-ossifying fibroma|9274/0
C0206640|T191|PT|302863006|SNOMEDCT_US|Cemento-ossifying fibroma|9274/0
C0206640|T191|PT|302862001|SNOMEDCT_US|Fibro-osteoma|9274/0
C0206640|T191|SY|25603007|SNOMEDCT_US|Fibro-osteoma|9274/0
C0206640|T191|PT|25603007|SNOMEDCT_US|Ossifying fibroma|9274/0
C0206640|T191|OAP|189896007|SNOMEDCT_US|Ossifying fibroma|9274/0
C0206640|T191|SY|302862001|SNOMEDCT_US|Ossifying fibroma|9274/0
C0206640|T191|SY|25603007|SNOMEDCT_US|Ossifying fibroma, calcified structure|9274/0
C3495361|T191|PT|MTHU015432|ICPC2ICD10ENG|cementoma; gigantiform|9275/0
C3495361|T191|PT|MTHU031979|ICPC2ICD10ENG|gigantiform; cementoma|9275/0
C3495361|T191|LLT|10081225|MDR|Familial gigantiform cementoma|9275/0
C3495361|T191|PT|10081225|MDR|Familial gigantiform cementoma|9275/0
C3495361|T191|CE|C563017|MSH|Cemental Dysplasia, Periapical|9275/0
C3495361|T191|CE|C563017|MSH|Cementomas, Familial Multiple|9275/0
C3495361|T191|NM|C563017|MSH|Gigantiform Cementoma, Familial|9275/0
C3495361|T191|PN|NOCODE|MTH|Gigantiform Cementoma, Familial|9275/0
C3495361|T191|SY|C8381|NCI|Florid Osseous Dysplasia|9275/0
C3495361|T191|PT|C8381|NCI|Gigantiform Cementoma|9275/0
C3495361|T191|OP|BBZ7.|RCD|Gigantiform cementoma|9275/0
C3495361|T191|SY|63937004|SNOMEDCT_US|Familial multiple cementoma|9275/0
C3495361|T191|OAP|189900005|SNOMEDCT_US|Gigantiform cementoma|9275/0
C3495361|T191|PT|63937004|SNOMEDCT_US|Gigantiform cementoma|9275/0
C0028882|T191|PT|0000008910|CHV|odontoma|9280/0
C0028882|T191|SY|0000008910|CHV|odontomas|9280/0
C0028882|T191|PT|HP:0011068|HPO|Odontoma|9280/0
C0028882|T191|ET|HP:0011068|HPO|Odontomas|9280/0
C0028882|T191|PT|MTHU053965|ICPC2ICD10ENG|odontoma|9280/0
C0028882|T191|PT|30770|MEDCIN|odontoma|9280/0
C0028882|T191|PM|D009810|MSH|Fibro Odontoma|9280/0
C0028882|T191|ET|D009810|MSH|Fibro-Odontoma|9280/0
C0028882|T191|PM|D009810|MSH|Fibro-Odontomas|9280/0
C0028882|T191|ET|D009810|MSH|Fibroodontoma|9280/0
C0028882|T191|PM|D009810|MSH|Fibroodontomas|9280/0
C0028882|T191|MH|D009810|MSH|Odontoma|9280/0
C0028882|T191|PM|D009810|MSH|Odontomas|9280/0
C0028882|T191|SY|C3287|NCI|Fibro-Odontoma|9280/0
C0028882|T191|SY|C3287|NCI|Fibroodontoma|9280/0
C0028882|T191|PT|C3287|NCI|Odontoma|9280/0
C0028882|T191|SY|C3287|NCI_CDISC|Fibro-Odontoma|9280/0
C0028882|T191|SY|C3287|NCI_CDISC|Fibroodontoma|9280/0
C0028882|T191|PT|C3287|NCI_CDISC|ODONTOMA, BENIGN|9280/0
C0028882|T191|PT|Xa9Ai|RCD|Odontoma|9280/0
C0028882|T191|OP|BBZ8.|RCDSY|Odontoma NOS|9280/0
C0028882|T191|PT|79074005|SNOMEDCT_US|Odontoma|9280/0
C0028882|T191|SY|79074005|SNOMEDCT_US|Odontoma, no ICD-O subtype|9280/0
C0028882|T191|SY|79074005|SNOMEDCT_US|Odontoma, no International Classification of Diseases for Oncology subtype|9280/0
C0028882|T191|IS|79074005|SNOMEDCT_US|Odontoma, NOS|9280/0
C0205866|T191|PT|MTHU065820|ICPC2ICD10ENG|compound; odontoma|9281/0
C0205866|T191|PT|MTHU053973|ICPC2ICD10ENG|odontoma; compound|9281/0
C0205866|T191|PM|D009810|MSH|Compound Odontoma|9281/0
C0205866|T191|PM|D009810|MSH|Compound Odontomas|9281/0
C0205866|T191|PEP|D009810|MSH|Odontoma, Compound|9281/0
C0205866|T191|PM|D009810|MSH|Odontomas, Compound|9281/0
C0205866|T191|PT|C3711|NCI|Compound Odontoma|9281/0
C0205866|T191|PT|BBZ9.|RCD|Compound odontoma|9281/0
C0205866|T191|PT|28733007|SNOMEDCT_US|Compound odontoma|9281/0
C0334563|T191|PT|MTHU017385|ICPC2ICD10ENG|complex; odontoma|9282/0
C0334563|T191|PT|MTHU053969|ICPC2ICD10ENG|odontoma; complex|9282/0
C0334563|T191|PT|C4309|NCI|Complex Odontoma|9282/0
C0334563|T191|PT|BBZA.|RCD|Complex odontoma|9282/0
C0334563|T191|PT|29020002|SNOMEDCT_US|Complex odontoma|9282/0
C0205865|T191|PT|MTHU028207|ICPC2ICD10ENG|fibro-odontoma; ameloblastic|9290/0
C0205865|T191|PT|MTHU028170|ICPC2ICD10ENG|fibroameloblastic; odontoma|9290/0
C0205865|T191|PT|MTHU053971|ICPC2ICD10ENG|odontoma; fibroameloblastic|9290/0
C0205865|T191|PM|D009810|MSH|Ameloblastic Fibro-odontoma|9290/0
C0205865|T191|PM|D009810|MSH|Ameloblastic Fibro-odontomas|9290/0
C0205865|T191|PM|D009810|MSH|Fibro odontoma, Ameloblastic|9290/0
C0205865|T191|PEP|D009810|MSH|Fibro-odontoma, Ameloblastic|9290/0
C0205865|T191|PM|D009810|MSH|Fibro-odontomas, Ameloblastic|9290/0
C0205865|T191|DSV|D009810|MSH|FIBROODONTOMA AMELOBLASTIC|9290/0
C0205865|T191|PT|C3710|NCI|Ameloblastic Fibro-Odontoma|9290/0
C0205865|T191|SY|C3710|NCI|Ameloblastic Fibroodontoma|9290/0
C0205865|T191|SY|C3710|NCI|Fibroameloblastic Odontoma|9290/0
C0205865|T191|SY|C3710|NCI_CDISC|Ameloblastic Fibroodontoma|9290/0
C0205865|T191|SY|C3710|NCI_CDISC|Fibroameloblastic Odontoma|9290/0
C0205865|T191|PT|C3710|NCI_CDISC|ODONTOMA, AMELOBLASTIC, BENIGN|9290/0
C0205865|T191|PT|BBZB.|RCD|Ameloblastic fibro-odontoma|9290/0
C0205865|T191|SY|BBZB.|RCD|Fibroameloblastic odontoma|9290/0
C0205865|T191|PT|84983008|SNOMEDCT_US|Ameloblastic fibro-odontoma|9290/0
C0205865|T191|SY|84983008|SNOMEDCT_US|Fibroameloblastic odontoma|9290/0
C0334573|T191|PT|MTHU005174|ICPC2ICD10ENG|ameloblastic; fibrosarcoma|9290/3
C0334573|T191|PT|MTHU005178|ICPC2ICD10ENG|ameloblastic; sarcoma|9290/3
C0334573|T191|PT|MTHU028226|ICPC2ICD10ENG|fibrosarcoma; ameloblastic|9290/3
C0334573|T191|PT|MTHU028231|ICPC2ICD10ENG|fibrosarcoma; odontogenic|9290/3
C0334573|T191|PT|MTHU053943|ICPC2ICD10ENG|odontogenic; fibrosarcoma|9290/3
C0334564|T191|PT|MTHU053976|ICPC2ICD10ENG|odontosarcoma; ameloblastic|9290/3
C0334573|T191|PT|MTHU065886|ICPC2ICD10ENG|sarcoma; ameloblastic|9290/3
C0334573|T191|PT|C4317|NCI|Ameloblastic Fibrosarcoma|9290/3
C0334573|T191|SY|C4317|NCI|Ameloblastic Sarcoma|9290/3
C0334573|T191|SY|C4317|NCI|Odontogenic Fibrosarcoma|9290/3
C0334573|T191|PT|BBZN.|RCD|Ameloblastic fibrosarcoma|9290/3
C0334564|T191|PT|BBZC.|RCD|Ameloblastic odontosarcoma|9290/3
C0334573|T191|SY|BBZN.|RCD|Ameloblastic sarcoma|9290/3
C0334573|T191|SY|BBZN.|RCD|Odontogenic fibrosarcoma|9290/3
C0334564|T191|SY|20380000|SNOMEDCT_US|Ameloblastic dentinosarcoma|9290/3
C0334564|T191|SY|20380000|SNOMEDCT_US|Ameloblastic fibro-odontosarcoma|9290/3
C0334564|T191|SY|20380000|SNOMEDCT_US|Ameloblastic fibrodentinosarcoma|9290/3
C0334573|T191|PT|27092008|SNOMEDCT_US|Ameloblastic fibrosarcoma|9290/3
C0334564|T191|PT|20380000|SNOMEDCT_US|Ameloblastic odontosarcoma|9290/3
C0334573|T191|SY|27092008|SNOMEDCT_US|Ameloblastic sarcoma|9290/3
C0334573|T191|SY|27092008|SNOMEDCT_US|Odontogenic fibrosarcoma|9290/3
C0334565|T191|PT|MTHU003364|ICPC2ICD10ENG|adenoameloblastoma|9300/0
C0334565|T191|PT|MTHU003457|ICPC2ICD10ENG|adenomatoid; odontogenic tumor|9300/0
C0334565|T191|PT|MTHU003459|ICPC2ICD10ENG|adenomatoid; tumor, odontogenic|9300/0
C0334565|T191|PT|MTHU053953|ICPC2ICD10ENG|odontogenic; tumor, adenomatoid|9300/0
C0334565|T191|PT|MTHU077009|ICPC2ICD10ENG|tumor; adenomatoid, odontogenic|9300/0
C0334565|T191|PT|MTHU077109|ICPC2ICD10ENG|tumor; odontogenic, adenomatoid|9300/0
C0334565|T191|NM|C538229|MSH|Adenoameloblastoma|9300/0
C0334565|T191|CE|C538229|MSH|Adenomatoid ameloblastoma|9300/0
C0334565|T191|CE|C538229|MSH|Adenomatoid odontogenic tumor|9300/0
C0334565|T191|CE|C538229|MSH|Pleomorphic adenomatoid tumor|9300/0
C0334565|T191|SY|C4310|NCI|Adenomatoid Odontogenic Neoplasm|9300/0
C0334565|T191|PT|C4310|NCI|Adenomatoid Odontogenic Tumor|9300/0
C0334565|T191|SY|BBZD.|RCD|Adenoameloblastoma|9300/0
C0334565|T191|PT|BBZD.|RCD|Adenomatoid odontogenic tumour|9300/0
C0334565|T191|PT|BBZD.|RCDAE|Adenomatoid odontogenic tumor|9300/0
C0334565|T191|SY|60599006|SNOMEDCT_US|Adenoameloblastoma|9300/0
C0334565|T191|PT|60599006|SNOMEDCT_US|Adenomatoid odontogenic tumor|9300/0
C0334565|T191|PTGB|60599006|SNOMEDCT_US|Adenomatoid odontogenic tumour|9300/0
C0206740|T190|PT|MTHU079883|ICPC2ICD10ENG|calcifying; cyst, odontogenic|9301/0
C0206740|T190|PT|MTHU079887|ICPC2ICD10ENG|calcifying; odontogenic cyst|9301/0
C0206740|T190|PT|MTHU020736|ICPC2ICD10ENG|cyst; calcifying odontogenic|9301/0
C0206740|T190|PM|D018333|MSH|Calcifying Odontogenic Cyst|9301/0
C0206740|T190|PM|D018333|MSH|Calcifying Odontogenic Cysts|9301/0
C0206740|T190|PM|D018333|MSH|Cyst, Calcifying Odontogenic|9301/0
C0206740|T190|PM|D018333|MSH|Cysts, Calcifying Odontogenic|9301/0
C0206740|T190|MH|D018333|MSH|Odontogenic Cyst, Calcifying|9301/0
C0206740|T190|PM|D018333|MSH|Odontogenic Cysts, Calcifying|9301/0
C0206740|T190|PN|NOCODE|MTH|Calcifying Odontogenic Cyst|9301/0
C0206740|T190|PT|C54319|NCI|Calcifying Cystic Odontogenic Tumor|9301/0
C0206740|T190|SY|C54319|NCI|Calcifying Odontogenic Cyst|9301/0
C0206740|T190|SY|C54319|NCI|Gorlin Cyst|9301/0
C0206740|T190|PT|BBZE.|RCD|Calcifying odontogenic cyst|9301/0
C0206740|T190|PT|75248003|SNOMEDCT_US|Calcifying odontogenic cyst|9301/0
C1704219|T191|PN|NOCODE|MTH|Dentinogenic Ghost Cell Tumor|9302/0
C1704219|T191|SY|C54323|NCI|Calcifying Ghost Cell Odontogenic Tumor|9302/0
C1704219|T191|SY|C54323|NCI|Dentinoameloblastoma|9302/0
C1704219|T191|PT|C54323|NCI|Dentinogenic Ghost Cell Tumor|9302/0
C1704219|T191|SY|C54323|NCI|Dentinoma|9302/0
C1704219|T191|SY|C54323|NCI|Odontogenic Ghost Cell Tumor|9302/0
C1704219|T191|DN|C54323|NCI_CTRP|Dentinogenic Ghost Cell Tumor|9302/0
C1704219|T191|SY|X77pE|RCD|Deninogenic ghost cell tumour|9302/0
C1704219|T191|PT|X77pE|RCD|Odontogenic ghost cell tumour|9302/0
C1704219|T191|SY|X77pE|RCDAE|Deninogenic ghost cell tumor|9302/0
C1704219|T191|PT|X77pE|RCDAE|Odontogenic ghost cell tumor|9302/0
C5229855|T191|SY|788590006|SNOMEDCT_US|Benign dentinogenic ghost cell neoplasm|9302/0
C5229855|T191|SY|788590006|SNOMEDCT_US|Benign dentinogenic ghost cell tumor|9302/0
C5229855|T191|SYGB|788590006|SNOMEDCT_US|Benign dentinogenic ghost cell tumour|9302/0
C5229855|T191|PT|788590006|SNOMEDCT_US|Benign odontogenic ghost cell neoplasm|9302/0
C5229855|T191|SY|788590006|SNOMEDCT_US|Benign odontogenic ghost cell tumor|9302/0
C5229855|T191|SYGB|788590006|SNOMEDCT_US|Benign odontogenic ghost cell tumour|9302/0
C1704219|T191|IS|67978001|SNOMEDCT_US|Deninogenic ghost cell tumor|9302/0
C1704219|T191|IS|67978001|SNOMEDCT_US|Deninogenic ghost cell tumour|9302/0
C1704219|T191|SY|788592003|SNOMEDCT_US|Dentinogenic ghost cell neoplasm|9302/0
C1704219|T191|OAS|67978001|SNOMEDCT_US|Dentinogenic ghost cell tumor|9302/0
C1704219|T191|SY|788592003|SNOMEDCT_US|Dentinogenic ghost cell tumor|9302/0
C1704219|T191|OAS|67978001|SNOMEDCT_US|Dentinogenic ghost cell tumour|9302/0
C1704219|T191|SYGB|788592003|SNOMEDCT_US|Dentinogenic ghost cell tumour|9302/0
C1704219|T191|PT|788592003|SNOMEDCT_US|Odontogenic ghost cell neoplasm|9302/0
C1704219|T191|OAP|67978001|SNOMEDCT_US|Odontogenic ghost cell tumor|9302/0
C1704219|T191|SY|788592003|SNOMEDCT_US|Odontogenic ghost cell tumor|9302/0
C1704219|T191|OAP|67978001|SNOMEDCT_US|Odontogenic ghost cell tumour|9302/0
C1704219|T191|SYGB|788592003|SNOMEDCT_US|Odontogenic ghost cell tumour|9302/0
C0334566|T191|PT|354170|MEDCIN|odontogenic ghost cell carcinoma|9302/3
C0334566|T191|PN|NOCODE|MTH|Ghost Cell Odontogenic Carcinoma|9302/3
C0334566|T191|PT|C4311|NCI|Ghost Cell Odontogenic Carcinoma|9302/3
C0334566|T191|SY|C4311|NCI|Odontogenic Ghost Cell Neoplasm|9302/3
C0334566|T191|AB|Xa0iB|RCD|Odontogenic ghost cell carc|9302/3
C0334566|T191|PT|Xa0iB|RCD|Odontogenic ghost cell carcinoma|9302/3
C1266170|T191|PT|110458000|SNOMEDCT_US|Malignant odontogenic ghost cell tumor|9302/3
C1266170|T191|PTGB|110458000|SNOMEDCT_US|Malignant odontogenic ghost cell tumour|9302/3
C0334566|T191|PT|788580003|SNOMEDCT_US|Odontogenic ghost cell carcinoma|9302/3
C0334566|T191|PT|134312002|SNOMEDCT_US|Odontogenic ghost cell carcinoma|9302/3
C0002448|T191|SY|0000000986|CHV|adamantinoma|9310/0
C0002448|T191|PT|0000000986|CHV|ameloblastoma|9310/0
C0002448|T191|ET|2013-2197|CSP|ameloblastoma|9310/0
C0002448|T191|SY|NOCODE|DXP|ADAMANTINOMA|9310/0
C0002448|T191|DI|U000076|DXP|AMELOBLASTOMA|9310/0
C0002448|T191|SY|NOCODE|DXP|EPITHELIOMA ADAMANTINUM|9310/0
C0002448|T191|PT|MTHU003257|ICPC2ICD10ENG|adamantinoma|9310/0
C0002448|T191|PT|MTHU005180|ICPC2ICD10ENG|ameloblastoma|9310/0
C0002448|T191|PT|10066796|MDR|Ameloblastoma|9310/0
C0002448|T191|LLT|10066796|MDR|Ameloblastoma|9310/0
C0002448|T191|MH|D000564|MSH|Ameloblastoma|9310/0
C0002448|T191|PM|D000564|MSH|Ameloblastomas|9310/0
C0002448|T191|PN|NOCODE|MTH|Ameloblastoma|9310/0
C0457531|T191|PT|C39754|NCI|Acanthomatous Ameloblastoma|9310/0
C0002448|T191|PT|C4313|NCI|Ameloblastoma|9310/0
C0457521|T191|SY|C39756|NCI|Cystogenic Ameloblastoma|9310/0
C0457533|T191|PT|C39758|NCI|Desmoplastic Ameloblastoma|9310/0
C0457530|T191|PT|C27397|NCI|Follicular Ameloblastoma|9310/0
C0457532|T191|PT|C27398|NCI|Granular Cell Ameloblastoma|9310/0
C0457529|T191|PT|C39753|NCI|Plexiform Ameloblastoma|9310/0
C0457521|T191|PT|C39756|NCI|Unicystic Ameloblastoma|9310/0
C0002448|T191|DN|C4313|NCI_CTRP|Ameloblastoma|9310/0
C0457531|T191|PT|Xa0hx|RCD|Acanthomatous ameloblastoma|9310/0
C0002448|T191|SY|Xa9Aj|RCD|Adamantinoma|9310/0
C0002448|T191|PT|Xa9Aj|RCD|Ameloblastoma|9310/0
C0457533|T191|PT|Xa0hz|RCD|Desmoplastic ameloblastoma|9310/0
C0457530|T191|PT|Xa0hw|RCD|Follicular ameloblastoma|9310/0
C0457532|T191|PT|Xa0hy|RCD|Granular cell ameloblastoma|9310/0
C0457534|T191|PT|Xa0i0|RCD|Keratoameloblastoma|9310/0
C0457540|T191|PT|Xa0i7|RCD|Mural unicystic ameloblastoma|9310/0
C0457536|T191|PT|Xa0i2|RCD|Peripheral ameloblastoma|9310/0
C0457539|T191|AB|Xa0i6|RCD|Plexif unicystic ameloblastoma|9310/0
C0457529|T191|PT|Xa0hv|RCD|Plexiform ameloblastoma|9310/0
C0457539|T191|PT|Xa0i6|RCD|Plexiform unicystic ameloblastoma|9310/0
C0457521|T191|PT|Xa0hj|RCD|Unicystic ameloblastoma|9310/0
C0002448|T191|OP|BBZF.|RCDSY|Ameloblastoma NOS|9310/0
C0457531|T191|PT|278399005|SNOMEDCT_US|Acanthomatous ameloblastoma|9310/0
C0002448|T191|SY|20462008|SNOMEDCT_US|Adamantinoma|9310/0
C0002448|T191|PT|20462008|SNOMEDCT_US|Ameloblastoma|9310/0
C0002448|T191|IS|20462008|SNOMEDCT_US|Ameloblastoma, NOS|9310/0
C0457533|T191|PT|278401004|SNOMEDCT_US|Desmoplastic ameloblastoma|9310/0
C0457530|T191|PT|278398002|SNOMEDCT_US|Follicular ameloblastoma|9310/0
C0457532|T191|PT|278400003|SNOMEDCT_US|Granular cell ameloblastoma|9310/0
C0457534|T191|PT|278402006|SNOMEDCT_US|Keratoameloblastoma|9310/0
C3698009|T191|PT|699226002|SNOMEDCT_US|Luminal unicystic ameloblastoma|9310/0
C0457540|T191|PT|278408005|SNOMEDCT_US|Mural unicystic ameloblastoma|9310/0
C0457536|T191|PT|278404007|SNOMEDCT_US|Peripheral ameloblastoma|9310/0
C0457529|T191|PT|278397007|SNOMEDCT_US|Plexiform ameloblastoma|9310/0
C0457539|T191|PT|278407000|SNOMEDCT_US|Plexiform unicystic ameloblastoma|9310/0
C0457521|T191|PT|278385006|SNOMEDCT_US|Unicystic ameloblastoma|9310/0
C0334567|T191|PT|MTHU003261|ICPC2ICD10ENG|adamantinoma; malignant|9310/3
C0334567|T191|PT|MTHU005184|ICPC2ICD10ENG|ameloblastoma; malignant|9310/3
C0334567|T191|PT|MTHU047261|ICPC2ICD10ENG|malignant; adamantinoma|9310/3
C0334567|T191|PT|MTHU047265|ICPC2ICD10ENG|malignant; ameloblastoma|9310/3
C0334567|T191|PT|271559|MEDCIN|malignant ameloblastoma|9310/3
C0334567|T191|PN|NOCODE|MTH|Malignant Ameloblastoma|9310/3
C0334567|T191|SY|C54297|NCI|Malignant Ameloblastoma|9310/3
C0334567|T191|PT|C54297|NCI|Metastasizing Ameloblastoma|9310/3
C0334567|T191|PT|C54297|NCI_CDISC|AMELOBLASTOMA, MALIGNANT|9310/3
C0334567|T191|SY|C54297|NCI_CDISC|Malignant Ameloblastoma|9310/3
C0334567|T191|SY|BBZG.|RCD|Malignant adamantinoma|9310/3
C0334567|T191|PT|BBZG.|RCD|Malignant ameloblastoma|9310/3
C0334567|T191|PT|88253001|SNOMEDCT_US|Ameloblastoma, malignant|9310/3
C0334567|T191|OAS|134171005|SNOMEDCT_US|Malignant adamantinoma|9310/3
C0334567|T191|SY|88253001|SNOMEDCT_US|Malignant adamantinoma|9310/3
C0334567|T191|SY|88253001|SNOMEDCT_US|Malignant ameloblastoma|9310/3
C0334567|T191|OAP|134171005|SNOMEDCT_US|Malignant ameloblastoma|9310/3
C4518376|T191|PT|734079001|SNOMEDCT_US|Multicystic ameloblastoma|9310/3
C1704220|T191|PT|MTHU005176|ICPC2ICD10ENG|ameloblastic; odontoma|9311/0
C1704220|T191|PT|MTHU053932|ICPC2ICD10ENG|odontoameloblastoma|9311/0
C1704220|T191|PT|MTHU053966|ICPC2ICD10ENG|odontoma; ameloblastic|9311/0
C1704220|T191|PN|NOCODE|MTH|Odontoameloblastoma|9311/0
C1704220|T191|SY|C54317|NCI|Ameloblastic Odontoma|9311/0
C1704220|T191|PT|C54317|NCI|Odontoameloblastoma|9311/0
C1704220|T191|SY|C54317|NCI|Odontoblastoma|9311/0
C1704220|T191|DN|C54317|NCI_CTRP|Odontoameloblastoma|9311/0
C1704220|T191|PT|BBZH.|RCD|Odontoameloblastoma|9311/0
C1704220|T191|SY|84983008|SNOMEDCT_US|Ameloblastic odontoma|9311/0
C1704220|T191|IS|84983008|SNOMEDCT_US|Odontoameloblastoma|9311/0
C1704220|T191|PT|49043004|SNOMEDCT_US|Odontoameloblastoma|9311/0
C1458142|T191|PT|0000057791|CHV|squamous odontogenic tumor|9312/0
C1458142|T191|SY|0000057791|CHV|squamous odontogenic tumour|9312/0
C1458142|T191|MH|D051527|MSH|Odontogenic Tumor, Squamous|9312/0
C1458142|T191|PM|D051527|MSH|Odontogenic Tumors, Squamous|9312/0
C1458142|T191|ET|D051527|MSH|Squamous Odontogenic Tumor|9312/0
C1458142|T191|PM|D051527|MSH|Squamous Odontogenic Tumors|9312/0
C1458142|T191|PM|D051527|MSH|Tumor, Squamous Odontogenic|9312/0
C1458142|T191|PM|D051527|MSH|Tumors, Squamous Odontogenic|9312/0
C1458142|T191|PN|NOCODE|MTH|Squamous odontogenic tumor|9312/0
C1458142|T191|SY|C7112|NCI|Squamous Odontogenic Neoplasm|9312/0
C1458142|T191|PT|C7112|NCI|Squamous Odontogenic Tumor|9312/0
C1458142|T191|PT|BBZJ.|RCD|Squamous odontogenic tumour|9312/0
C1458142|T191|PT|BBZJ.|RCDAE|Squamous odontogenic tumor|9312/0
C1458142|T191|PT|9155002|SNOMEDCT_US|Squamous odontogenic tumor|9312/0
C1458142|T191|PTGB|9155002|SNOMEDCT_US|Squamous odontogenic tumour|9312/0
C0334569|T191|PT|MTHU051311|ICPC2ICD10ENG|myxoma; odontogenic|9320/0
C0334569|T191|PT|MTHU053948|ICPC2ICD10ENG|odontogenic; myxoma|9320/0
C0334569|T191|PT|C7501|NCI|Odontogenic Myxoma|9320/0
C0334569|T191|PT|BBZK.|RCD|Odontogenic myxoma|9320/0
C0334569|T191|PT|34941004|SNOMEDCT_US|Odontogenic myxoma|9320/0
C1260966|T191|PT|MTHU028213|ICPC2ICD10ENG|fibroma; odontogenic|9321/0
C1260966|T191|PT|MTHU053939|ICPC2ICD10ENG|odontogenic; fibroma|9321/0
C1260966|T191|SY|C4314|NCI|Central Odontogenic Fibroma|9321/0
C1260966|T191|PT|C4314|NCI|Odontogenic Fibroma|9321/0
C1260966|T191|SY|C4314|NCI_CDISC|Central Odontogenic Fibroma|9321/0
C1260966|T191|PT|C4314|NCI_CDISC|FIBROMA, ODONTOGENIC, BENIGN|9321/0
C1260966|T191|PT|Xa9Ak|RCD|Central odontogenic fibroma|9321/0
C1260966|T191|SY|Xa9Ak|RCD|Odontogenic fibroma|9321/0
C1260966|T191|OP|BBZL.|RCDSY|Odontogenic fibroma NOS|9321/0
C1260966|T191|PT|88686005|SNOMEDCT_US|Central odontogenic fibroma|9321/0
C1260966|T191|SY|88686005|SNOMEDCT_US|Odontogenic fibroma|9321/0
C1260966|T191|IS|88686005|SNOMEDCT_US|Odontogenic fibroma, NOS|9321/0
C0334571|T191|PT|MTHU028215|ICPC2ICD10ENG|fibroma; odontogenic, peripheral|9322/0
C0334571|T191|PT|MTHU053941|ICPC2ICD10ENG|odontogenic; fibroma, peripheral|9322/0
C0334571|T191|PN|NOCODE|MTH|Peripheral Odontogenic Fibroma|9322/0
C0334571|T191|PT|C4315|NCI|Peripheral Odontogenic Fibroma|9322/0
C0334571|T191|PT|X77pF|RCD|Peripheral odontogenic fibroma|9322/0
C0334571|T191|PT|75914009|SNOMEDCT_US|Peripheral odontogenic fibroma|9322/0
C0334572|T191|PT|MTHU005172|ICPC2ICD10ENG|ameloblastic; fibroma|9330/0
C0334572|T191|PT|MTHU028209|ICPC2ICD10ENG|fibroma; ameloblastic|9330/0
C0334572|T191|PT|C4316|NCI|Ameloblastic Fibroma|9330/0
C0334572|T191|SY|C4316|NCI|Fibrodentinoma|9330/0
C0334572|T191|PT|BBZM.|RCD|Ameloblastic fibroma|9330/0
C0457541|T191|AB|Xa0i8|RCD|Granul cell ameloblast fibroma|9330/0
C0457541|T191|PT|Xa0i8|RCD|Granular cell ameloblastic fibroma|9330/0
C0334572|T191|PT|11063000|SNOMEDCT_US|Ameloblastic fibroma|9330/0
C0457541|T191|PT|278409002|SNOMEDCT_US|Granular cell ameloblastic fibroma|9330/0
C0334573|T191|PT|MTHU005174|ICPC2ICD10ENG|ameloblastic; fibrosarcoma|9330/3
C0334573|T191|PT|MTHU005178|ICPC2ICD10ENG|ameloblastic; sarcoma|9330/3
C0334573|T191|PT|MTHU028226|ICPC2ICD10ENG|fibrosarcoma; ameloblastic|9330/3
C0334573|T191|PT|MTHU028231|ICPC2ICD10ENG|fibrosarcoma; odontogenic|9330/3
C0334573|T191|PT|MTHU053943|ICPC2ICD10ENG|odontogenic; fibrosarcoma|9330/3
C0334573|T191|PT|MTHU065886|ICPC2ICD10ENG|sarcoma; ameloblastic|9330/3
C0334573|T191|PT|C4317|NCI|Ameloblastic Fibrosarcoma|9330/3
C0334573|T191|SY|C4317|NCI|Ameloblastic Sarcoma|9330/3
C0334573|T191|SY|C4317|NCI|Odontogenic Fibrosarcoma|9330/3
C0334573|T191|PT|BBZN.|RCD|Ameloblastic fibrosarcoma|9330/3
C0334573|T191|SY|BBZN.|RCD|Ameloblastic sarcoma|9330/3
C0334573|T191|SY|BBZN.|RCD|Odontogenic fibrosarcoma|9330/3
C0334573|T191|PT|27092008|SNOMEDCT_US|Ameloblastic fibrosarcoma|9330/3
C0334573|T191|SY|27092008|SNOMEDCT_US|Ameloblastic sarcoma|9330/3
C0334573|T191|SY|27092008|SNOMEDCT_US|Odontogenic fibrosarcoma|9330/3
C0334574|T191|PT|MTHU079885|ICPC2ICD10ENG|calcifying; epithelial neoplasm, odontogenic|9340/0
C0334574|T191|PT|MTHU079888|ICPC2ICD10ENG|calcifying; odontogenic epithelial tumor|9340/0
C0334574|T191|PT|MTHU026828|ICPC2ICD10ENG|epithelial; tumor, calcifying, odontogenic|9340/0
C0334574|T191|PT|MTHU053961|ICPC2ICD10ENG|odontogenic; tumor, calcifying epithelial|9340/0
C0334574|T191|PT|MTHU059665|ICPC2ICD10ENG|Pindborg|9340/0
C0334574|T191|PT|MTHU059667|ICPC2ICD10ENG|Pindborg; tumor|9340/0
C0334574|T191|PT|MTHU077177|ICPC2ICD10ENG|tumor; calcifying epithelial odontogenic|9340/0
C0334574|T191|PT|MTHU077118|ICPC2ICD10ENG|tumor; odontogenic, calcifying epithelial|9340/0
C0334574|T191|PT|MTHU077137|ICPC2ICD10ENG|tumor; Pindborg|9340/0
C0334574|T191|NM|C537961|MSH|Calcifying Epithelial Odontogenic Tumor|9340/0
C0334574|T191|CE|C537961|MSH|Pindborg tumor|9340/0
C0334574|T191|PT|C54301|NCI|Calcifying Epithelial Odontogenic Tumor|9340/0
C0334574|T191|SY|C54301|NCI|Pindborg Tumor|9340/0
C0334574|T191|DN|C54301|NCI_CTRP|Calcifying Epithelial Odontogenic Tumor|9340/0
C0334574|T191|PT|CDR0000762523|PDQ|calcifying epithelial odontogenic tumor|9340/0
C0334574|T191|SY|CDR0000762523|PDQ|Pindborg tumor|9340/0
C0334574|T191|AB|BBZP.|RCD|Calcif epithel odontogenic tum|9340/0
C0334574|T191|PT|BBZP.|RCD|Calcifying epithelial odontogenic tumour|9340/0
C0334574|T191|SY|BBZP.|RCD|CEOT - Calcifying epithelial odontogenic tumour|9340/0
C0334574|T191|AB|BBZP.|RCD|CEOT-Calc epith odontogen tum|9340/0
C0334574|T191|SY|BBZP.|RCD|Pindborg tumour|9340/0
C0334574|T191|PT|BBZP.|RCDAE|Calcifying epithelial odontogenic tumor|9340/0
C0334574|T191|SY|BBZP.|RCDAE|CEOT - Calcifying epithelial odontogenic tumor|9340/0
C0334574|T191|SY|BBZP.|RCDAE|Pindborg tumor|9340/0
C0334574|T191|PT|83048004|SNOMEDCT_US|Calcifying epithelial odontogenic tumor|9340/0
C0334574|T191|PTGB|83048004|SNOMEDCT_US|Calcifying epithelial odontogenic tumour|9340/0
C0334574|T191|SY|83048004|SNOMEDCT_US|CEOT - Calcifying epithelial odontogenic tumor|9340/0
C0334574|T191|SYGB|83048004|SNOMEDCT_US|CEOT - Calcifying epithelial odontogenic tumour|9340/0
C0334574|T191|SY|83048004|SNOMEDCT_US|Pindborg tumor|9340/0
C0334574|T191|SYGB|83048004|SNOMEDCT_US|Pindborg tumour|9340/0
C4316837|T191|PN|NOCODE|MTH|Clear cell odontogenic carcinoma|9341/1
C0475829|T191|PN|NOCODE|MTH|Clear cell odontogenic tumor|9341/1
C4316837|T191|SY|C54300|NCI|Clear Cell Ameloblastoma|9341/1
C4316837|T191|PT|C54300|NCI|Clear Cell Odontogenic Carcinoma|9341/1
C4316837|T191|SY|C54300|NCI|Clear Cell Odontogenic Tumor|9341/1
C0475829|T191|PT|Xa0hh|RCD|Clear cell odontogenic tumour|9341/1
C0475829|T191|PT|Xa0hh|RCDAE|Clear cell odontogenic tumor|9341/1
C4316837|T191|PT|734032001|SNOMEDCT_US|Clear cell odontogenic carcinoma|9341/1
C0475829|T191|OAP|134310005|SNOMEDCT_US|Clear cell odontogenic tumor|9341/1
C0475829|T191|PT|128779001|SNOMEDCT_US|Clear cell odontogenic tumor|9341/1
C0475829|T191|OAP|134310005|SNOMEDCT_US|Clear cell odontogenic tumour|9341/1
C0475829|T191|PTGB|128779001|SNOMEDCT_US|Clear cell odontogenic tumour|9341/1
C4316837|T191|PN|NOCODE|MTH|Clear cell odontogenic carcinoma|9341/3
C4316837|T191|SY|C54300|NCI|Clear Cell Ameloblastoma|9341/3
C4316837|T191|PT|C54300|NCI|Clear Cell Odontogenic Carcinoma|9341/3
C4316837|T191|SY|C54300|NCI|Clear Cell Odontogenic Tumor|9341/3
C4316837|T191|PT|734032001|SNOMEDCT_US|Clear cell odontogenic carcinoma|9341/3
C0334558|T191|PT|MTHU014805|ICPC2ICD10ENG|carcinoma; odontogenic|9342/3
C0334558|T191|PT|MTHU053936|ICPC2ICD10ENG|odontogenic; carcinoma|9342/3
C0334558|T191|PT|MTHU053957|ICPC2ICD10ENG|odontogenic; tumor, malignant|9342/3
C0334558|T191|PT|MTHU077114|ICPC2ICD10ENG|tumor; odontogenic, malignant|9342/3
C0334558|T191|PN|NOCODE|MTH|Malignant odontogenic tumor|9342/3
C0334558|T191|PT|C4812|NCI|Malignant Odontogenic Neoplasm|9342/3
C0334558|T191|SY|C4812|NCI|Malignant Odontogenic Tumor|9342/3
C0334558|T191|SY|C4812|NCI|Odontogenic Carcinoma|9342/3
C0334558|T191|SY|C4812|NCI|Odontogenic Carcinosarcoma|9342/3
C0334558|T191|SY|C4812|NCI_CDISC|Malignant Odontogenic Tumor|9342/3
C0334558|T191|SY|C4812|NCI_CDISC|Odontogenic Carcinoma|9342/3
C0334558|T191|SY|C4812|NCI_CDISC|Odontogenic Carcinosarcoma|9342/3
C0334558|T191|PT|C4812|NCI_CDISC|ODONTOMA, MALIGNANT|9342/3
C0334558|T191|DN|C4812|NCI_CTRP|Malignant Odontogenic Tumor|9342/3
C0334558|T191|PT|BBZ2.|RCD|Malignant odontogenic tumour|9342/3
C0334558|T191|PT|Xa0hk|RCD|Odontogenic carcinoma|9342/3
C0334558|T191|PT|BBZ2.|RCDAE|Malignant odontogenic tumor|9342/3
C0334558|T191|SY|128780003|SNOMEDCT_US|Ameloblastic carcinosarcoma|9342/3
C0334558|T191|SY|26888009|SNOMEDCT_US|Carcinoma arising in an odontogenic cyst|9342/3
C0334558|T191|SY|26888009|SNOMEDCT_US|Malignant odontogenic tumor|9342/3
C0334558|T191|SYGB|26888009|SNOMEDCT_US|Malignant odontogenic tumour|9342/3
C0334558|T191|SY|26888009|SNOMEDCT_US|Odontogenic carcinoma|9342/3
C0334558|T191|OAP|278386007|SNOMEDCT_US|Odontogenic carcinoma|9342/3
C0334558|T191|OF|278386007|SNOMEDCT_US|Odontogenic carcinoma|9342/3
C0334558|T191|PT|128780003|SNOMEDCT_US|Odontogenic carcinosarcoma|9342/3
C0334558|T191|PT|26888009|SNOMEDCT_US|Odontogenic tumor, malignant|9342/3
C0334558|T191|PTGB|26888009|SNOMEDCT_US|Odontogenic tumour, malignant|9342/3
C0010276|T191|ET|0000004638|AOD|craniopharyngioma|9350/1
C0010276|T191|PT|0059189|CCPSS|CRANIOPHARYNGIOMA|9350/1
C0010276|T191|PT|0000003431|CHV|craniopharyngioma|9350/1
C0010276|T191|SY|0000003431|CHV|craniopharyngiomas|9350/1
C0010276|T191|SY|0000003431|CHV|rathke pouch tumor|9350/1
C0010276|T191|SY|0000003431|CHV|rathke's pouch tumour|9350/1
C0010276|T191|PT|NOCODE|COSTAR|Craniopharyngioma|9350/1
C0010276|T191|GT|NEOPL CNS|CST|CRANIOPHARYNGIOMA|9350/1
C0010276|T191|SY|NOCODE|DXP|ADAMANTINOMA, PITUITARY|9350/1
C0010276|T191|SY|NOCODE|DXP|BRAIN TUMOR, CRANIOPHARYNGIOMA|9350/1
C0010276|T191|DI|U000414|DXP|CRANIOPHARYNGIOMA|9350/1
C0010276|T191|SY|NOCODE|DXP|INTRACRANIAL NEOPLASM, CRANIOPHARYNGIOMA|9350/1
C0010276|T191|SY|NOCODE|DXP|PITUITARY EPIDERMOID TUMOR|9350/1
C0010276|T191|SY|NOCODE|DXP|RATHKE POUCH TUMOR|9350/1
C0010276|T191|PT|HP:0030062|HPO|Craniopharyngioma|9350/1
C0010276|T191|PT|MTHU019894|ICPC2ICD10ENG|craniopharyngioma|9350/1
C0010276|T191|PT|MTHU063690|ICPC2ICD10ENG|Rathke's pouch; tumor|9350/1
C0010276|T191|PT|MTHU077144|ICPC2ICD10ENG|tumor; Rathke's pouch|9350/1
C0010276|T191|PT|10011318|MDR|Craniopharyngioma|9350/1
C0010276|T191|LLT|10011318|MDR|Craniopharyngioma|9350/1
C0010276|T191|PT|31936|MEDCIN|craniopharyngioma|9350/1
C0010276|T191|MH|D003397|MSH|Craniopharyngioma|9350/1
C0010276|T191|PM|D003397|MSH|Craniopharyngiomas|9350/1
C0010276|T191|DEV|D003397|MSH|NEOPL RATHKE CLEFT|9350/1
C0010276|T191|DEV|D003397|MSH|NEOPL RATHKES CLEFT|9350/1
C0010276|T191|ET|D003397|MSH|Neoplasm, Rathke Cleft|9350/1
C0010276|T191|ET|D003397|MSH|Neoplasm, Rathke's Cleft|9350/1
C0010276|T191|PM|D003397|MSH|Neoplasm, Rathkes Cleft|9350/1
C0010276|T191|DEV|D003397|MSH|RATHKE CLEFT NEOPL|9350/1
C0010276|T191|ET|D003397|MSH|Rathke Cleft Neoplasm|9350/1
C0010276|T191|ET|D003397|MSH|Rathke Pouch Tumor|9350/1
C0010276|T191|ET|D003397|MSH|Rathke's Cleft Neoplasm|9350/1
C0010276|T191|ET|D003397|MSH|Rathke's Pouch Tumor|9350/1
C0010276|T191|DEV|D003397|MSH|RATHKES CLEFT NEOPL|9350/1
C0010276|T191|PM|D003397|MSH|Rathkes Cleft Neoplasm|9350/1
C0010276|T191|PM|D003397|MSH|Rathkes Pouch Tumor|9350/1
C0010276|T191|PM|D003397|MSH|Tumor, Rathke Pouch|9350/1
C0010276|T191|PM|D003397|MSH|Tumor, Rathke's Pouch|9350/1
C0010276|T191|PN|NOCODE|MTH|Craniopharyngioma|9350/1
C0010276|T191|PT|C2964|NCI|Craniopharyngioma|9350/1
C0010276|T191|SY|TCGA|NCI|Craniopharyngioma|9350/1
C0010276|T191|SY|C2964|NCI|Neoplasm of Rathke's Pouch|9350/1
C0010276|T191|SY|C2964|NCI|Rathke Pouch Neoplasm|9350/1
C0010276|T191|SY|C2964|NCI|Rathke Pouch Tumor|9350/1
C0010276|T191|SY|C2964|NCI|Rathke's Pouch Neoplasm|9350/1
C0010276|T191|SY|C2964|NCI|Rathke's Pouch Tumor|9350/1
C0010276|T191|SY|C2964|NCI|Tumor of Rathke's Pouch|9350/1
C0010276|T191|PT|C2964|NCI_CDISC|CRANIOPHARYNGIOMA, BENIGN|9350/1
C0010276|T191|SY|C2964|NCI_CDISC|Cystoma|9350/1
C0010276|T191|SY|C2964|NCI_CDISC|Neoplasm of Rathke's Pouch|9350/1
C0010276|T191|SY|C2964|NCI_CDISC|Rathke Pouch Neoplasm|9350/1
C0010276|T191|SY|C2964|NCI_CDISC|Rathke Pouch Tumor|9350/1
C0010276|T191|SY|C2964|NCI_CDISC|Rathke's Pouch Neoplasm|9350/1
C0010276|T191|SY|C2964|NCI_CDISC|Rathke's Pouch Tumor|9350/1
C0010276|T191|SY|C2964|NCI_CDISC|Tumor of Rathke's Pouch|9350/1
C0010276|T191|PT|C2964|NCI_CPTAC|Craniopharyngioma|9350/1
C0010276|T191|PT|10011318|NCI_CTEP-SDC|Craniopharyngioma|9350/1
C0010276|T191|PT|CDR0000046131|NCI_NCI-GLOSS|craniopharyngioma|9350/1
C0010276|T191|PT|C2964|NCI_NICHD|Craniopharyngioma|9350/1
C0010276|T191|PT|R0121571|QMR|CRANIOPHARYNGIOMA|9350/1
C0010276|T191|PT|B7H21|RCD|Craniopharyngioma|9350/1
C0010276|T191|SY|BBa0.|RCDSA|Rathke's pouch tumor|9350/1
C0010276|T191|PT|BBa0.|RCDSY|Craniopharyngioma|9350/1
C0010276|T191|SY|BBa0.|RCDSY|Rathke's pouch tumour|9350/1
C0010276|T191|PT|189179009|SNOMEDCT_US|Craniopharyngioma|9350/1
C0010276|T191|PT|40009002|SNOMEDCT_US|Craniopharyngioma|9350/1
C0010276|T191|SY|40009002|SNOMEDCT_US|Rathke's pouch tumor|9350/1
C0010276|T191|SYGB|40009002|SNOMEDCT_US|Rathke's pouch tumour|9350/1
C0010276|T191|PT|1550|WHO|CRANIOPHARYNGIOMA|9350/1
C0431129|T191|PM|D003397|MSH|Adamantinous Craniopharyngioma|9351/1
C0431129|T191|PM|D003397|MSH|Adamantinous Craniopharyngiomas|9351/1
C0431129|T191|PEP|D003397|MSH|Craniopharyngioma, Adamantinous|9351/1
C0431129|T191|PM|D003397|MSH|Craniopharyngiomas, Adamantinous|9351/1
C0431129|T191|PN|NOCODE|MTH|Adamantinous Craniopharyngioma|9351/1
C0431129|T191|AB|C4726|NCI|ACP|9351/1
C0431129|T191|PT|C4726|NCI|Adamantinomatous Craniopharyngioma|9351/1
C0431129|T191|SY|TCGA|NCI|Adamantinomatous Craniopharyngioma|9351/1
C0431129|T191|SY|C4726|NCI|Adamantinous Craniopharyngioma|9351/1
C0431129|T191|SY|C4726|NCI|Adamantinous Neoplasm of Rathke's Pouch|9351/1
C0431129|T191|SY|C4726|NCI|Adamantinous Rathke's Pouch Neoplasm|9351/1
C0431129|T191|SY|C4726|NCI|Adamantinous Rathke's Pouch Tumor|9351/1
C0431129|T191|SY|C4726|NCI|Adamantinous Tumor of Rathke's Pouch|9351/1
C0431129|T191|PT|X77q2|RCD|Adamantinous craniopharyngioma|9351/1
C0431129|T191|SY|128781004|SNOMEDCT_US|Adamantinous craniopharyngioma|9351/1
C0431129|T191|OAP|134216001|SNOMEDCT_US|Adamantinous craniopharyngioma|9351/1
C0431129|T191|PT|128781004|SNOMEDCT_US|Craniopharyngioma, adamantinomatous|9351/1
C0431128|T191|PEP|D003397|MSH|Craniopharyngioma, Papillary|9352/1
C0431128|T191|PM|D003397|MSH|Craniopharyngiomas, Papillary|9352/1
C0431128|T191|PM|D003397|MSH|Papillary Craniopharyngioma|9352/1
C0431128|T191|PM|D003397|MSH|Papillary Craniopharyngiomas|9352/1
C0431128|T191|PN|NOCODE|MTH|Papillary craniopharyngioma|9352/1
C0431128|T191|SY|TCGA|NCI|Papillary Craniopharyngioma|9352/1
C0431128|T191|PT|C4725|NCI|Papillary Craniopharyngioma|9352/1
C0431128|T191|SY|C4725|NCI|Papillary Neoplasm of Rathke's Pouch|9352/1
C0431128|T191|SY|C4725|NCI|Papillary Rathke Pouch Neoplasm|9352/1
C0431128|T191|SY|C4725|NCI|Papillary Rathke's Pouch Neoplasm|9352/1
C0431128|T191|SY|C4725|NCI|Papillary Rathke's Pouch Tumor|9352/1
C0431128|T191|SY|C4725|NCI|Papillary Tumor of Rathke's Pouch|9352/1
C0431128|T191|AB|C4725|NCI|PCP|9352/1
C0431128|T191|PT|X77q1|RCD|Papillary craniopharyngioma|9352/1
C0431128|T191|PT|128782006|SNOMEDCT_US|Craniopharyngioma, papillary|9352/1
C0431128|T191|OAP|134215002|SNOMEDCT_US|Papillary craniopharyngioma|9352/1
C0431128|T191|SY|128782006|SNOMEDCT_US|Papillary craniopharyngioma|9352/1
C0031941|T191|SY|0000009743|CHV|gland pineal tumor|9360/1
C0031941|T191|SY|0000009743|CHV|gland pineal tumors|9360/1
C0031941|T191|SY|0000009743|CHV|gland pineal tumours|9360/1
C0031941|T191|SY|0000009743|CHV|pineal gland tumor|9360/1
C0031941|T191|SY|0000009743|CHV|pineal gland tumour|9360/1
C0031941|T191|SY|0000009743|CHV|pineal region tumor|9360/1
C0031941|T191|SY|0000009743|CHV|pineal region tumors|9360/1
C0031941|T191|PT|0000009743|CHV|pineal tumor|9360/1
C0031941|T191|SY|0000009743|CHV|pineal tumors|9360/1
C0031941|T191|SY|0000009743|CHV|pinealoma|9360/1
C0031941|T191|PT|NOCODE|COSTAR|Pinealoma|9360/1
C0031941|T191|PT|2006-6484|CSP|pineal body neoplasm|9360/1
C0031941|T191|ET|2006-6484|CSP|pinealoma|9360/1
C0031941|T191|SY|NOCODE|DXP|BRAIN TUMOR, PINEAL GLAND|9360/1
C0031941|T191|SY|NOCODE|DXP|INTRACRANIAL NEOPLASM, PINEAL GLAND|9360/1
C0031941|T191|DI|U001502|DXP|PINEAL GLAND, TUMOR|9360/1
C0031941|T191|PT|HP:0030694|HPO|Pineal parenchymal cell neoplasm|9360/1
C0031941|T191|SY|HP:0030693|HPO|Pineal parenchymal tumor|9360/1
C0031941|T191|SY|HP:0030693|HPO|Pineal parenchymal tumour|9360/1
C0031941|T191|PT|HP:0010799|HPO|Pinealoma|9360/1
C0031941|T191|PT|MTHU059669|ICPC2ICD10ENG|pinealoma|9360/1
C0031941|T191|PT|sh85102234|LCH_NW|Pineal gland--Tumors|9360/1
C0031941|T191|PT|10061348|MDR|Pineal neoplasm|9360/1
C0031941|T191|LLT|10061348|MDR|Pineal neoplasm|9360/1
C0031941|T191|LLT|10035053|MDR|Pineal neoplasm NOS|9360/1
C0031941|T191|LLT|10035057|MDR|Pinealoma|9360/1
C0031941|T191|PT|10035057|MDR|Pinealoma|9360/1
C0031941|T191|PT|31940|MEDCIN|benign pinealoma|9360/1
C0031941|T191|SY|355521|MEDCIN|neoplasm of endocrine gland pineal|9360/1
C0031941|T191|PT|355521|MEDCIN|Neoplasm of pineal gland|9360/1
C0031941|T191|SY|355648|MEDCIN|neoplasm uncertain behavior pinealoma|9360/1
C0031941|T191|PT|355648|MEDCIN|pinealoma|9360/1
C0031941|T191|DEV|D010871|MSH|NEOPL PINEAL|9360/1
C0031941|T191|PM|D010871|MSH|Neoplasm, Pineal|9360/1
C0031941|T191|ET|D010871|MSH|Neoplasms, Pineal|9360/1
C0031941|T191|ET|D010871|MSH|Pineal Gland Tumor|9360/1
C0031941|T191|PM|D010871|MSH|Pineal Gland Tumors|9360/1
C0031941|T191|DEV|D010871|MSH|PINEAL NEOPL|9360/1
C0031941|T191|PM|D010871|MSH|Pineal Neoplasm|9360/1
C0031941|T191|ET|D010871|MSH|Pineal Neoplasms|9360/1
C0031941|T191|PM|D010871|MSH|Pineal Parenchymal Tumor|9360/1
C0031941|T191|ET|D010871|MSH|Pineal Parenchymal Tumors|9360/1
C0031941|T191|PM|D010871|MSH|Pineal Tumor|9360/1
C0031941|T191|ET|D010871|MSH|Pineal Tumors|9360/1
C0031941|T191|MH|D010871|MSH|Pinealoma|9360/1
C0031941|T191|PM|D010871|MSH|Pinealomas|9360/1
C0031941|T191|PM|D010871|MSH|Tumor, Pineal|9360/1
C0031941|T191|PM|D010871|MSH|Tumor, Pineal Gland|9360/1
C0031941|T191|PM|D010871|MSH|Tumor, Pineal Parenchymal|9360/1
C0031941|T191|PM|D010871|MSH|Tumors, Pineal|9360/1
C0031941|T191|PM|D010871|MSH|Tumors, Pineal Gland|9360/1
C0031941|T191|PM|D010871|MSH|Tumors, Pineal Parenchymal|9360/1
C0031941|T191|PN|NOCODE|MTH|Pineal Gland Neoplasm|9360/1
C0031941|T191|SY|C6965|NCI|Neoplasm of Pineal Gland|9360/1
C0031941|T191|SY|C6965|NCI|Neoplasm of the Pineal Gland|9360/1
C0031941|T191|SY|C6965|NCI|Pineal Gland Neoplasm|9360/1
C0031941|T191|SY|C6965|NCI|Pineal Gland Tumor|9360/1
C0031941|T191|PT|C6965|NCI|Pineal Parenchymal Cell Neoplasm|9360/1
C0031941|T191|SY|C6965|NCI|Pineal Parenchymal Cell Tumor|9360/1
C0031941|T191|SY|C6965|NCI|Pineal Parenchymal Neoplasm|9360/1
C0031941|T191|SY|C6965|NCI|Pineal Parenchymal Tumor|9360/1
C0031941|T191|SY|C6965|NCI|Pineocytic Neoplasm|9360/1
C0031941|T191|SY|C6965|NCI|Pineocytic Tumor|9360/1
C0031941|T191|SY|C6965|NCI|Tumor of Pineal Gland|9360/1
C0031941|T191|SY|C6965|NCI|Tumor of the Pineal Gland|9360/1
C0031941|T191|PT|10035054|NCI_CTEP-SDC|Pineal parenchymal tumor|9360/1
C0031941|T191|SY|X40P4|RCD|Pineal tumour|9360/1
C0031941|T191|SY|X40P4|RCD|Pinealoma|9360/1
C0031941|T191|PT|X40P4|RCD|Tumour of pineal gland|9360/1
C0031941|T191|SY|X40P4|RCDAE|Pineal tumor|9360/1
C0031941|T191|PT|X40P4|RCDAE|Tumor of pineal gland|9360/1
C0031941|T191|PT|127026004|SNOMEDCT_US|Neoplasm of pineal gland|9360/1
C0031941|T191|SY|127026004|SNOMEDCT_US|Pineal tumor|9360/1
C0031941|T191|SYGB|127026004|SNOMEDCT_US|Pineal tumour|9360/1
C0031941|T191|OAP|47598005|SNOMEDCT_US|Pinealoma|9360/1
C0031941|T191|PT|359619007|SNOMEDCT_US|Pinealoma|9360/1
C0031941|T191|SY|127026004|SNOMEDCT_US|Tumor of pineal gland|9360/1
C0031941|T191|SYGB|127026004|SNOMEDCT_US|Tumour of pineal gland|9360/1
C0917890|T191|SY|0000052373|CHV|pinealocytoma|9361/1
C0917890|T191|PT|0000052373|CHV|pineocytoma|9361/1
C0917890|T191|SY|0000052373|CHV|pineocytomas|9361/1
C0917890|T191|PT|HP:0030407|HPO|Pineocytoma|9361/1
C0917890|T191|PT|MTHU059671|ICPC2ICD10ENG|pineocytoma|9361/1
C0917890|T191|LLT|10035059|MDR|Pineocytoma|9361/1
C0917890|T191|PT|10035059|MDR|Pineocytoma|9361/1
C0917890|T191|PT|35001|MEDCIN|pineocytoma|9361/1
C0917890|T191|PEP|D010871|MSH|Pinealocytoma|9361/1
C0917890|T191|PM|D010871|MSH|Pinealocytomas|9361/1
C0917890|T191|ET|D010871|MSH|Pineocytoma|9361/1
C0917890|T191|PM|D010871|MSH|Pineocytomas|9361/1
C0917890|T191|PN|NOCODE|MTH|Pineocytoma|9361/1
C0917890|T191|SY|TCGA|NCI|Pineocytoma|9361/1
C0917890|T191|PT|C6966|NCI|Pineocytoma|9361/1
C0917890|T191|SY|C6966|NCI_CDISC|Benign Pinealoma|9361/1
C0917890|T191|PT|C6966|NCI_CDISC|PINEOCYTOMA, BENIGN|9361/1
C0917890|T191|PT|CDR0000046228|NCI_NCI-GLOSS|pineocytoma|9361/1
C0917890|T191|SY|C6966|NCI_NICHD|Benign Pinealoma|9361/1
C0917890|T191|SY|C6966|NCI_NICHD|Pinealocytoma|9361/1
C0917890|T191|PT|C6966|NCI_NICHD|Pineocytoma|9361/1
C0917890|T191|PT|X78dZ|RCD|Benign pinealoma|9361/1
C0917890|T191|PT|BBa2.|RCD|Pineocytoma|9361/1
C0917890|T191|OAP|255045009|SNOMEDCT_US|Benign pinealoma|9361/1
C0917890|T191|PT|89096009|SNOMEDCT_US|Pineocytoma|9361/1
C0205898|T191|SY|0000020745|CHV|pinealblastoma|9362/3
C0205898|T191|SY|0000020745|CHV|pinealoblastoma|9362/3
C0205898|T191|PT|0000020745|CHV|pineoblastoma|9362/3
C0205898|T191|SY|HP:0030408|HPO|Pinealoblastoma|9362/3
C0205898|T191|PT|HP:0030408|HPO|Pineoblastoma|9362/3
C0205898|T191|PT|MTHU059670|ICPC2ICD10ENG|pineoblastoma|9362/3
C0205898|T191|LLT|10035056|MDR|Pinealblastoma|9362/3
C0205898|T191|LLT|10050487|MDR|Pinealoblastoma|9362/3
C0205898|T191|PT|10050487|MDR|Pinealoblastoma|9362/3
C0205898|T191|LLT|10035058|MDR|Pineoblastoma|9362/3
C0205898|T191|SY|35000|MEDCIN|pineoblastoma|9362/3
C0205898|T191|PT|35000|MEDCIN|pineoblastoma of pineal body|9362/3
C0205898|T191|PEP|D010871|MSH|Pineoblastoma|9362/3
C0205898|T191|PM|D010871|MSH|Pineoblastomas|9362/3
C1367859|T191|PN|NOCODE|MTH|Pineal parenchymal tumor of intermediate differentiation|9362/3
C0205898|T191|PN|NOCODE|MTH|pineoblastoma|9362/3
C0205898|T191|SY|C9344|NCI|Pineal Gland PNET|9362/3
C0205898|T191|SY|C9344|NCI|Pineal Gland Primitive Neuroectodermal Neoplasm|9362/3
C0205898|T191|SY|C9344|NCI|Pineal Gland Primitive Neuroectodermal Tumor|9362/3
C1367859|T191|PT|C6967|NCI|Pineal Parenchymal Tumor of Intermediate Differentiation|9362/3
C1367859|T191|SY|TCGA|NCI|Pineal Parenchymal Tumor of Intermediate Differentiation|9362/3
C0205898|T191|SY|C9344|NCI|Pineal PNET|9362/3
C0205898|T191|SY|C9344|NCI|Pineal Primitive Neuroectodermal Neoplasm|9362/3
C0205898|T191|SY|C9344|NCI|Pineal Primitive Neuroectodermal Tumor|9362/3
C0205898|T191|SY|TCGA|NCI|Pineoblastoma|9362/3
C0205898|T191|PT|C9344|NCI|Pineoblastoma|9362/3
C0205898|T191|SY|C9344|NCI|PNET of Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI|PNET of the Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI|Primitive Neuroectodermal Neoplasm of Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI|Primitive Neuroectodermal Neoplasm of the Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI|Primitive Neuroectodermal Tumor of Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI|Primitive Neuroectodermal Tumor of the Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Pineal Gland PNET|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Pineal Gland Primitive Neuroectodermal Neoplasm|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Pineal Gland Primitive Neuroectodermal Tumor|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Pineal PNET|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Pineal Primitive Neuroectodermal Neoplasm|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Pineal Primitive Neuroectodermal Tumor|9362/3
C0205898|T191|PT|C9344|NCI_CDISC|PINEOBLASTOMA, MALIGNANT|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|PNET of Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|PNET of the Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Primitive Neuroectodermal Neoplasm of Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Primitive Neuroectodermal Neoplasm of the Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Primitive Neuroectodermal Tumor of Pineal Gland|9362/3
C0205898|T191|SY|C9344|NCI_CDISC|Primitive Neuroectodermal Tumor of the Pineal Gland|9362/3
C0205898|T191|PT|C9344|NCI_CPTAC|Pineoblastoma|9362/3
C0205898|T191|DN|C9344|NCI_CTRP|Pineoblastoma|9362/3
C0205898|T191|PT|C9344|NCI_CTRP|Pineoblastoma|9362/3
C0205898|T191|PT|CDR0000046227|NCI_NCI-GLOSS|pineoblastoma|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Pineal Gland PNET|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Pineal Gland Primitive Neuroectodermal Neoplasm|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Pineal Gland Primitive Neuroectodermal Tumor|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Pineal PNET|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Pineal Primitive Neuroectodermal Neoplasm|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Pineal Primitive Neuroectodermal Tumor|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Pineoblastoma|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|PNET of Pineal Gland|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|PNET of the Pineal Gland|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Primitive Neuroectodermal Neoplasm of Pineal Gland|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Primitive Neuroectodermal Neoplasm of the Pineal Gland|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Primitive Neuroectodermal Tumor of Pineal Gland|9362/3
C0205898|T191|SY|CDR0000562070|PDQ|Primitive Neuroectodermal Tumor of the Pineal Gland|9362/3
C0205898|T191|PT|BBa3.|RCD|Pineoblastoma|9362/3
C1367859|T191|SY|31671006|SNOMEDCT_US|Pineal parenchymal tumor of intermediate differentiation|9362/3
C1367859|T191|PT|715904005|SNOMEDCT_US|Pineal parenchymal tumor of intermediate differentiation|9362/3
C1367859|T191|PT|397379005|SNOMEDCT_US|Pineal parenchymal tumor of intermediate differentiation|9362/3
C1367859|T191|PTGB|715904005|SNOMEDCT_US|Pineal parenchymal tumour of intermediate differentiation|9362/3
C1367859|T191|PTGB|397379005|SNOMEDCT_US|Pineal parenchymal tumour of intermediate differentiation|9362/3
C1367859|T191|SYGB|31671006|SNOMEDCT_US|Pineal parenchymal tumour of intermediate differentiation|9362/3
C0205898|T191|PT|767448007|SNOMEDCT_US|Pineoblastoma|9362/3
C0205898|T191|PT|31671006|SNOMEDCT_US|Pineoblastoma|9362/3
C0206094|T191|SY|0000020806|CHV|melanoameloblastoma|9363/0
C0206094|T191|PT|0000020806|CHV|melanotic neuroectodermal tumor|9363/0
C0206094|T191|SY|0000020806|CHV|melanotic neuroectodermal tumour|9363/0
C0206094|T191|PM|D017600|MSH|Anlage Tumor, Retinal|9363/0
C0206094|T191|PM|D017600|MSH|Anlage Tumors, Retinal|9363/0
C0206094|T191|ET|D017600|MSH|Melanoameloblastoma|9363/0
C0206094|T191|PM|D017600|MSH|Melanoameloblastomas|9363/0
C0206094|T191|PM|D017600|MSH|Melanotic Neuroectodermal Tumor|9363/0
C0206094|T191|PM|D017600|MSH|Melanotic Neuroectodermal Tumors|9363/0
C0206094|T191|PM|D017600|MSH|Melanotic Progonoma|9363/0
C0206094|T191|PM|D017600|MSH|Melanotic Progonomas|9363/0
C0206094|T191|MH|D017600|MSH|Neuroectodermal Tumor, Melanotic|9363/0
C0206094|T191|PM|D017600|MSH|Neuroectodermal Tumors, Melanotic|9363/0
C0206094|T191|ET|D017600|MSH|Progonoma, Melanotic|9363/0
C0206094|T191|PM|D017600|MSH|Progonomas, Melanotic|9363/0
C0206094|T191|ET|D017600|MSH|Retinal Anlage Tumor|9363/0
C0206094|T191|PM|D017600|MSH|Retinal Anlage Tumors|9363/0
C0206094|T191|PM|D017600|MSH|Tumor, Melanotic Neuroectodermal|9363/0
C0206094|T191|PM|D017600|MSH|Tumor, Retinal Anlage|9363/0
C0206094|T191|PM|D017600|MSH|Tumors, Melanotic Neuroectodermal|9363/0
C0206094|T191|PM|D017600|MSH|Tumors, Retinal Anlage|9363/0
C0206094|T191|SY|C3717|NCI|Infantile Melanotic Neuroectodermal Neoplasm|9363/0
C0206094|T191|PT|C3717|NCI|Melanotic Neuroectodermal Tumor|9363/0
C0206094|T191|SY|C3717|NCI|Melanotic Neuroectodermal Tumor of Infancy|9363/0
C0206094|T191|SY|C3717|NCI|Melanotic Progonoma|9363/0
C0206094|T191|AB|C3717|NCI|MNTI|9363/0
C0206094|T191|SY|C3717|NCI|Pigmented Neuroectodermal Tumor|9363/0
C0206094|T191|SY|C3717|NCI|Retinal Anlage Neoplasm|9363/0
C0206094|T191|SY|BBa4.|RCD|Melanomeloblastoma|9363/0
C0206094|T191|AB|BBa4.|RCD|Melanotic neuroectodermal tum|9363/0
C0206094|T191|PT|BBa4.|RCD|Melanotic neuroectodermal tumour|9363/0
C0206094|T191|PT|X77pb|RCD|Melanotic neuroectodermal tumour of infancy|9363/0
C0206094|T191|SY|BBa4.|RCD|Melanotic progonoma|9363/0
C0206094|T191|SY|X77pb|RCD|Melanotic progonoma of skin|9363/0
C0206094|T191|AB|X77pb|RCD|Primi neuroectoderm tum infan|9363/0
C0206094|T191|SY|BBa4.|RCD|Retinal anlage tumour|9363/0
C0206094|T191|PT|BBa4.|RCDAE|Melanotic neuroectodermal tumor|9363/0
C0206094|T191|PT|X77pb|RCDAE|Melanotic neuroectodermal tumor of infancy|9363/0
C0206094|T191|SY|BBa4.|RCDAE|Retinal anlage tumor|9363/0
C0206094|T191|SY|1513001|SNOMEDCT_US|Melanoameloblastoma|9363/0
C0206094|T191|IS|1513001|SNOMEDCT_US|Melanomeloblastoma|9363/0
C0206094|T191|PT|1513001|SNOMEDCT_US|Melanotic neuroectodermal tumor|9363/0
C0206094|T191|OAP|253076000|SNOMEDCT_US|Melanotic neuroectodermal tumor of infancy|9363/0
C0206094|T191|PT|767047005|SNOMEDCT_US|Melanotic neuroectodermal tumor of infancy|9363/0
C0206094|T191|PTGB|1513001|SNOMEDCT_US|Melanotic neuroectodermal tumour|9363/0
C0206094|T191|PTGB|767047005|SNOMEDCT_US|Melanotic neuroectodermal tumour of infancy|9363/0
C0206094|T191|OAP|253076000|SNOMEDCT_US|Melanotic neuroectodermal tumour of infancy|9363/0
C0206094|T191|SY|404042005|SNOMEDCT_US|Melanotic progonoma|9363/0
C0206094|T191|SY|1513001|SNOMEDCT_US|Melanotic progonoma|9363/0
C0206094|T191|OAS|253076000|SNOMEDCT_US|Melanotic progonoma of skin|9363/0
C0206094|T191|SY|767047005|SNOMEDCT_US|MNTI - melanotic neuroectodermal tumor of infancy|9363/0
C0206094|T191|SYGB|767047005|SNOMEDCT_US|MNTI - melanotic neuroectodermal tumour of infancy|9363/0
C0206094|T191|SYGB|767047005|SNOMEDCT_US|MNTI-melanotic neuroectodermal tumour of infancy|9363/0
C0206094|T191|PT|404042005|SNOMEDCT_US|Pigmented neuroectodermal tumor of infancy|9363/0
C0206094|T191|PTGB|404042005|SNOMEDCT_US|Pigmented neuroectodermal tumour of infancy|9363/0
C0206094|T191|SY|404042005|SNOMEDCT_US|Retinal anlage tumor|9363/0
C0206094|T191|SY|1513001|SNOMEDCT_US|Retinal anlage tumor|9363/0
C0206094|T191|SYGB|404042005|SNOMEDCT_US|Retinal anlage tumour|9363/0
C0206094|T191|SYGB|1513001|SNOMEDCT_US|Retinal anlage tumour|9363/0
C0553580|T191|SY|0000039089|CHV|ewing sarcoma|9364/3
C0553580|T191|SY|0000039089|CHV|ewing tumor|9364/3
C0684337|T191|PT|0000043998|CHV|Ewing tumor of bone|9364/3
C0553580|T191|PT|0000039089|CHV|ewing's sarcoma|9364/3
C0553580|T191|SY|0000039089|CHV|ewing's tumor|9364/3
C0553580|T191|SY|0000039089|CHV|ewing's tumors|9364/3
C0553580|T191|SY|0000039089|CHV|ewings sarcoma|9364/3
C0553580|T191|SY|0000039089|CHV|ewings tumor|9364/3
C0553580|T191|SY|0000039089|CHV|ewings tumors|9364/3
C0553580|T191|SY|0000039089|CHV|ewings's sarcoma|9364/3
C0684337|T191|SY|0000043998|CHV|peripheral neuroectodermal tumor|9364/3
C0684337|T191|SY|0000043998|CHV|pnet|9364/3
C0553580|T191|SY|0000039089|CHV|sarcoma ewing|9364/3
C0553580|T191|SY|0000039089|CHV|sarcoma ewing's|9364/3
C0553580|T191|SY|0000039089|CHV|sarcoma ewings|9364/3
C0553580|T191|PT|NOCODE|COSTAR|Ewing's Sarcoma|9364/3
C0553580|T191|ET|2008-4746|CSP|Ewing's sarcoma|9364/3
C0553580|T191|PT|2008-4746|CSP|Ewing's tumor|9364/3
C0553580|T191|SY|NOCODE|DXP|EWING TUMOR|9364/3
C0553580|T191|DI|U001700|DXP|SARCOMA, EWING|9364/3
C0553580|T191|PT|HP:0012254|HPO|Ewing sarcoma|9364/3
C0553580|T191|SY|HP:0012254|HPO|Ewing sarcoma|9364/3
C0553580|T191|SY|HP:0012254|HPO|Ewing's sarcoma|9364/3
C0684337|T191|PT|HP:0030067|HPO|Peripheral primitive neuroectodermal neoplasm|9364/3
C0553580|T191|PT|sh85046050|LCH_NW|Ewing's sarcoma|9364/3
C0553580|T191|LLT|10015560|MDR|Ewing's sarcoma|9364/3
C0553580|T191|PT|10015560|MDR|Ewing's sarcoma|9364/3
C0553580|T191|LLT|10015563|MDR|Ewing's sarcoma NOS|9364/3
C0553580|T191|LLT|10015565|MDR|Ewing's sarcoma stage unspecified|9364/3
C0553580|T191|LLT|10015566|MDR|Ewing's tumor|9364/3
C0553580|T191|LLT|10015570|MDR|Ewing's tumour|9364/3
C0684337|T191|SY|354546|MEDCIN|malignant neoplasm primary peripheral neuroectodermal tumor|9364/3
C0684337|T191|PT|354546|MEDCIN|peripheral neuroectodermal tumor|9364/3
C0553580|T191|ET|169|MEDLINEPLUS|Ewing's Sarcoma|9364/3
C0553580|T191|ET|169|MEDLINEPLUS|Sarcoma, Ewing's|9364/3
C0553580|T191|ET|D012512|MSH|Ewing Sarcoma|9364/3
C0553580|T191|ET|D012512|MSH|Ewing Tumor|9364/3
C0553580|T191|ET|D012512|MSH|Ewing's Sarcoma|9364/3
C0553580|T191|ET|D012512|MSH|Ewing's Tumor|9364/3
C0553580|T191|PM|D012512|MSH|Ewings Sarcoma|9364/3
C0553580|T191|PM|D012512|MSH|Ewings Tumor|9364/3
C0684337|T191|ET|D018241|MSH|Extracranial Primitive Neuroectodermal Tumor|9364/3
C0684337|T191|DEV|D018241|MSH|NEUROECTODERMAL NEOPL PERIPHERAL PRIMITIVE|9364/3
C0684337|T191|ET|D018241|MSH|Neuroectodermal Neoplasm, Peripheral Primitive|9364/3
C0684337|T191|ET|D018241|MSH|Neuroectodermal Tumor, Peripheral|9364/3
C0684337|T191|ET|D018241|MSH|Neuroectodermal Tumor, Peripheral Primitive|9364/3
C0684337|T191|PM|D018241|MSH|Neuroectodermal Tumors, Peripheral|9364/3
C0684337|T191|MH|D018241|MSH|Neuroectodermal Tumors, Primitive, Peripheral|9364/3
C0684337|T191|ET|D018241|MSH|Neuroepithelioma, Peripheral|9364/3
C0684337|T191|PM|D018241|MSH|Neuroepitheliomas, Peripheral|9364/3
C0684337|T191|PM|D018241|MSH|Peripheral Neuroectodermal Tumor|9364/3
C0684337|T191|PM|D018241|MSH|Peripheral Neuroectodermal Tumors|9364/3
C0684337|T191|PM|D018241|MSH|Peripheral Neuroepithelioma|9364/3
C0684337|T191|PM|D018241|MSH|Peripheral Neuroepitheliomas|9364/3
C0684337|T191|DEV|D018241|MSH|PERIPHERAL PRIMITIVE NEUROECTODERMAL NEOPL|9364/3
C0684337|T191|ET|D018241|MSH|Peripheral Primitive Neuroectodermal Neoplasm|9364/3
C0684337|T191|ET|D018241|MSH|Peripheral Primitive Neuroectodermal Tumors|9364/3
C0684337|T191|ET|D018241|MSH|Primitive Neuroectodermal Tumor, Extracranial|9364/3
C0553580|T191|MH|D012512|MSH|Sarcoma, Ewing|9364/3
C0553580|T191|ET|D012512|MSH|Sarcoma, Ewing's|9364/3
C0553580|T191|PM|D012512|MSH|Sarcoma, Ewings|9364/3
C0553580|T191|PM|D012512|MSH|Tumor, Ewing|9364/3
C0553580|T191|PM|D012512|MSH|Tumor, Ewing's|9364/3
C0684337|T191|PM|D018241|MSH|Tumor, Peripheral Neuroectodermal|9364/3
C0684337|T191|PM|D018241|MSH|Tumors, Peripheral Neuroectodermal|9364/3
C0553580|T191|PN|NOCODE|MTH|Ewings sarcoma|9364/3
C0553580|T191|SY|C4817|NCI|ES|9364/3
C0553580|T191|PT|C4817|NCI|Ewing Sarcoma|9364/3
C0553580|T191|SY|C4817|NCI|Ewing's Sarcoma|9364/3
C0553580|T191|SY|C4817|NCI|Ewing's Tumor|9364/3
C0684337|T191|SY|C9341|NCI|Peripheral Neuroectodermal Neoplasm|9364/3
C0684337|T191|SY|C9341|NCI|Peripheral Neuroectodermal Tumor|9364/3
C0684337|T191|SY|C9341|NCI|Peripheral Neuroepithelioma|9364/3
C0684337|T191|SY|C9341|NCI|Peripheral PNET|9364/3
C0684337|T191|SY|C9341|NCI|Peripheral Primitive Neuroectodermal Neoplasm|9364/3
C0684337|T191|PT|C9341|NCI|Peripheral Primitive Neuroectodermal Tumor|9364/3
C0684337|T191|AB|C9341|NCI|pPNET|9364/3
C0553580|T191|PT|C4817|NCI_CPTAC|Ewing Sarcoma|9364/3
C0553580|T191|DN|C4817|NCI_CTRP|Ewing Sarcoma|9364/3
C0553580|T191|PT|C4817|NCI_CTRP|Ewing Sarcoma|9364/3
C0684337|T191|DN|C9341|NCI_CTRP|Peripheral Primitive Neuroectodermal Tumor|9364/3
C0553580|T191|PT|CDR0000046031|NCI_NCI-GLOSS|Ewing sarcoma|9364/3
C0684337|T191|PT|CDR0000045848|NCI_NCI-GLOSS|peripheral primitive neuroectodermal tumor|9364/3
C0684337|T191|PT|CDR0000520410|NCI_NCI-GLOSS|pPNET|9364/3
C0553580|T191|PT|C4817|NCI_NICHD|Ewing Sarcoma|9364/3
C0553580|T191|PT|CDR0000546979|PDQ|Ewing sarcoma|9364/3
C0684337|T191|ET|CDR0000039466|PDQ|Ewing sarcoma/PNET|9364/3
C0684337|T191|OP|CDR0000043409|PDQ|Ewing's family of tumors|9364/3
C0684337|T191|SY|CDR0000039466|PDQ|Ewing's family of tumors|9364/3
C0553580|T191|SY|CDR0000546979|PDQ|Ewing's Sarcoma|9364/3
C0553580|T191|SY|CDR0000546979|PDQ|Ewing's Tumor|9364/3
C0684337|T191|SY|CDR0000546986|PDQ|Peripheral Neuroectodermal Neoplasm|9364/3
C0684337|T191|SY|CDR0000546986|PDQ|Peripheral Neuroectodermal Tumor|9364/3
C0684337|T191|SY|CDR0000039466|PDQ|peripheral neuroectodermal tumor|9364/3
C0684337|T191|SY|CDR0000546986|PDQ|Peripheral Neuroepithelioma|9364/3
C0684337|T191|SY|CDR0000546986|PDQ|Peripheral PNET|9364/3
C0684337|T191|SY|CDR0000546986|PDQ|Peripheral Primitive Neuroectodermal Neoplasm|9364/3
C0684337|T191|PT|CDR0000546986|PDQ|peripheral primitive neuroectodermal tumor|9364/3
C0684337|T191|SY|CDR0000546986|PDQ|Peripheral Primitive Neuroectodermal Tumors|9364/3
C0684337|T191|SY|CDR0000039466|PDQ|pPNET|9364/3
C0684337|T191|AB|CDR0000546986|PDQ|pPNET|9364/3
C0684337|T191|SY|CDR0000039466|PDQ|primitive neuroectodermal tumor, peripheral|9364/3
C0684337|T191|SY|CDR0000039466|PDQ|primitive peripheral neuroectodermal tumor|9364/3
C0684337|T191|SY|CDR0000039466|PDQ|sarcoma, Ewing's|9364/3
C0553580|T191|PT|BBY0.|RCD|Ewing's sarcoma|9364/3
C0553580|T191|SY|BBY0.|RCD|Ewing's tumour|9364/3
C0684337|T191|AB|X77q4|RCD|Peripheral neuroectodermal tum|9364/3
C0684337|T191|PT|X77q4|RCD|Peripheral neuroectodermal tumour|9364/3
C0553580|T191|SY|BBY0.|RCDAE|Ewing's tumor|9364/3
C0684337|T191|PT|X77q4|RCDAE|Peripheral neuroectodermal tumor|9364/3
C0553580|T191|SY|76909002|SNOMEDCT_US|Ewing sarcoma|9364/3
C0684337|T191|PT|703707001|SNOMEDCT_US|Ewing sarcoma / peripheral neuroectodermal tumor|9364/3
C0684337|T191|PTGB|703707001|SNOMEDCT_US|Ewing sarcoma / peripheral neuroectodermal tumour|9364/3
C0684337|T191|SY|703707001|SNOMEDCT_US|Ewing sarcoma / PNET|9364/3
C0553580|T191|PT|76909002|SNOMEDCT_US|Ewing's sarcoma|9364/3
C0553580|T191|SY|76909002|SNOMEDCT_US|Ewing's tumor|9364/3
C0553580|T191|SYGB|76909002|SNOMEDCT_US|Ewing's tumour|9364/3
C0684337|T191|PT|73676002|SNOMEDCT_US|Peripheral neuroectodermal tumor|9364/3
C0684337|T191|PT|253096008|SNOMEDCT_US|Peripheral neuroectodermal tumor|9364/3
C0684337|T191|PTGB|73676002|SNOMEDCT_US|Peripheral neuroectodermal tumour|9364/3
C0684337|T191|PTGB|253096008|SNOMEDCT_US|Peripheral neuroectodermal tumour|9364/3
C0684337|T191|SY|73676002|SNOMEDCT_US|Peripheral primitive neuroectodermal tumor|9364/3
C0684337|T191|SYGB|73676002|SNOMEDCT_US|Peripheral primitive neuroectodermal tumour|9364/3
C0684337|T191|SY|73676002|SNOMEDCT_US|PPNET|9364/3
C0877849|T191|SY|0000051935|CHV|askin tumor|9365/3
C0877849|T191|PT|0000051935|CHV|askin's tumor|9365/3
C0877849|T191|SY|0000051935|CHV|askin's tumors|9365/3
C0877849|T191|LLT|10057657|MDR|Askin's tumor|9365/3
C0877849|T191|LLT|10057656|MDR|Askin's tumour|9365/3
C0877849|T191|NM|C563168|MSH|Askin Tumor|9365/3
C0877849|T191|PN|NOCODE|MTH|Askin's tumor|9365/3
C0877849|T191|PT|C7542|NCI|Askin Tumor|9365/3
C0877849|T191|SY|C7542|NCI|Askin's Tumor|9365/3
C0877849|T191|SY|C7542|NCI|Peripheral Neuroectodermal Tumor of Thoracopulmonary Region|9365/3
C0877849|T191|SY|C7542|NCI|PNET of Thoracopulmonary Region|9365/3
C0877849|T191|SY|C7542|NCI|Small Cell Tumor of Thoracopulmonary Region|9365/3
C0877849|T191|DN|C7542|NCI_CTRP|Askin Tumor|9365/3
C0877849|T191|PT|CDR0000546988|PDQ|Askin tumor|9365/3
C0877849|T191|SY|CDR0000546988|PDQ|Askin's Tumor|9365/3
C0877849|T191|SY|CDR0000546988|PDQ|Peripheral Neuroectodermal Tumor of Thoracopulmonary Region|9365/3
C0877849|T191|SY|CDR0000546988|PDQ|PNET of chest wall|9365/3
C0877849|T191|SY|CDR0000546988|PDQ|PNET of Thoracopulmonary Region|9365/3
C0877849|T191|SY|CDR0000546988|PDQ|Small Cell Tumor of Thoracopulmonary Region|9365/3
C0877849|T191|PT|X77oU|RCD|Askin's tumour|9365/3
C0877849|T191|PT|X77oU|RCDAE|Askin's tumor|9365/3
C0877849|T191|IS|128783001|SNOMEDCT_US|Askin tumor|9365/3
C0877849|T191|PT|128783001|SNOMEDCT_US|Askin tumor|9365/3
C0877849|T191|PTGB|128783001|SNOMEDCT_US|Askin tumour|9365/3
C0877849|T191|IS|73506006|SNOMEDCT_US|Askin's tumor|9365/3
C0877849|T191|OAP|134210007|SNOMEDCT_US|Askin's tumor|9365/3
C0877849|T191|SY|128783001|SNOMEDCT_US|Askin's tumor|9365/3
C0877849|T191|OAP|134210007|SNOMEDCT_US|Askin's tumour|9365/3
C0877849|T191|SYGB|128783001|SNOMEDCT_US|Askin's tumour|9365/3
C3839583|T191|PT|703708006|SNOMEDCT_US|Benign notochordal tumor|9370/0
C3839583|T191|PTGB|703708006|SNOMEDCT_US|Benign notochordal tumour|9370/0
C0008487|T191|PT|0000002906|CHV|chordoma|9370/3
C0008487|T191|SY|0000002906|CHV|chordomas|9370/3
C0008487|T191|PT|2000-4323|CSP|chordoma|9370/3
C0008487|T191|ET|2000-4323|CSP|notochordoma|9370/3
C0008487|T191|PT|HP:0010762|HPO|Chordoma|9370/3
C0008487|T191|PT|U000997|LCH|Chordoma|9370/3
C0008487|T191|PT|sh85024739|LCH_NW|Chordoma|9370/3
C0008487|T191|PT|10008747|MDR|Chordoma|9370/3
C0008487|T191|LLT|10008747|MDR|Chordoma|9370/3
C0008487|T191|PT|271560|MEDCIN|chordoma|9370/3
C0008487|T191|MH|D002817|MSH|Chordoma|9370/3
C0008487|T191|PM|D002817|MSH|Chordomas|9370/3
C0008487|T191|PT|C2947|NCI|Chordoma|9370/3
C0008487|T191|PT|C2947|NCI_CDISC|CHORDOMA, MALIGNANT|9370/3
C0008487|T191|PT|C2947|NCI_CPTAC|Chordoma|9370/3
C0008487|T191|DN|C2947|NCI_CTRP|Chordoma|9370/3
C0008487|T191|PT|C2947|NCI_CTRP|Chordoma|9370/3
C0008487|T191|PT|CDR0000045297|NCI_NCI-GLOSS|chordoma|9370/3
C0008487|T191|PSC|CDR0000040402|PDQ|chordoma|9370/3
C0008487|T191|ET|CDR0000040402|PDQ|Chordoma|9370/3
C0008487|T191|PT|BBa5.|RCD|Chordoma|9370/3
C0008487|T191|PT|50007008|SNOMEDCT_US|Chordoma|9370/3
C1266173|T191|PT|271561|MEDCIN|chondroid chordoma|9371/3
C1266173|T191|PT|C6902|NCI|Chondroid Chordoma|9371/3
C1266173|T191|PT|128784007|SNOMEDCT_US|Chondroid chordoma|9371/3
C1266174|T191|PT|271562|MEDCIN|dedifferentiated chordoma|9372/3
C1266174|T191|PT|C48876|NCI|Dedifferentiated Chordoma|9372/3
C1266174|T191|SY|C48876|NCI|Sarcomatoid Chordoma|9372/3
C1266174|T191|PT|128785008|SNOMEDCT_US|Dedifferentiated chordoma|9372/3
C1266175|T191|PT|C6581|NCI|Parachordoma|9373/0
C1266175|T191|PT|128786009|SNOMEDCT_US|Parachordoma|9373/0
C1266175|T191|PT|404086000|SNOMEDCT_US|Parachordoma|9373/0
C1266175|T191|PT|C6581|NCI|Parachordoma|9373/1
C1266175|T191|PT|404086000|SNOMEDCT_US|Parachordoma|9373/1
C1266175|T191|PT|128786009|SNOMEDCT_US|Parachordoma|9373/1
C0555198|T191|PT|0000039208|CHV|malignant glioma|9380/3
C0555198|T191|SY|0000039208|CHV|malignant gliomas|9380/3
C0555198|T191|MTH_HT|10018335|MDR|Glial tumors malignant|9380/3
C0555198|T191|HT|10018335|MDR|Glial tumours malignant|9380/3
C0555198|T191|PT|10065443|MDR|Malignant glioma|9380/3
C0555198|T191|LLT|10065443|MDR|Malignant glioma|9380/3
C0555198|T191|PM|D005910|MSH|Glioma, Malignant|9380/3
C0555198|T191|PM|D005910|MSH|Gliomas, Malignant|9380/3
C0555198|T191|PEP|D005910|MSH|Malignant Glioma|9380/3
C0555198|T191|PM|D005910|MSH|Malignant Gliomas|9380/3
C4722099|T191|PN|NOCODE|MTH|High grade glioma|9380/3
C0555198|T191|PN|NOCODE|MTH|Malignant Glioma|9380/3
C4289688|T191|PT|C129309|NCI|Diffuse Midline Glioma, H3 K27M-Mutant|9380/3
C0555198|T191|SY|C4822|NCI|High Grade Glioma|9380/3
C0555198|T191|SY|C4822|NCI|High-Grade Glioma|9380/3
C0555198|T191|SY|C4822|NCI|Malignant Glial Neoplasm|9380/3
C0555198|T191|SY|C4822|NCI|Malignant Glial Tumor|9380/3
C0555198|T191|PT|C4822|NCI|Malignant Glioma|9380/3
C0555198|T191|SY|C4822|NCI|Malignant Neuroglial Neoplasm|9380/3
C0555198|T191|SY|C4822|NCI|Malignant Neuroglial Tumor|9380/3
C0555198|T191|PT|C4822|NCI_CDISC|GLIOMA, MALIGNANT|9380/3
C0555198|T191|SY|C4822|NCI_CDISC|Malignant Glial Neoplasm|9380/3
C0555198|T191|SY|C4822|NCI_CDISC|Malignant Glial Tumor|9380/3
C0555198|T191|SY|C4822|NCI_CDISC|Malignant Neuroglial Neoplasm|9380/3
C0555198|T191|SY|C4822|NCI_CDISC|Malignant Neuroglial Tumor|9380/3
C0555198|T191|PT|C4822|NCI_CTRP|Malignant Glioma|9380/3
C0555198|T191|DN|C4822|NCI_CTRP|Malignant Glioma|9380/3
C0555198|T191|OP|XE1wa|RCD|Malignant glioma|9380/3
C4289688|T191|SY|733862004|SNOMEDCT_US|Diffuse midline glioma, H3 K27M-mutant|9380/3
C4289688|T191|PT|733862004|SNOMEDCT_US|Diffuse midline glioma, point mutation K27M in histone H3|9380/3
C4518387|T191|PT|734093008|SNOMEDCT_US|Embryonal neoplasm with multilayered rosettes|9380/3
C4518388|T191|PT|734087000|SNOMEDCT_US|Embryonal neoplasm with multilayered rosettes with C19MC-altered|9380/3
C0555198|T191|SY|74532006|SNOMEDCT_US|Glioma, malignant|9380/3
C0555198|T191|PT|74532006|SNOMEDCT_US|Glioma, malignant, no ICD-O subtype|9380/3
C4722099|T191|PT|772292003|SNOMEDCT_US|High grade glioma|9380/3
C4722099|T191|SY|772292003|SNOMEDCT_US|High-grade glioma|9380/3
C0555198|T191|OAP|269505000|SNOMEDCT_US|Malignant glioma|9380/3
C0555198|T191|SY|74532006|SNOMEDCT_US|Malignant glioma|9380/3
C0555198|T191|PT|416500007|SNOMEDCT_US|Malignant glioma - category|9380/3
C0334576|T191|PT|MTHU032165|ICPC2ICD10ENG|gliomatosis; cerebri|9381/3
C0334576|T191|PT|10066254|MDR|Gliomatosis cerebri|9381/3
C0334576|T191|LLT|10066254|MDR|Gliomatosis cerebri|9381/3
C0334576|T191|PEP|D018302|MSH|Gliomatosis Cerebri|9381/3
C0334576|T191|PN|NOCODE|MTH|Gliomatosis cerebri|9381/3
C0334576|T191|SY|C4318|NCI|Astrocytosis cerebri|9381/3
C0334576|T191|SY|C4318|NCI|Gliomatosis|9381/3
C0334576|T191|PT|C4318|NCI|Gliomatosis Cerebri|9381/3
C0334576|T191|PT|BBb1.|RCD|Gliomatosis cerebri|9381/3
C0334576|T191|PT|26138003|SNOMEDCT_US|Gliomatosis cerebri|9381/3
C0431108|T191|SY|0000034148|CHV|anaplastic oligoastrocytoma|9382/3
C0259783|T191|SY|0000025233|CHV|glial mixed tumor|9382/3
C0259783|T191|PT|0000025233|CHV|mixed glioma|9382/3
C0547065|T191|SY|0000038901|CHV|mixed oligo-astrocytoma|9382/3
C0547065|T191|PT|0000038901|CHV|mixed oligoastrocytoma|9382/3
C0259783|T191|LLT|10074669|MDR|Mixed glioma|9382/3
C0547065|T191|LLT|10027769|MDR|Mixed oligo-astrocytoma|9382/3
C0259783|T191|PT|351510|MEDCIN|mixed glioma|9382/3
C0259783|T191|PM|D005910|MSH|Glioma, Mixed|9382/3
C0259783|T191|PM|D005910|MSH|Gliomas, Mixed|9382/3
C0259783|T191|PEP|D005910|MSH|Mixed Glioma|9382/3
C0259783|T191|PM|D005910|MSH|Mixed Gliomas|9382/3
C0547065|T191|PM|D001254|MSH|Mixed Oligoastrocytoma|9382/3
C0547065|T191|PM|D001254|MSH|Mixed Oligoastrocytomas|9382/3
C0547065|T191|PEP|D001254|MSH|Oligoastrocytoma, Mixed|9382/3
C0547065|T191|PM|D001254|MSH|Oligoastrocytomas, Mixed|9382/3
C0431108|T191|PN|NOCODE|MTH|Anaplastic Oligoastrocytoma|9382/3
C0259783|T191|PN|NOCODE|MTH|mixed gliomas|9382/3
C0547065|T191|PN|NOCODE|MTH|Mixed oligoastrocytoma|9382/3
C0431108|T191|SY|C6959|NCI|Anaplastic Mixed Glioma|9382/3
C0431108|T191|SY|TCGA|NCI|Anaplastic Oligoastrocytoma|9382/3
C0431108|T191|PT|C6959|NCI|Anaplastic Oligoastrocytoma|9382/3
C0431108|T191|SY|C129324|NCI|Anaplastic Oligoastrocytoma, NOS|9382/3
C0431108|T191|PT|C129324|NCI|Anaplastic Oligoastrocytoma, Not Otherwise Specified|9382/3
C0259783|T191|SY|C3903|NCI|Mixed Glial Neoplasm|9382/3
C0259783|T191|SY|C3903|NCI|Mixed Glial Tumor|9382/3
C0259783|T191|PT|C3903|NCI|Mixed Glioma|9382/3
C0259783|T191|SY|C3903|NCI|Mixed Neuroglial Neoplasm|9382/3
C0259783|T191|SY|C3903|NCI|Mixed Neuroglial Tumor|9382/3
C0431108|T191|SY|C6959|NCI|WHO Grade III Mixed Glioma|9382/3
C0259783|T191|SY|C3903|NCI_CDISC|Glioma, Mixed|9382/3
C0259783|T191|PT|C3903|NCI_CDISC|GLIOMA, MIXED, MALIGNANT|9382/3
C0259783|T191|SY|C3903|NCI_CDISC|Mixed Glial Neoplasm|9382/3
C0259783|T191|SY|C3903|NCI_CDISC|Mixed Glial Tumor|9382/3
C0259783|T191|SY|C3903|NCI_CDISC|Mixed Neuroglial Neoplasm|9382/3
C0259783|T191|SY|C3903|NCI_CDISC|Mixed Neuroglial Tumor|9382/3
C0431108|T191|PT|C6959|NCI_CPTAC|Anaplastic Oligoastrocytoma|9382/3
C0431108|T191|PT|C129324|NCI_CPTAC|Anaplastic Oligoastrocytoma, NOS|9382/3
C0259783|T191|PT|C3903|NCI_CTRP|Mixed Glioma|9382/3
C0259783|T191|DN|C3903|NCI_CTRP|Mixed Glioma|9382/3
C0259783|T191|PT|CDR0000045344|NCI_NCI-GLOSS|mixed glioma|9382/3
C0431108|T191|PT|X77pT|RCD|Anaplastic oligoastrocytoma|9382/3
C0259783|T191|PT|BBb2.|RCD|Mixed glioma|9382/3
C0547065|T191|PT|X77pS|RCD|Mixed oligoastrocytoma|9382/3
C0431108|T191|PT|253072003|SNOMEDCT_US|Anaplastic oligoastrocytoma|9382/3
C0431108|T191|SY|22217002|SNOMEDCT_US|Anaplastic oligoastrocytoma|9382/3
C0259783|T191|PT|443937008|SNOMEDCT_US|Mixed glioma|9382/3
C0259783|T191|PT|22217002|SNOMEDCT_US|Mixed glioma|9382/3
C0547065|T191|PT|716647001|SNOMEDCT_US|Mixed oligoastrocytoma|9382/3
C0547065|T191|PT|253071005|SNOMEDCT_US|Mixed oligoastrocytoma|9382/3
C0547065|T191|IS|22217002|SNOMEDCT_US|Mixed oligoastrocytoma|9382/3
C0206725|T191|SY|0000021049|CHV|astrocytoma subependymal|9383/1
C0206725|T191|SY|0000021049|CHV|subependymal astrocytoma|9383/1
C0206725|T191|SY|0000021049|CHV|subependymal glioma|9383/1
C0206725|T191|PT|0000021049|CHV|subependymoma|9383/1
C0206725|T191|PT|MTHU008890|ICPC2ICD10ENG|astrocytoma; subependymal|9383/1
C0206725|T191|PT|MTHU071276|ICPC2ICD10ENG|subependymal; astrocytoma|9383/1
C0206725|T191|PM|D018315|MSH|Astrocytoma, Subependymal|9383/1
C0206725|T191|PM|D018315|MSH|Astrocytomas, Subependymal|9383/1
C0206725|T191|MH|D018315|MSH|Glioma, Subependymal|9383/1
C0206725|T191|PM|D018315|MSH|Gliomas, Subependymal|9383/1
C0206725|T191|ET|D018315|MSH|Subependymal Astrocytoma|9383/1
C0206725|T191|PM|D018315|MSH|Subependymal Astrocytomas|9383/1
C0206725|T191|ET|D018315|MSH|Subependymal Glioma|9383/1
C0206725|T191|PM|D018315|MSH|Subependymal Gliomas|9383/1
C0206725|T191|ET|D018315|MSH|Subependymoma|9383/1
C0206725|T191|PM|D018315|MSH|Subependymomas|9383/1
C0206725|T191|PN|NOCODE|MTH|Subependymal Glioma|9383/1
C0206725|T191|SY|C3795|NCI|Subependymal Astrocytoma|9383/1
C0206725|T191|SY|C3795|NCI|Subependymal Glioma|9383/1
C0206725|T191|SY|TCGA|NCI|Subependymoma|9383/1
C0206725|T191|PT|C3795|NCI|Subependymoma|9383/1
C0206725|T191|SY|C3795|NCI|WHO Grade I Ependymal Neoplasm|9383/1
C0206725|T191|SY|C3795|NCI|WHO Grade I Ependymal Tumor|9383/1
C0206725|T191|SY|C3795|NCI_CDISC|Subependymal Glioma|9383/1
C0206725|T191|PT|C3795|NCI_CDISC|SUBEPENDYMOMA, BENIGN|9383/1
C0206725|T191|SY|C3795|NCI_CDISC|Who Grade I Ependymal Neoplasm|9383/1
C0206725|T191|SY|C3795|NCI_CDISC|Who Grade I Ependymal Tumor|9383/1
C0206725|T191|IS|Xa07D|RCD|Subependymoma|9383/1
C0206725|T191|OP|Xa07D|RCDSY|Subependymal astrocytoma NOS|9383/1
C0206725|T191|OA|Xa07D|RCDSY|Subependyml astrocytoma NOS|9383/1
C0206725|T191|SY|4553004|SNOMEDCT_US|Mixed subependymoma-ependymoma|9383/1
C0206725|T191|SY|4553004|SNOMEDCT_US|Subependymal astrocytoma|9383/1
C0206725|T191|IS|4553004|SNOMEDCT_US|Subependymal astrocytoma, NOS|9383/1
C0206725|T191|PT|4553004|SNOMEDCT_US|Subependymal glioma|9383/1
C0206725|T191|SY|4553004|SNOMEDCT_US|Subependymoma|9383/1
C0205768|T191|PT|HP:0009718|HPO|Subependymal giant-cell astrocytoma|9384/1
C0205768|T191|LLT|10073233|MDR|Subependymal giant cell astrocytoma|9384/1
C0205768|T191|SY|31903|MEDCIN|CNS mass lesions ventricle subependymal giant cell astrocytoma|9384/1
C0205768|T191|PT|31903|MEDCIN|subependymal giant cell astrocytoma|9384/1
C0205768|T191|PEP|D001254|MSH|Astrocytoma, Subependymal Giant Cell|9384/1
C0205768|T191|ET|D001254|MSH|Subependymal Giant Cell Astrocytoma|9384/1
C0205768|T191|PN|NOCODE|MTH|Subependymal Giant Cell Astrocytoma|9384/1
C0205768|T191|SY|C3696|NCI|SEGA|9384/1
C0205768|T191|SY|C3696|NCI|Subependymal Giant Cell Astrocytic Neoplasm|9384/1
C0205768|T191|SY|C3696|NCI|Subependymal Giant Cell Astrocytic Tumor|9384/1
C0205768|T191|PT|C3696|NCI|Subependymal Giant Cell Astrocytoma|9384/1
C0205768|T191|AB|BBb4.|RCD|Subepend giant cell astrocytom|9384/1
C0205768|T191|SY|BBb4.|RCD|Subependymal giant cell astrocytoma|9384/1
C0205768|T191|AB|BBb4.|RCDSY|Subepend.giant astrocytoma|9384/1
C0205768|T191|SY|449799008|SNOMEDCT_US|SEGA - Subependymal giant cell astrocytoma|9384/1
C0205768|T191|PT|449799008|SNOMEDCT_US|Subependymal giant cell astrocytoma|9384/1
C0205768|T191|PT|1586004|SNOMEDCT_US|Subependymal giant cell astrocytoma|9384/1
C0205770|T191|PT|0000020713|CHV|choroid plexus papilloma|9390/0
C0205770|T191|SY|0000020713|CHV|choroid plexus papillomas|9390/0
C0205770|T191|SY|NOCODE|DXP|BRAIN TUMOR, CHOROID PLEXUS PAPILLOMA|9390/0
C0205770|T191|DI|U000351|DXP|CHOROID PLEXUS, PAPILLOMA|9390/0
C0205770|T191|SY|NOCODE|DXP|INTRACRANIAL NEOPLASM, CHOROID PLEXUS PAPILLOMA|9390/0
C0205770|T191|PT|HP:0200022|HPO|Choroid plexus papilloma|9390/0
C0205770|T191|PT|MTHU084549|ICPC2ICD10ENG|choroid plexus; papilloma|9390/0
C0205770|T191|PT|MTHU057343|ICPC2ICD10ENG|papilloma; choroid plexus|9390/0
C0205770|T191|PT|MTHU060165|ICPC2ICD10ENG|plexus choroideus; papilloma|9390/0
C0205770|T191|LLT|10008777|MDR|Choroid plexus papilloma|9390/0
C0205770|T191|PT|10008777|MDR|Choroid plexus papilloma|9390/0
C0205770|T191|PT|31929|MEDCIN|papilloma of choroid plexus|9390/0
C0205770|T191|ET|D020288|MSH|Choroid Plexus Papilloma|9390/0
C0205770|T191|PM|D020288|MSH|Choroid Plexus Papillomas|9390/0
C0205770|T191|ET|D020288|MSH|Papilloma of Choroid Plexus|9390/0
C0205770|T191|MH|D020288|MSH|Papilloma, Choroid Plexus|9390/0
C0205770|T191|PM|D020288|MSH|Papillomas, Choroid Plexus|9390/0
C0205770|T191|PN|NOCODE|MTH|Choroid Plexus Papilloma|9390/0
C0205770|T191|SY|TCGA|NCI|Choroid Plexus Papilloma|9390/0
C0205770|T191|PT|C3698|NCI|Choroid Plexus Papilloma|9390/0
C0205770|T191|SY|C3698|NCI|Papilloma of Choroid Plexus|9390/0
C0205770|T191|SY|C3698|NCI|Papilloma of the Choroid Plexus|9390/0
C0205770|T191|SY|C3698|NCI_CDISC|Papilloma of Choroid Plexus|9390/0
C0205770|T191|SY|C3698|NCI_CDISC|Papilloma of the Choroid Plexus|9390/0
C0205770|T191|PT|C3698|NCI_CDISC|PAPILLOMA, CHOROID PLEXUS, BENIGN|9390/0
C0205770|T191|SY|CDR0000043274|PDQ|choroid plexus papilloma|9390/0
C0205770|T191|PT|Xa992|RCD|Choroid plexus papilloma|9390/0
C0205770|T191|OA|BBb5.|RCDSY|Choroid plexus papillom.NOS|9390/0
C0205770|T191|OP|BBb5.|RCDSY|Choroid plexus papilloma NOS|9390/0
C0205770|T191|PT|18021007|SNOMEDCT_US|Choroid plexus papilloma|9390/0
C0205770|T191|SY|18021007|SNOMEDCT_US|Choroid plexus papilloma, no ICD-O subtype|9390/0
C0205770|T191|SY|18021007|SNOMEDCT_US|Choroid plexus papilloma, no International Classification of Diseases for Oncology subtype|9390/0
C0205770|T191|IS|18021007|SNOMEDCT_US|Choroid plexus papilloma, NOS|9390/0
C1266176|T191|PT|C53686|NCI|Atypical Choroid Plexus Papilloma|9390/1
C1266176|T191|PT|128904001|SNOMEDCT_US|Atypical choroid plexus papilloma|9390/1
C0431109|T191|PT|HP:0030392|HPO|Choroid plexus carcinoma|9390/3
C0431109|T191|PT|MTHU005661|ICPC2ICD10ENG|anaplastic; papilloma choroid plexus|9390/3
C0431109|T191|PT|MTHU084548|ICPC2ICD10ENG|choroid plexus; papilloma, anaplastic|9390/3
C0431109|T191|PT|MTHU057344|ICPC2ICD10ENG|papilloma; choroid plexus, anaplastic|9390/3
C0431109|T191|PT|MTHU060166|ICPC2ICD10ENG|plexus choroideus; papilloma, anaplastic|9390/3
C0431109|T191|LLT|10002225|MDR|Anaplastic choroid plexus papilloma|9390/3
C0431109|T191|LLT|10067478|MDR|Choroid plexus carcinoma|9390/3
C0431109|T191|PT|10067478|MDR|Choroid plexus carcinoma|9390/3
C0431109|T191|PT|31930|MEDCIN|carcinoma of choroid plexus|9390/3
C0431109|T191|NM|C562943|MSH|Choroid Plexus Carcinoma|9390/3
C0431109|T191|PN|NOCODE|MTH|Choroid Plexus Carcinoma|9390/3
C0431109|T191|OP|C4715|NCI|Anaplastic Choroid Plexus Papilloma|9390/3
C0431109|T191|SY|C4715|NCI|Cancer of Choroid Plexus|9390/3
C0431109|T191|SY|C4715|NCI|Cancer of the Choroid Plexus|9390/3
C0431109|T191|SY|C4715|NCI|Carcinoma of Choroid Plexus|9390/3
C0431109|T191|SY|C4715|NCI|Carcinoma of the Choroid Plexus|9390/3
C0431109|T191|SY|C4715|NCI|Choroid Plexus Cancer|9390/3
C0431109|T191|PT|C4715|NCI|Choroid Plexus Carcinoma|9390/3
C0431109|T191|SY|TCGA|NCI|Choroid Plexus Carcinoma|9390/3
C0431109|T191|SY|C4715|NCI_CDISC|Anaplastic Choroid Plexus Papilloma|9390/3
C0431109|T191|SY|C4715|NCI_CDISC|Cancer of Choroid Plexus|9390/3
C0431109|T191|SY|C4715|NCI_CDISC|Cancer of the Choroid Plexus|9390/3
C0431109|T191|SY|C4715|NCI_CDISC|Carcinoma of Choroid Plexus|9390/3
C0431109|T191|SY|C4715|NCI_CDISC|Carcinoma of the Choroid Plexus|9390/3
C0431109|T191|PT|C4715|NCI_CDISC|CARCINOMA, CHOROID PLEXUS, MALIGNANT|9390/3
C0431109|T191|SY|C4715|NCI_CDISC|Choroid Plexus Cancer|9390/3
C0431109|T191|PT|C4715|NCI_CPTAC|Choroid Plexus Carcinoma|9390/3
C0431109|T191|PT|90600120|NCI_CTEP-SDC|Choroid plexus carcinoma|9390/3
C0431109|T191|DN|C4715|NCI_CTRP|Choroid Plexus Cancer|9390/3
C0431109|T191|PT|C4715|NCI_CTRP|Choroid Plexus Carcinoma|9390/3
C0431109|T191|SY|CDR0000043274|PDQ|choroid plexus carcinoma|9390/3
C0431109|T191|PT|Xa993|RCD|Choroid plexus carcinoma|9390/3
C0431109|T191|PT|88252006|SNOMEDCT_US|Choroid plexus carcinoma|9390/3
C0431109|T191|SY|88252006|SNOMEDCT_US|Choroid plexus papilloma, anaplastic|9390/3
C0014474|T191|ET|0000004652|AOD|ependymoma|9391/3
C1384403|T191|SY|0000004535|CHV|cellular ependymoma|9391/3
C0014474|T191|PT|0000004535|CHV|ependymoma|9391/3
C0014474|T191|SY|0000004535|CHV|ependymomas|9391/3
C1370500|T191|SY|0000004535|CHV|tanycytic ependymoma|9391/3
C0014474|T191|PT|NOCODE|COSTAR|Ependymoma|9391/3
C0014474|T191|PT|2012-5783|CSP|ependymoma|9391/3
C0014474|T191|PT|HP:0002888|HPO|Ependymoma|9391/3
C0014474|T191|PT|MTHU026460|ICPC2ICD10ENG|ependymoma; unspecified site|9391/3
C0014474|T191|PT|10014967|MDR|Ependymoma|9391/3
C0014474|T191|LLT|10014967|MDR|Ependymoma|9391/3
C1384403|T191|PEP|D004806|MSH|Cellular Ependymoma|9391/3
C1384403|T191|ET|D004806|MSH|Clear Cell Ependymoma|9391/3
C0014474|T191|MH|D004806|MSH|Ependymoma|9391/3
C0014474|T191|PM|D004806|MSH|Ependymomas|9391/3
C1384403|T191|PN|NOCODE|MTH|Cellular Ependymoma|9391/3
C0014474|T191|PN|NOCODE|MTH|Ependymoma|9391/3
C1370500|T191|PN|NOCODE|MTH|Tanycytic ependymoma|9391/3
C1384403|T191|PT|C4713|NCI|Cellular Ependymoma|9391/3
C1384403|T191|PT|C4714|NCI|Clear Cell Ependymoma|9391/3
C0014474|T191|PT|C3017|NCI|Ependymoma|9391/3
C0014474|T191|SY|TCGA|NCI|Ependymoma|9391/3
C4289581|T191|PT|C129351|NCI|Ependymoma, RELA Fusion-Positive|9391/3
C1370500|T191|PT|C6903|NCI|Tanycytic Ependymoma|9391/3
C1370500|T191|SY|TCGA|NCI|Tanycytic Ependymoma|9391/3
C0014474|T191|SY|C3017|NCI|WHO Grade II Ependymal Neoplasm|9391/3
C0014474|T191|SY|C3017|NCI|WHO Grade II Ependymal Tumor|9391/3
C0014474|T191|PT|C3017|NCI_CPTAC|Ependymoma|9391/3
C0014474|T191|PT|10014967|NCI_CTEP-SDC|Ependymoma, NOS|9391/3
C0014474|T191|PT|CDR0000046432|NCI_NCI-GLOSS|ependymoma|9391/3
C0014474|T191|PT|C3017|NCI_NICHD|Ependymoma|9391/3
C1384403|T191|PT|X77pP|RCD|Cellular ependymoma|9391/3
C1384403|T191|PT|X77pQ|RCD|Clear cell ependymoma|9391/3
C0014474|T191|PT|Xa994|RCD|Ependymoma|9391/3
C0014474|T191|OP|X77pO|RCD|Epithelial ependymoma|9391/3
C0014474|T191|OP|BBb7.|RCDSY|Ependymoma NOS|9391/3
C1384403|T191|PT|827053007|SNOMEDCT_US|Cellular ependymoma|9391/3
C1384403|T191|IS|57706008|SNOMEDCT_US|Cellular ependymoma|9391/3
C1384403|T191|OAP|253067007|SNOMEDCT_US|Cellular ependymoma|9391/3
C1384403|T191|OF|253067007|SNOMEDCT_US|Cellular ependymoma|9391/3
C1384403|T191|IS|57706008|SNOMEDCT_US|Clear cell ependymoma|9391/3
C1384403|T191|OF|253068002|SNOMEDCT_US|Clear cell ependymoma|9391/3
C1384403|T191|PT|253068002|SNOMEDCT_US|Clear cell ependymoma|9391/3
C0014474|T191|PT|57706008|SNOMEDCT_US|Ependymoma|9391/3
C0014474|T191|PT|443643007|SNOMEDCT_US|Ependymoma|9391/3
C0014474|T191|SY|57706008|SNOMEDCT_US|Ependymoma, no ICD-O subtype|9391/3
C0014474|T191|SY|57706008|SNOMEDCT_US|Ependymoma, no International Classification of Diseases for Oncology subtype|9391/3
C0014474|T191|IS|57706008|SNOMEDCT_US|Ependymoma, NOS|9391/3
C1370500|T191|IS|397378002|SNOMEDCT_US|Ependymoma, tancytic|9391/3
C1370500|T191|PT|397378002|SNOMEDCT_US|Ependymoma, tanycytic|9391/3
C0014474|T191|OAP|253066003|SNOMEDCT_US|Epithelial ependymoma|9391/3
C0014474|T191|OF|253066003|SNOMEDCT_US|Epithelial ependymoma|9391/3
C0014474|T191|SY|57706008|SNOMEDCT_US|Epithelial ependymoma|9391/3
C4289581|T191|PT|733868000|SNOMEDCT_US|RELA fusion-positive ependymoma|9391/3
C1370500|T191|IS|57706008|SNOMEDCT_US|Tanycytic ependymoma|9391/3
C1370500|T191|SY|397378002|SNOMEDCT_US|Tanycytic ependymoma|9391/3
C0280788|T191|LLT|10002226|MDR|Anaplastic ependymoma|9392/3
C0280788|T191|PT|10014968|MDR|Ependymoma malignant|9392/3
C0280788|T191|LLT|10014968|MDR|Ependymoma malignant|9392/3
C0280788|T191|SY|350016|MEDCIN|CNS neoplasm malignant ependymoma|9392/3
C0280788|T191|PT|350016|MEDCIN|malignant ependymoma|9392/3
C0280788|T191|PEP|D004806|MSH|Anaplastic Ependymoma|9392/3
C0280788|T191|PM|D004806|MSH|Anaplastic Ependymomas|9392/3
C0280788|T191|PM|D004806|MSH|Ependymoma, Anaplastic|9392/3
C0280788|T191|PM|D004806|MSH|Ependymomas, Anaplastic|9392/3
C0280788|T191|PN|NOCODE|MTH|Anaplastic Ependymoma|9392/3
C0280788|T191|SY|C4049|NCI|Anaplastic Ependymal Neoplasm|9392/3
C0280788|T191|SY|C4049|NCI|Anaplastic Ependymal Tumor|9392/3
C0280788|T191|PT|C4049|NCI|Anaplastic Ependymoma|9392/3
C0280788|T191|SY|TCGA|NCI|Anaplastic Ependymoma|9392/3
C0280788|T191|SY|C4049|NCI|Malignant Ependymoma|9392/3
C0280788|T191|SY|C4049|NCI|Undifferentiated Ependymal Neoplasm|9392/3
C0280788|T191|SY|C4049|NCI|Undifferentiated Ependymal Tumor|9392/3
C0280788|T191|SY|C4049|NCI|Undifferentiated Ependymoma|9392/3
C0280788|T191|SY|C4049|NCI|WHO Grade III Ependymal Neoplasm|9392/3
C0280788|T191|SY|C4049|NCI|WHO Grade III Ependymal Tumor|9392/3
C0280788|T191|PT|C4049|NCI_CPTAC|Anaplastic Ependymoma|9392/3
C0280788|T191|PT|BBb8.|RCD|Anaplastic ependymoma|9392/3
C0280788|T191|OAP|134172003|SNOMEDCT_US|Anaplastic ependymoma|9392/3
C0280788|T191|PT|21589007|SNOMEDCT_US|Ependymoma, anaplastic|9392/3
C0334578|T191|PT|MTHU026461|ICPC2ICD10ENG|ependymoma; papillary|9393/3
C0334578|T191|PT|MTHU026462|ICPC2ICD10ENG|ependymoma; papillary, unspecified site|9393/3
C0334578|T191|PT|MTHU057306|ICPC2ICD10ENG|papillary; ependymoma|9393/3
C0334578|T191|PT|MTHU057307|ICPC2ICD10ENG|papillary; ependymoma, unspecified site|9393/3
C0334578|T191|PEP|D004806|MSH|Ependymoma, Papillary|9393/3
C0334578|T191|PM|D004806|MSH|Ependymomas, Papillary|9393/3
C0334578|T191|ET|D004806|MSH|Papillary Ependymoma|9393/3
C0334578|T191|PM|D004806|MSH|Papillary Ependymomas|9393/3
C0334578|T191|PN|NOCODE|MTH|Papillary ependymoma|9393/3
C0334578|T191|PT|C4319|NCI|Papillary Ependymoma|9393/3
C0334578|T191|PT|BBb9.|RCD|Papillary ependymoma|9393/3
C0334578|T191|OAP|112686007|SNOMEDCT_US|Papillary ependymoma|9393/3
C0334578|T191|PT|128839002|SNOMEDCT_US|Papillary ependymoma|9393/3
C0334578|T191|IS|112686007|SNOMEDCT_US|Papillary ependymoma -RETIRED-|9393/3
C0334578|T191|OF|112686007|SNOMEDCT_US|Papillary ependymoma -RETIRED-|9393/3
C0205769|T191|PT|MTHU026458|ICPC2ICD10ENG|ependymoma; myxopapillary|9394/1
C0205769|T191|PT|MTHU026459|ICPC2ICD10ENG|ependymoma; myxopapillary, unspecified site|9394/1
C0205769|T191|PT|MTHU051313|ICPC2ICD10ENG|myxopapillary; ependymoma, unspecified site|9394/1
C0205769|T191|LLT|10014969|MDR|Ependymoma benign|9394/1
C0205769|T191|PT|10014969|MDR|Ependymoma benign|9394/1
C0205769|T191|PEP|D004806|MSH|Ependymoma, Myxopapillary|9394/1
C0205769|T191|PM|D004806|MSH|Ependymomas, Myxopapillary|9394/1
C0205769|T191|PM|D004806|MSH|Myxopapillary Ependymoma|9394/1
C0205769|T191|PM|D004806|MSH|Myxopapillary Ependymomas|9394/1
C0205769|T191|PN|NOCODE|MTH|Myxopapillary ependymoma|9394/1
C0205769|T191|PT|C3697|NCI|Myxopapillary Ependymoma|9394/1
C0205769|T191|SY|TCGA|NCI|Myxopapillary Ependymoma|9394/1
C0205769|T191|PT|C3697|NCI_CDISC|EPENDYMOMA, BENIGN|9394/1
C0205769|T191|PT|BBbA.|RCD|Myxopapillary ependymoma|9394/1
C0205769|T191|PT|1623000|SNOMEDCT_US|Myxopapillary ependymoma|9394/1
C2985219|T191|PT|C92624|NCI|Papillary Tumor of the Pineal Region|9395/3
C2985219|T191|PT|450899004|SNOMEDCT_US|Papillary tumor of the pineal region|9395/3
C2985219|T191|PTGB|450899004|SNOMEDCT_US|Papillary tumour of the pineal region|9395/3
C0004114|T191|ET|0000004651|AOD|astrocytoma|9400/3
C0004114|T191|PT|0000001546|CHV|astrocytoma|9400/3
C0280785|T191|SY|0000057639|CHV|astrocytoma diffuse|9400/3
C0004114|T191|SY|0000001546|CHV|astrocytomas|9400/3
C0004114|T191|SY|0000001546|CHV|astroglioma|9400/3
C0004114|T191|SY|0000001546|CHV|astrogliomas|9400/3
C0280785|T191|PT|0000057639|CHV|diffuse astrocytoma|9400/3
C0004114|T191|PT|U000052|COSTAR|ASTROCYTOMA|9400/3
C0004114|T191|ET|2012-6768|CSP|astrocytic glioma|9400/3
C0004114|T191|PT|2012-6768|CSP|astrocytoma|9400/3
C0004114|T191|ET|2012-6768|CSP|astroglioma|9400/3
C0004114|T191|PT|HP:0009592|HPO|Astrocytoma|9400/3
C0004114|T191|PTN|N74001|ICPC2P|astrocytoma|9400/3
C0004114|T191|PT|N74001|ICPC2P|Astrocytoma|9400/3
C0004114|T191|PT|sh92001188|LCH_NW|Astrocytomas|9400/3
C0004114|T191|PT|10003571|MDR|Astrocytoma|9400/3
C0004114|T191|LLT|10003571|MDR|Astrocytoma|9400/3
C0004114|T191|PM|D001254|MSH|Astrocytic Glioma|9400/3
C0004114|T191|PM|D001254|MSH|Astrocytic Gliomas|9400/3
C0004114|T191|MH|D001254|MSH|Astrocytoma|9400/3
C0280785|T191|PEP|D001254|MSH|Astrocytoma, Grade II|9400/3
C0004114|T191|PM|D001254|MSH|Astrocytomas|9400/3
C0280785|T191|PM|D001254|MSH|Astrocytomas, Grade II|9400/3
C0004114|T191|ET|D001254|MSH|Astroglioma|9400/3
C0004114|T191|PM|D001254|MSH|Astrogliomas|9400/3
C0004114|T191|ET|D001254|MSH|Glioma, Astrocytic|9400/3
C0004114|T191|PM|D001254|MSH|Gliomas, Astrocytic|9400/3
C0280785|T191|PM|D001254|MSH|Grade II Astrocytoma|9400/3
C0280785|T191|PM|D001254|MSH|Grade II Astrocytomas|9400/3
C0004114|T191|PN|NOCODE|MTH|Astrocytoma|9400/3
C0280785|T191|PN|NOCODE|MTH|Diffuse Astrocytoma|9400/3
C0004114|T191|SY|C6958|NCI|Astrocytic Neoplasm|9400/3
C0004114|T191|PT|C6958|NCI|Astrocytic Tumor|9400/3
C0004114|T191|SY|TCGA|NCI|Astrocytoma|9400/3
C0004114|T191|PT|C60781|NCI|Astrocytoma|9400/3
C0004114|T191|SY|C6958|NCI|Astroglioma|9400/3
C0280785|T191|PT|C7173|NCI|Diffuse Astrocytoma|9400/3
C0280785|T191|SY|TCGA|NCI|Diffuse Astrocytoma|9400/3
C0280785|T191|SY|C129277|NCI|Diffuse Astrocytoma, NOS|9400/3
C0280785|T191|PT|C129277|NCI|Diffuse Astrocytoma, Not Otherwise Specified|9400/3
C0280785|T191|SY|C7173|NCI|Grade II Astrocytic Neoplasm|9400/3
C0280785|T191|SY|C7173|NCI|Grade II Astrocytic Tumor|9400/3
C0280785|T191|SY|C7173|NCI|Grade II Astrocytoma|9400/3
C0280785|T191|SY|C7173|NCI|WHO Grade II Astrocytoma|9400/3
C0280785|T191|SY|C7173|NCI_CDISC|Astrocytoma, Diffuse|9400/3
C0280785|T191|PT|C7173|NCI_CDISC|ASTROCYTOMA, DIFFUSE, MALIGNANT|9400/3
C0004114|T191|PT|C60781|NCI_CPTAC|Astrocytoma|9400/3
C0280785|T191|PT|C129277|NCI_CPTAC|Diffuse Astrocytoma, NOS|9400/3
C0280785|T191|PT|10003571|NCI_CTEP-SDC|Low-grade astrocytoma, NOS|9400/3
C0004114|T191|PT|C60781|NCI_CTRP|Astrocytoma|9400/3
C0004114|T191|DN|C60781|NCI_CTRP|Astrocytoma|9400/3
C0004114|T191|PT|CDR0000045602|NCI_NCI-GLOSS|astrocytoma|9400/3
C0004114|T191|PT|C60781|NCI_NICHD|Astrocytoma|9400/3
C0280785|T191|SY|CDR0000041743|PDQ|diffuse astrocytoma|9400/3
C0004114|T191|PT|Xa995|RCD|Astrocytoma|9400/3
C0004114|T191|SY|Xa995|RCDSY|Astrocytoma NOS|9400/3
C0004114|T191|SY|38713004|SNOMEDCT_US|Astrocytic glioma|9400/3
C0004114|T191|OAP|189914005|SNOMEDCT_US|Astrocytoma|9400/3
C0004114|T191|OF|189914005|SNOMEDCT_US|Astrocytoma|9400/3
C0004114|T191|PT|38713004|SNOMEDCT_US|Astrocytoma|9400/3
C0004114|T191|SY|38713004|SNOMEDCT_US|Astrocytoma, no ICD-O subtype|9400/3
C0004114|T191|SY|38713004|SNOMEDCT_US|Astrocytoma, no International Classification of Diseases for Oncology subtype|9400/3
C0004114|T191|IS|38713004|SNOMEDCT_US|Astrocytoma, NOS|9400/3
C0004114|T191|SY|38713004|SNOMEDCT_US|Astroglioma|9400/3
C0280785|T191|PT|397381007|SNOMEDCT_US|Diffuse astrocytoma|9400/3
C0280785|T191|SY|38713004|SNOMEDCT_US|Diffuse astrocytoma|9400/3
C0280785|T191|SY|38713004|SNOMEDCT_US|Diffuse astrocytoma, low grade|9400/3
C4518200|T191|PT|733842007|SNOMEDCT_US|Isocitrate dehydrogenase mutant diffuse astrocytoma|9400/3
C4518199|T191|PT|733841000|SNOMEDCT_US|Isocitrate dehydrogenase wild-type diffuse astrocytoma|9400/3
C0004114|T191|PT|1777|WHO|ASTROCYTOMA|9400/3
C0334579|T191|PT|0000030007|CHV|anaplastic astrocytoma|9401/3
C0334579|T191|SY|0000030007|CHV|anaplastic astrocytomas|9401/3
C0334579|T191|SY|0000030007|CHV|astrocytoma grade iii|9401/3
C0334579|T191|SY|0000030007|CHV|malignant astrocytoma|9401/3
C0334579|T191|ET|2012-6768|CSP|anaplastic astrocytoma|9401/3
C0334579|T191|ET|2012-6410|CSP|anaplastic astrocytoma|9401/3
C0334579|T191|LLT|10002224|MDR|Anaplastic astrocytoma|9401/3
C0334579|T191|PT|10002224|MDR|Anaplastic astrocytoma|9401/3
C0334579|T191|LLT|10060971|MDR|Astrocytoma malignant|9401/3
C0334579|T191|PT|10060971|MDR|Astrocytoma malignant|9401/3
C0334579|T191|LLT|10003572|MDR|Astrocytoma malignant NOS|9401/3
C0334579|T191|PEP|D001254|MSH|Anaplastic Astrocytoma|9401/3
C0334579|T191|PM|D001254|MSH|Anaplastic Astrocytomas|9401/3
C0334579|T191|PM|D001254|MSH|Astrocytoma, Anaplastic|9401/3
C0334579|T191|ET|D001254|MSH|Astrocytoma, Grade III|9401/3
C0334579|T191|PM|D001254|MSH|Astrocytomas, Anaplastic|9401/3
C0334579|T191|PM|D001254|MSH|Astrocytomas, Grade III|9401/3
C0334579|T191|PM|D001254|MSH|Grade III Astrocytoma|9401/3
C0334579|T191|PM|D001254|MSH|Grade III Astrocytomas|9401/3
C0334579|T191|PN|NOCODE|MTH|Anaplastic astrocytoma|9401/3
C0334579|T191|PT|C9477|NCI|Anaplastic Astrocytoma|9401/3
C0334579|T191|SY|TCGA|NCI|Anaplastic Astrocytoma|9401/3
C0334579|T191|SY|C129292|NCI|Anaplastic Astrocytoma, NOS|9401/3
C0334579|T191|PT|C129292|NCI|Anaplastic Astrocytoma, Not Otherwise Specified|9401/3
C0334579|T191|SY|C9477|NCI|Grade III Astrocytic Neoplasm|9401/3
C0334579|T191|SY|C9477|NCI|Grade III Astrocytic Tumor|9401/3
C0334579|T191|SY|C9477|NCI|Grade III Astrocytoma|9401/3
C0334579|T191|SY|C9477|NCI|Malignant Astrocytoma|9401/3
C0334579|T191|PT|C9477|NCI_CPTAC|Anaplastic Astrocytoma|9401/3
C0334579|T191|PT|C129292|NCI_CPTAC|Anaplastic Astrocytoma, NOS|9401/3
C0334579|T191|PT|10002224|NCI_CTEP-SDC|Anaplastic astrocytoma|9401/3
C0334579|T191|PT|10008093|NCI_CTEP-SDC|High-grade astrocytoma, NOS|9401/3
C0334579|T191|PT|BBbC.|RCD|Anaplastic astrocytoma|9401/3
C0334579|T191|SY|BBbC.|RCD|Malignant astrocytoma|9401/3
C0334579|T191|SY|55353007|SNOMEDCT_US|Anaplastic astrocytoma|9401/3
C0334579|T191|PT|55353007|SNOMEDCT_US|Astrocytoma, anaplastic|9401/3
C4518197|T191|PT|733832005|SNOMEDCT_US|Isocitrate dehydrogenase mutant anaplastic astrocytoma|9401/3
C4518198|T191|PT|733840004|SNOMEDCT_US|Isocitrate dehydrogenase wild-type anaplastic astrocytoma|9401/3
C0334579|T191|SY|55353007|SNOMEDCT_US|Malignant astrocytoma|9401/3
C0334580|T191|PEP|D001254|MSH|Astrocytoma, Protoplasmic|9410/3
C0334580|T191|PM|D001254|MSH|Astrocytomas, Protoplasmic|9410/3
C0334580|T191|PM|D001254|MSH|Protoplasmic Astrocytoma|9410/3
C0334580|T191|PM|D001254|MSH|Protoplasmic Astrocytomas|9410/3
C0334580|T191|PN|NOCODE|MTH|Protoplasmic astrocytoma|9410/3
C0334580|T191|PT|C4320|NCI|Protoplasmic Astrocytoma|9410/3
C0334580|T191|PT|BBbD.|RCD|Protoplasmic astrocytoma|9410/3
C0334580|T191|PT|55094006|SNOMEDCT_US|Protoplasmic astrocytoma|9410/3
C0334581|T191|PM|D001254|MSH|Astrocytoma, Gemistocytic|9411/3
C0334581|T191|PM|D001254|MSH|Astrocytomas, Gemistocytic|9411/3
C0334581|T191|PEP|D001254|MSH|Gemistocytic Astrocytoma|9411/3
C0334581|T191|PM|D001254|MSH|Gemistocytic Astrocytomas|9411/3
C0334581|T191|PN|NOCODE|MTH|Gemistocytic astrocytoma|9411/3
C0334581|T191|PT|C4321|NCI|Gemistocytic Astrocytoma|9411/3
C0334581|T191|SY|C4321|NCI|Gemistocytoma|9411/3
C0334581|T191|PT|BBbE.|RCD|Gemistocytic astrocytoma|9411/3
C0334581|T191|PT|73982001|SNOMEDCT_US|Gemistocytic astrocytoma|9411/3
C4518230|T191|PT|733891001|SNOMEDCT_US|Gemistocytic astrocytoma isocitrate dehydrogenase mutation|9411/3
C0334581|T191|SY|73982001|SNOMEDCT_US|Gemistocytoma|9411/3
C0457179|T191|PN|NOCODE|MTH|Desmoplastic infantile astrocytoma|9412/1
C0457179|T191|SY|C9476|NCI|Desmoplastic Astrocytoma of Infancy|9412/1
C0457179|T191|PT|C9476|NCI|Desmoplastic Infantile Astrocytoma|9412/1
C0457179|T191|AB|C9476|NCI|DIA|9412/1
C0457179|T191|PT|C9476|NCI_NICHD|Desmoplastic Infantile Astrocytoma|9412/1
C0457179|T191|PT|128787000|SNOMEDCT_US|Desmoplastic infantile astrocytoma|9412/1
C1266177|T191|MTH_LLT|10072677|MDR|Dysembryoplastic neurepithelial tumor|9413/0
C1266177|T191|MTH_LLT|10072668|MDR|Dysembryoplastic neurepithelial tumor|9413/0
C1266177|T191|LLT|10072668|MDR|Dysembryoplastic neuroepithelial tumor|9413/0
C1266177|T191|LLT|10072677|MDR|Dysembryoplastic neuroepithelial tumour|9413/0
C1266177|T191|PN|NOCODE|MTH|Dysembryoplastic neuroepithelial tumor|9413/0
C1266177|T191|OP|C9505|NCI|DNET|9413/0
C1266177|T191|AB|C9505|NCI|DNT|9413/0
C1266177|T191|SY|C9505|NCI|Dysembryoplastic Neuroepithelial Neoplasm|9413/0
C1266177|T191|PT|C9505|NCI|Dysembryoplastic Neuroepithelial Tumor|9413/0
C1266177|T191|SY|TCGA|NCI|Dysembryoplastic Neuroepithelial Tumor|9413/0
C1266177|T191|PT|87211000119104|SNOMEDCT_US|Dysembryoplastic neuroepithelial tumor|9413/0
C1266177|T191|PT|128788005|SNOMEDCT_US|Dysembryoplastic neuroepithelial tumor|9413/0
C1266177|T191|PTGB|87211000119104|SNOMEDCT_US|Dysembryoplastic neuroepithelial tumour|9413/0
C1266177|T191|PTGB|128788005|SNOMEDCT_US|Dysembryoplastic neuroepithelial tumour|9413/0
C0334582|T191|PT|0000030008|CHV|fibrillary astrocytoma|9420/3
C0334582|T191|PT|MTHU008883|ICPC2ICD10ENG|astrocytoma; fibrillary, unspecified site|9420/3
C0334582|T191|PT|MTHU008882|ICPC2ICD10ENG|astrocytoma; fibrous, unspecified site|9420/3
C0334582|T191|PT|MTHU028125|ICPC2ICD10ENG|fibrillary; astrocytoma, unspecified site|9420/3
C0334582|T191|PT|MTHU028107|ICPC2ICD10ENG|fibrous; astrocytoma, unspecified site|9420/3
C0334582|T191|LLT|10065889|MDR|Fibrillary astrocytoma|9420/3
C0334582|T191|PM|D001254|MSH|Astrocytoma, Fibrillary|9420/3
C0334582|T191|PM|D001254|MSH|Astrocytomas, Fibrillary|9420/3
C0334582|T191|PEP|D001254|MSH|Fibrillary Astrocytoma|9420/3
C0334582|T191|PM|D001254|MSH|Fibrillary Astrocytomas|9420/3
C0334582|T191|PN|NOCODE|MTH|Fibrillary Astrocytoma|9420/3
C0334582|T191|PT|C4322|NCI|Fibrillary Astrocytoma|9420/3
C0334582|T191|PT|10065889|NCI_CTEP-SDC|Fibrillary astrocytoma|9420/3
C0334582|T191|PT|BBbF.|RCD|Fibrillary astrocytoma|9420/3
C0334582|T191|OP|X77pJ|RCD|Fibrous astrocytoma|9420/3
C0334582|T191|PT|71314006|SNOMEDCT_US|Fibrillary astrocytoma|9420/3
C0334582|T191|OAP|253063006|SNOMEDCT_US|Fibrous astrocytoma|9420/3
C0334582|T191|SY|71314006|SNOMEDCT_US|Fibrous astrocytoma|9420/3
C0334583|T191|SY|0000030009|CHV|astrocytoma pilocytic|9421/1
C0334583|T191|PT|0000030009|CHV|pilocytic astrocytoma|9421/1
C0334583|T191|SY|0000030009|CHV|pilocytic astrocytomas|9421/1
C1321865|T191|PT|MTHU008885|ICPC2ICD10ENG|astrocytoma; juvenile, unspecified site|9421/1
C1321865|T191|PT|MTHU040678|ICPC2ICD10ENG|juvenile; astrocytoma, unspecified site|9421/1
C0334583|T191|PM|D001254|MSH|Astrocytoma, Pilocytic|9421/1
C0334583|T191|PM|D001254|MSH|Astrocytomas, Pilocytic|9421/1
C0334583|T191|PEP|D001254|MSH|Pilocytic Astrocytoma|9421/1
C0334583|T191|PM|D001254|MSH|Pilocytic Astrocytomas|9421/1
C1321865|T191|PN|NOCODE|MTH|Juvenile astrocytoma|9421/1
C0334583|T191|PN|NOCODE|MTH|Pilocytic Astrocytoma|9421/1
C1321865|T191|SY|C9022|NCI|Astrocytic Tumors, Childhood|9421/1
C1321865|T191|SY|C9022|NCI|Childhood Astrocytic Neoplasm|9421/1
C1321865|T191|PT|C9022|NCI|Childhood Astrocytic Tumor|9421/1
C1321865|T191|SY|C9022|NCI|Childhood Astrocytic Tumour|9421/1
C0334583|T191|SY|C4047|NCI|Grade I Astrocytic Neoplasm|9421/1
C0334583|T191|SY|C4047|NCI|Grade I Astrocytic Tumor|9421/1
C0334583|T191|SY|C4047|NCI|Grade I Astrocytoma|9421/1
C1321865|T191|SY|C9022|NCI|Pediatric Astrocytic Neoplasm|9421/1
C1321865|T191|SY|C9022|NCI|Pediatric Astrocytic Tumor|9421/1
C0334583|T191|PT|C4047|NCI|Pilocytic Astrocytoma|9421/1
C0334583|T191|SY|TCGA|NCI|Pilocytic Astrocytoma|9421/1
C0334583|T191|PT|90600112|NCI_CTEP-SDC|Pilocytic astrocytoma|9421/1
C1321865|T191|DN|C9022|NCI_CTRP|Astrocytic Tumor|9421/1
C1321865|T191|PT|C9022|NCI_NICHD|Childhood Astrocytic Tumor|9421/1
C1321865|T191|OP|X77pL|RCD|Juvenile astrocytoma|9421/1
C0334583|T191|PT|BBbG.|RCD|Pilocytic astrocytoma|9421/1
C0334583|T191|OP|X77pK|RCD|Piloid astrocytoma|9421/1
C1321865|T191|SY|128854008|SNOMEDCT_US|Juvenile astrocytoma|9421/1
C1321865|T191|IS|67859002|SNOMEDCT_US|Juvenile astrocytoma|9421/1
C1321865|T191|OAP|253065004|SNOMEDCT_US|Juvenile astrocytoma|9421/1
C0334583|T191|PT|763865009|SNOMEDCT_US|Pilocytic astrocytoma|9421/1
C0334583|T191|OAP|67859002|SNOMEDCT_US|Pilocytic astrocytoma|9421/1
C0334583|T191|PT|128854008|SNOMEDCT_US|Pilocytic astrocytoma|9421/1
C0334583|T191|OAP|189915006|SNOMEDCT_US|Pilocytic astrocytoma|9421/1
C0334583|T191|IS|67859002|SNOMEDCT_US|Pilocytic astrocytoma -RETIRED-|9421/1
C0334583|T191|OF|67859002|SNOMEDCT_US|Pilocytic astrocytoma -RETIRED-|9421/1
C0334583|T191|OAP|253064000|SNOMEDCT_US|Piloid astrocytoma|9421/1
C0334583|T191|OF|253064000|SNOMEDCT_US|Piloid astrocytoma|9421/1
C0334583|T191|SY|128854008|SNOMEDCT_US|Piloid astrocytoma|9421/1
C0334583|T191|IS|67859002|SNOMEDCT_US|Piloid astrocytoma|9421/1
C0555199|T191|PT|MTHU060715|ICPC2ICD10ENG|polare; spongioblastoma, unspecified site|9423/3
C0555199|T191|PT|MTHU069101|ICPC2ICD10ENG|spongioblastoma; polare, unspecified site|9423/3
C0555199|T191|PM|D018302|MSH|Polar Spongioblastoma|9423/3
C0555199|T191|PM|D018302|MSH|Polar Spongioblastomas|9423/3
C0555199|T191|PEP|D018302|MSH|Spongioblastoma, Polar|9423/3
C0555199|T191|PM|D018302|MSH|Spongioblastomas, Polar|9423/3
C0555199|T191|PT|C66801|NCI|Polar Spongioblastoma|9423/3
C0555199|T191|OP|C66801|NCI|Polar Spongioblastoma|9423/3
C0555199|T191|OP|Xa997|RCD|Polar spongioblastoma|9423/3
C0334589|T191|OA|BBbP.|RCD|Primitiv polar spongioblastoma|9423/3
C0334589|T191|OP|BBbP.|RCD|Primitive polar spongioblastoma|9423/3
C0555199|T191|OP|BBbJ.|RCD|Spongioblastoma polare|9423/3
C0555199|T191|OAP|134322008|SNOMEDCT_US|Polar spongioblastoma|9423/3
C0555199|T191|OF|134322008|SNOMEDCT_US|Polar spongioblastoma|9423/3
C0555199|T191|PT|12943006|SNOMEDCT_US|Polar spongioblastoma|9423/3
C0334589|T191|OAP|74843007|SNOMEDCT_US|Primitive polar spongioblastoma|9423/3
C0334589|T191|PT|189919000|SNOMEDCT_US|Primitive polar spongioblastoma|9423/3
C0334589|T191|OF|74843007|SNOMEDCT_US|Primitive polar spongioblastoma -RETIRED-|9423/3
C0334589|T191|IS|74843007|SNOMEDCT_US|Primitive polar spongioblastoma -RETIRED-|9423/3
C0555199|T191|SY|12943006|SNOMEDCT_US|Spongioblastoma polare|9423/3
C4283858|T191|PN|NOCODE|MTH|Anaplastic Pleomorphic Xanthoastrocytoma|9424/3
C0334586|T191|PN|NOCODE|MTH|Pleomorphic Xanthoastrocytoma|9424/3
C4283858|T191|PT|C129327|NCI|Anaplastic Pleomorphic Xanthoastrocytoma|9424/3
C4283858|T191|AB|C129327|NCI|APX|9424/3
C0334586|T191|SY|C4323|NCI|Pleomorphic Xantho-Astrocytoma|9424/3
C0334586|T191|SY|TCGA|NCI|Pleomorphic Xanthoastrocytoma|9424/3
C0334586|T191|PT|C4323|NCI|Pleomorphic Xanthoastrocytoma|9424/3
C4283858|T191|SY|C129327|NCI|WHO Grade III Pleomorphic Xanthoastrocytoma|9424/3
C0334586|T191|PT|X77pM|RCD|Pleomorphic xanthoastrocytoma|9424/3
C0334586|T191|AB|X77pM|RCDSY|Pleomorphic xanthoastrocyt|9424/3
C4283858|T191|PT|733848006|SNOMEDCT_US|Anaplastic pleomorphic xanthoastrocytoma|9424/3
C0334586|T191|PT|78838008|SNOMEDCT_US|Pleomorphic xanthoastrocytoma|9424/3
C0334586|T191|OAP|189924002|SNOMEDCT_US|Pleomorphic xanthoastrocytoma|9424/3
C0334586|T191|OF|189924002|SNOMEDCT_US|Pleomorphic xanthoastrocytoma|9424/3
C1519086|T191|PN|NOCODE|MTH|Pilomyxoid astrocytoma|9425/3
C1519086|T191|PT|C40315|NCI|Pilomyxoid Astrocytoma|9425/3
C1519086|T191|IS|388600004|SNOMEDCT_US|Pilomxyoid astrocytoma|9425/3
C1519086|T191|PT|388600004|SNOMEDCT_US|Pilomyxoid astrocytoma|9425/3
C0334587|T191|PT|0000030010|CHV|astroblastoma|9430/3
C0334587|T191|PT|10079366|MDR|Astroblastoma|9430/3
C0334587|T191|LLT|10079366|MDR|Astroblastoma|9430/3
C0334587|T191|PEP|D018302|MSH|Astroblastoma|9430/3
C0334587|T191|PM|D018302|MSH|Astroblastomas|9430/3
C0334587|T191|PN|NOCODE|MTH|Astroblastoma|9430/3
C0334587|T191|PT|C4324|NCI|Astroblastoma|9430/3
C0334587|T191|PT|BBbK.|RCD|Astroblastoma|9430/3
C0334587|T191|PT|48952003|SNOMEDCT_US|Astroblastoma|9430/3
C2363903|T191|LLT|10073129|MDR|Angiocentric glioma|9431/1
C2363903|T191|PT|10073129|MDR|Angiocentric glioma|9431/1
C2363903|T191|MTH_LLT|10068603|MDR|Angiocentric neurepithelial tumor|9431/1
C2363903|T191|MTH_LLT|10068604|MDR|Angiocentric neurepithelial tumor|9431/1
C2363903|T191|LLT|10068603|MDR|Angiocentric neuroepithelial tumor|9431/1
C2363903|T191|LLT|10068604|MDR|Angiocentric neuroepithelial tumour|9431/1
C2363903|T191|PT|C92552|NCI|Angiocentric Glioma|9431/1
C2363903|T191|SY|C92552|NCI|Angiocentric Neuroepithelial Tumor|9431/1
C2363903|T191|SY|C92552|NCI|Monomorphus Angiocentric Glioma|9431/1
C2363903|T191|PT|450900009|SNOMEDCT_US|Angiocentric glioma|9431/1
C2986550|T191|PT|HP:0011754|HPO|Pituicytoma|9432/1
C2986550|T191|PT|C94524|NCI|Pituicytoma|9432/1
C2986550|T191|SY|C94524|NCI|Posterior Pituitary Astrocytoma|9432/1
C2986550|T191|PT|C94524|NCI_CDISC|PITUICYTOMA, BENIGN|9432/1
C2986550|T191|PT|450901008|SNOMEDCT_US|Pituicytoma|9432/1
C2986550|T191|PT|608817003|SNOMEDCT_US|Pituicytoma|9432/1
C0017636|T191|PT|0000005523|CHV|glioblastoma|9440/3
C0017636|T191|SY|0000031708|CHV|glioblastoma|9440/3
C0017636|T191|SY|0000005523|CHV|glioblastomas|9440/3
C0017636|T191|SY|0000031708|CHV|grade iv astrocytoma|9440/3
C0017636|T191|ET|2012-6410|CSP|glioblastoma|9440/3
C0017636|T191|SY|NOCODE|DXP|ASTROCYTOMA, GRADES 3-4|9440/3
C0017636|T191|OP|HP:0100843|HPO|obsolete Glioblastoma|9440/3
C0017636|T191|PT|MTHU032163|ICPC2ICD10ENG|glioblastoma; unspecified site|9440/3
C0017636|T191|PTN|N74012|ICPC2P|glioblastoma|9440/3
C0017636|T191|PT|N74012|ICPC2P|Glioblastoma|9440/3
C0017636|T191|LLT|10018336|MDR|Glioblastoma|9440/3
C0017636|T191|PT|10018336|MDR|Glioblastoma|9440/3
C0017636|T191|ET|D005909|MSH|Astrocytoma, Grade IV|9440/3
C0017636|T191|PM|D005909|MSH|Astrocytomas, Grade IV|9440/3
C0017636|T191|MH|D005909|MSH|Glioblastoma|9440/3
C0017636|T191|PM|D005909|MSH|Glioblastomas|9440/3
C0017636|T191|PM|D005909|MSH|Grade IV Astrocytoma|9440/3
C0017636|T191|PM|D005909|MSH|Grade IV Astrocytomas|9440/3
C0017636|T191|PN|NOCODE|MTH|Glioblastoma|9440/3
C4289580|T191|PT|C129293|NCI|Epithelioid Glioblastoma|9440/3
C0017636|T191|AB|C3058|NCI|GBM|9440/3
C0017636|T191|PT|C3058|NCI|Glioblastoma|9440/3
C0017636|T191|SY|TCGA|NCI|Glioblastoma|9440/3
C0017636|T191|SY|C129295|NCI|Glioblastoma, NOS|9440/3
C0017636|T191|PT|C129295|NCI|Glioblastoma, Not Otherwise Specified|9440/3
C0017636|T191|SY|C3058|NCI|Grade IV Astrocytic Neoplasm|9440/3
C0017636|T191|SY|C3058|NCI|Grade IV Astrocytic Tumor|9440/3
C1272516|T191|PT|C125890|NCI|Small Cell Glioblastoma|9440/3
C0017636|T191|SY|C3058|NCI|WHO Grade IV Glioma|9440/3
C0017636|T191|PT|C3058|NCI_CPTAC|Glioblastoma|9440/3
C0017636|T191|PT|10018337|NCI_CTEP-SDC|Glioblastoma multiforme|9440/3
C0017636|T191|PT|CDR0000539131|NCI_NCI-GLOSS|GBM|9440/3
C0017636|T191|PT|CDR0000045698|NCI_NCI-GLOSS|glioblastoma|9440/3
C0017636|T191|PT|CDR0000044407|NCI_NCI-GLOSS|grade IV astrocytoma|9440/3
C0017636|T191|SY|XM0B6|RCD|Glioblastoma|9440/3
C0017636|T191|OP|XE1wb|RCDSY|Glioblastoma NOS|9440/3
C4289580|T191|PT|733837004|SNOMEDCT_US|Epithelioid glioblastoma|9440/3
C0017636|T191|PT|63634009|SNOMEDCT_US|Glioblastoma|9440/3
C2733135|T191|PT|443811009|SNOMEDCT_US|Glioblastoma - category|9440/3
C4518228|T191|PT|733888001|SNOMEDCT_US|Glioblastoma isocitrate dehydrogenase 1 mutation|9440/3
C4518227|T191|SY|733889009|SNOMEDCT_US|Glioblastoma isocitrate dehydrogenase wild-type|9440/3
C4518227|T191|PT|733889009|SNOMEDCT_US|Glioblastoma isocitrate dehydrogenase wildtype|9440/3
C2733135|T191|SY|443811009|SNOMEDCT_US|Glioblastoma multiforme - category|9440/3
C0017636|T191|SY|63634009|SNOMEDCT_US|Glioblastoma, no ICD-O subtype|9440/3
C0017636|T191|SY|63634009|SNOMEDCT_US|Glioblastoma, no International Classification of Diseases for Oncology subtype|9440/3
C0017636|T191|IS|63634009|SNOMEDCT_US|Glioblastoma, NOS|9440/3
C1272516|T191|PT|384992008|SNOMEDCT_US|Small cell glioblastoma|9440/3
C1272516|T191|SY|384992008|SNOMEDCT_US|Small-cell glioblastoma|9440/3
C0334588|T191|ET|2012-6410|CSP|giant cell glioblastoma|9441/3
C0334588|T191|PT|MTHU064701|ICPC2ICD10ENG|giant cell; glioblastoma, unspecified site|9441/3
C0334588|T191|PT|MTHU032164|ICPC2ICD10ENG|glioblastoma; giant cell, unspecified site|9441/3
C0334588|T191|PEP|D005909|MSH|Giant Cell Glioblastoma|9441/3
C0334588|T191|PM|D005909|MSH|Giant Cell Glioblastomas|9441/3
C0334588|T191|PM|D005909|MSH|Glioblastoma, Giant Cell|9441/3
C0334588|T191|PM|D005909|MSH|Glioblastomas, Giant Cell|9441/3
C0334588|T191|PN|NOCODE|MTH|Giant Cell Glioblastoma|9441/3
C0334588|T191|PT|C4325|NCI|Giant Cell Glioblastoma|9441/3
C0334588|T191|PT|BBbM.|RCD|Giant cell glioblastoma|9441/3
C0334593|T191|PT|BBbX.|RCD|Monstrocellular sarcoma|9441/3
C0334588|T191|PT|44529004|SNOMEDCT_US|Giant cell glioblastoma|9441/3
C0334593|T191|OAP|33556008|SNOMEDCT_US|Monstrocellular sarcoma|9441/3
C0334593|T191|PT|189923008|SNOMEDCT_US|Monstrocellular sarcoma|9441/3
C0334593|T191|IS|33556008|SNOMEDCT_US|Monstrocellular sarcoma -RETIRED-|9441/3
C0334593|T191|OF|33556008|SNOMEDCT_US|Monstrocellular sarcoma -RETIRED-|9441/3
C1266178|T191|PT|C5419|NCI|Gliofibroma|9442/1
C1266178|T191|PT|128909006|SNOMEDCT_US|Gliofibroma|9442/1
C0206726|T191|PT|0000021050|CHV|gliosarcoma|9442/3
C0206726|T191|ET|2012-6589|CSP|gliosarcoma|9442/3
C0206726|T191|PT|MTHU032171|ICPC2ICD10ENG|gliosarcoma; unspecified site|9442/3
C0206726|T191|PT|10018340|MDR|Gliosarcoma|9442/3
C0206726|T191|LLT|10018340|MDR|Gliosarcoma|9442/3
C0206726|T191|ET|D018316|MSH|Glioblastoma with Sarcomatous Component|9442/3
C0206726|T191|PM|D018316|MSH|Glioma, Sarcomatous|9442/3
C0206726|T191|PM|D018316|MSH|Gliomas, Sarcomatous|9442/3
C0206726|T191|MH|D018316|MSH|Gliosarcoma|9442/3
C0206726|T191|PM|D018316|MSH|Gliosarcomas|9442/3
C0206726|T191|ET|D018316|MSH|Sarcomatous Glioma|9442/3
C0206726|T191|PM|D018316|MSH|Sarcomatous Gliomas|9442/3
C0206726|T191|PN|NOCODE|MTH|gliosarcoma|9442/3
C0206726|T191|SY|C3796|NCI|Glioblastoma with a Sarcomatous Component|9442/3
C0206726|T191|PT|C3796|NCI|Gliosarcoma|9442/3
C0206726|T191|SY|TCGA|NCI|Gliosarcoma|9442/3
C0206726|T191|PT|CDR0000045701|NCI_NCI-GLOSS|gliosarcoma|9442/3
C0206726|T191|OA|BBbN.|RCD|Glioblastoma sarcoma component|9442/3
C0206726|T191|OP|BBbN.|RCD|Glioblastoma with sarcomatous component|9442/3
C0206726|T191|PT|X77pN|RCD|Gliosarcoma|9442/3
C0206726|T191|SY|35262004|SNOMEDCT_US|Glioblastoma with sarcomatous component|9442/3
C0206726|T191|OAP|189918008|SNOMEDCT_US|Glioblastoma with sarcomatous component|9442/3
C0206726|T191|OF|189918008|SNOMEDCT_US|Glioblastoma with sarcomatous component|9442/3
C0206726|T191|PT|35262004|SNOMEDCT_US|Gliosarcoma|9442/3
C1322252|T191|PN|NOCODE|MTH|Chordoid Glioma of the Third Ventricle|9444/1
C1322252|T191|SY|C5592|NCI|Chordoid Glioma|9444/1
C1322252|T191|SY|C5592|NCI|Chordoid Glioma of 3rd Ventricle|9444/1
C1322252|T191|SY|C5592|NCI|Chordoid Glioma of the 3rd Ventricle|9444/1
C1322252|T191|PT|C5592|NCI|Chordoid Glioma of the Third Ventricle|9444/1
C1322252|T191|SY|C5592|NCI|Chordoid Glioma of Third Ventricle|9444/1
C1322252|T191|SY|C5592|NCI|Third Ventricle Chordoid Glioma|9444/1
C1322252|T191|PT|715900001|SNOMEDCT_US|Chordoid glioma|9444/1
C1322252|T191|PT|128789002|SNOMEDCT_US|Chordoid glioma|9444/1
C1322252|T191|SY|128789002|SNOMEDCT_US|Chordoid glioma of third ventricle|9444/1
C0751396|T191|PT|0000008930|CHV|oligodendroglioma|9450/3
C0751396|T191|SY|0000008930|CHV|oligodendrogliomas|9450/3
C0751396|T191|ET|2012-6589|CSP|oligodendroglioma|9450/3
C0751396|T191|LLT|10030286|MDR|Oligodendroglioma|9450/3
C0751396|T191|PT|10030286|MDR|Oligodendroglioma|9450/3
C0028945|T191|MH|D009837|MSH|Oligodendroglioma|9450/3
C0751396|T191|DEV|D009837|MSH|OLIGODENDROGLIOMA WELL DIFFER|9450/3
C0751396|T191|PM|D009837|MSH|Oligodendroglioma, Well Differentiated|9450/3
C0751396|T191|PEP|D009837|MSH|Oligodendroglioma, Well-Differentiated|9450/3
C0028945|T191|PM|D009837|MSH|Oligodendrogliomas|9450/3
C0751396|T191|PM|D009837|MSH|Oligodendrogliomas, Well-Differentiated|9450/3
C0751396|T191|DEV|D009837|MSH|WELL DIFFER OLIGODENDROGLIOMA|9450/3
C0751396|T191|PM|D009837|MSH|Well Differentiated Oligodendroglioma|9450/3
C0751396|T191|ET|D009837|MSH|Well-Differentiated Oligodendroglioma|9450/3
C0751396|T191|PM|D009837|MSH|Well-Differentiated Oligodendrogliomas|9450/3
C0028945|T191|PN|NOCODE|MTH|oligodendroglioma|9450/3
C0751396|T191|PN|NOCODE|MTH|Well Differentiated Oligodendroglioma|9450/3
C0751396|T191|SY|TCGA|NCI|Oligodendroglioma|9450/3
C0751396|T191|PT|C3288|NCI|Oligodendroglioma|9450/3
C0028945|T191|SY|C129319|NCI|Oligodendroglioma, NOS|9450/3
C0028945|T191|PT|C129319|NCI|Oligodendroglioma, Not Otherwise Specified|9450/3
C0751396|T191|SY|C3288|NCI|Well Differentiated Oligodendroglial Tumor|9450/3
C0751396|T191|SY|C3288|NCI|Well Differentiated Oligodendroglioma|9450/3
C0751396|T191|SY|C3288|NCI|WHO Grade II Oligodendroglial Neoplasm|9450/3
C0751396|T191|SY|C3288|NCI|WHO Grade II Oligodendroglial Tumor|9450/3
C0028945|T191|PT|C129319|NCI_CPTAC|Oligodendroglioma, NOS|9450/3
C0751396|T191|PT|10030286|NCI_CTEP-SDC|Oligodendroglioma, NOS|9450/3
C0751396|T191|PT|CDR0000046257|NCI_NCI-GLOSS|oligodendroglioma|9450/3
C0751396|T191|PT|Xa998|RCD|Oligodendroglioma|9450/3
C0751396|T191|OP|BBbQ.|RCDSY|Oligodendroglioma NOS|9450/3
C0028945|T191|SY|73348003|SNOMEDCT_US|Oligodendroglioma|9450/3
C0751396|T191|PT|443936004|SNOMEDCT_US|Oligodendroglioma|9450/3
C2732301|T191|PT|443565000|SNOMEDCT_US|Oligodendroglioma - category|9450/3
C4518383|T191|PT|734086009|SNOMEDCT_US|Oligodendroglioma with isocitrate dehydrogenase mutant and 1p/19q-codeleted|9450/3
C0028945|T191|PT|73348003|SNOMEDCT_US|Oligodendroglioma, no ICD-O subtype|9450/3
C0028945|T191|SY|73348003|SNOMEDCT_US|Oligodendroglioma, no International Classification of Diseases for Oncology subtype|9450/3
C0028945|T191|IS|73348003|SNOMEDCT_US|Oligodendroglioma, NOS|9450/3
C0334590|T191|PT|0000030011|CHV|anaplastic oligodendroglioma|9451/3
C0334590|T191|SY|0000030011|CHV|anaplastic oligodendrogliomas|9451/3
C0334590|T191|PT|10073128|MDR|Anaplastic oligodendroglioma|9451/3
C0334590|T191|LLT|10073128|MDR|Anaplastic oligodendroglioma|9451/3
C0334590|T191|LLT|10026659|MDR|Malignant oligodendroglioma|9451/3
C0334590|T191|PT|10026659|MDR|Malignant oligodendroglioma|9451/3
C0334590|T191|LLT|10030288|MDR|Oligodendroglioma malignant|9451/3
C0334590|T191|SY|350017|MEDCIN|CNS neoplasm malignant oligodendroglioma|9451/3
C0334590|T191|PT|350017|MEDCIN|malignant oligodendroglioma|9451/3
C0334590|T191|PEP|D009837|MSH|Anaplastic Oligodendroglioma|9451/3
C0334590|T191|PM|D009837|MSH|Anaplastic Oligodendrogliomas|9451/3
C0334590|T191|PM|D009837|MSH|Oligodendroglioma, Anaplastic|9451/3
C0334590|T191|PM|D009837|MSH|Oligodendrogliomas, Anaplastic|9451/3
C0334590|T191|PN|NOCODE|MTH|Anaplastic Oligodendroglioma|9451/3
C0334590|T191|SY|TCGA|NCI|Anaplastic Oligodendroglioma|9451/3
C0334590|T191|PT|C4326|NCI|Anaplastic Oligodendroglioma|9451/3
C0334590|T191|SY|C129322|NCI|Anaplastic Oligodendroglioma, NOS|9451/3
C0334590|T191|PT|C129322|NCI|Anaplastic Oligodendroglioma, Not Otherwise Specified|9451/3
C0334590|T191|SY|C4326|NCI|Malignant Oligodendroglioma|9451/3
C0334590|T191|SY|C4326|NCI|Oligodendroglioma, Malignant|9451/3
C0334590|T191|SY|C4326|NCI|Undifferentiated Oligodendroglioma|9451/3
C0334590|T191|SY|C4326|NCI|WHO Grade III Oligodendroglial Neoplasm|9451/3
C0334590|T191|SY|C4326|NCI|WHO Grade III Oligodendroglial Tumor|9451/3
C0334590|T191|PT|C129322|NCI_CPTAC|Anaplastic Oligodendroglioma, NOS|9451/3
C0334590|T191|PT|10026659|NCI_CTEP-SDC|Anaplastic oligodendroglioma|9451/3
C0334590|T191|PT|BBbR.|RCD|Anaplastic oligodendroglioma|9451/3
C0334590|T191|SY|3102004|SNOMEDCT_US|Anaplastic oligodendroglioma|9451/3
C4518384|T191|PT|733843002|SNOMEDCT_US|Anaplastic oligodendroglioma with isocitrate dehydrogenase mutant and 1p/19q-codeleted|9451/3
C0334590|T191|PT|3102004|SNOMEDCT_US|Oligodendroglioma, anaplastic|9451/3
C0344461|T191|PEP|D009837|MSH|Oligodendroblastoma|9460/3
C0344461|T191|PM|D009837|MSH|Oligodendroblastomas|9460/3
C0344461|T191|PT|C66802|NCI|Oligodendroblastoma|9460/3
C0344461|T191|OP|C66802|NCI|Oligodendroblastoma|9460/3
C0344461|T191|OP|BBbS.|RCD|Oligodendroblastoma|9460/3
C0344461|T191|PT|80061003|SNOMEDCT_US|Oligodendroblastoma|9460/3
C0025149|T191|ET|0000004649|AOD|medulloblastoma|9470/3
C0025149|T191|SY|0000007877|CHV|brain medulloblastoma tumors|9470/3
C0025149|T191|PT|0000007877|CHV|medulloblastoma|9470/3
C0025149|T191|SY|0000007877|CHV|medulloblastoma brain tumor|9470/3
C0025149|T191|SY|0000007877|CHV|medulloblastomas|9470/3
C0025149|T191|PT|2006-5547|CSP|medulloblastoma|9470/3
C0025149|T191|SY|NOCODE|DXP|BRAIN TUMOR, MEDULLOBLASTOMA|9470/3
C0025149|T191|DI|U000241|DXP|BRAIN, MEDULLOBLASTOMA|9470/3
C0025149|T191|SY|NOCODE|DXP|INTRACRANIAL NEOPLASM, MEDULLOBLASTOMA|9470/3
C0025149|T191|PT|HP:0002885|HPO|Medulloblastoma|9470/3
C0025149|T191|PT|U002880|LCH|Medulloblastoma|9470/3
C0025149|T191|PT|sh85083247|LCH_NW|Medulloblastoma|9470/3
C0025149|T191|LLT|10027107|MDR|Medulloblastoma|9470/3
C0025149|T191|PT|10027107|MDR|Medulloblastoma|9470/3
C0025149|T191|SY|31905|MEDCIN|central nervous system mass lesions cerebellum medulloblastoma|9470/3
C0025149|T191|PT|358400|MEDCIN|medulloblastoma|9470/3
C0025149|T191|PT|31905|MEDCIN|medulloblastoma of cerebellum|9470/3
C0025149|T191|SY|358400|MEDCIN|neuroendocrine tumor medulloblastoma|9470/3
C0025149|T191|MH|D008527|MSH|Medulloblastoma|9470/3
C1275668|T191|PM|D008527|MSH|Medulloblastoma, Melanocytic|9470/3
C0025149|T191|PM|D008527|MSH|Medulloblastomas|9470/3
C1275668|T191|PM|D008527|MSH|Medulloblastomas, Melanocytic|9470/3
C1275668|T191|PEP|D008527|MSH|Melanocytic Medulloblastoma|9470/3
C1275668|T191|PM|D008527|MSH|Melanocytic Medulloblastomas|9470/3
C0025149|T191|PN|NOCODE|MTH|Medulloblastoma|9470/3
C1275668|T191|PN|NOCODE|MTH|Melanotic medulloblastoma|9470/3
C1707400|T191|PT|C54039|NCI|Classic Medulloblastoma|9470/3
C0025149|T191|SY|TCGA|NCI|Medulloblastoma|9470/3
C0025149|T191|PT|C3222|NCI|Medulloblastoma|9470/3
C1275668|T191|PT|C9497|NCI|Medulloblastoma with Melanotic Differentiation|9470/3
C1275668|T191|SY|TCGA|NCI|Medulloblastoma with Melanotic Differentiation|9470/3
C1275668|T191|SY|C9497|NCI|Melanocytic Medulloblastoma|9470/3
C1275668|T191|SY|C9497|NCI|Melanotic Medulloblastoma|9470/3
C0025149|T191|PT|C3222|NCI_CDISC|MEDULLOBLASTOMA, MALIGNANT|9470/3
C0025149|T191|SY|C3222|NCI_CDISC|Medulloblastomas|9470/3
C0025149|T191|PT|10027107|NCI_CTEP-SDC|Medulloblastoma|9470/3
C0025149|T191|PT|CDR0000045780|NCI_NCI-GLOSS|medulloblastoma|9470/3
C0025149|T191|PT|C3222|NCI_NICHD|Medulloblastoma|9470/3
C0025149|T191|SY|Xa999|RCD|MDB - Medulloblastoma|9470/3
C0025149|T191|PT|Xa999|RCD|Medulloblastoma|9470/3
C0025149|T191|OP|BBbT.|RCDSY|Medulloblastoma NOS|9470/3
C1707400|T191|PT|699703008|SNOMEDCT_US|Classic medulloblastoma|9470/3
C1707400|T191|PT|699704002|SNOMEDCT_US|Classic medulloblastoma|9470/3
C0025149|T191|SY|83217000|SNOMEDCT_US|MDB - Medulloblastoma|9470/3
C0025149|T191|PT|443333004|SNOMEDCT_US|Medulloblastoma|9470/3
C0025149|T191|PT|83217000|SNOMEDCT_US|Medulloblastoma|9470/3
C2732566|T191|PT|443334005|SNOMEDCT_US|Medulloblastoma - category|9470/3
C1275668|T191|PT|397380008|SNOMEDCT_US|Medulloblastoma, melanotic|9470/3
C0025149|T191|SY|83217000|SNOMEDCT_US|Medulloblastoma, no ICD-O subtype|9470/3
C0025149|T191|SY|83217000|SNOMEDCT_US|Medulloblastoma, no International Classification of Diseases for Oncology subtype|9470/3
C0025149|T191|IS|83217000|SNOMEDCT_US|Medulloblastoma, NOS|9470/3
C1275668|T191|SY|83217000|SNOMEDCT_US|Melanotic medulloblastoma|9470/3
C1275668|T191|SY|397380008|SNOMEDCT_US|Melanotic medulloblastoma|9470/3
C4518406|T191|PT|734073000|SNOMEDCT_US|Non-wingless and non-sonic hedgehog medulloblastoma|9470/3
C4518214|T191|PT|733872001|SNOMEDCT_US|Sonic hedgehog pathway activated and tumor protein p53 mutant medulloblastoma|9470/3
C4518214|T191|PTGB|733872001|SNOMEDCT_US|Sonic hedgehog pathway activated and tumour protein p53 mutant medulloblastoma|9470/3
C4518357|T191|PT|733909005|SNOMEDCT_US|Wingless-activated medulloblastoma|9470/3
C0751291|T191|PT|MTHU022673|ICPC2ICD10ENG|desmoplastic; medulloblastoma|9471/3
C0751291|T191|PT|MTHU048017|ICPC2ICD10ENG|medulloblastoma; desmoplastic|9471/3
C0751291|T191|PEP|D008527|MSH|Arachnoidal Cerebellar Sarcoma, Circumscribed|9471/3
C0751291|T191|PM|D008527|MSH|Desmoplastic Medulloblastoma|9471/3
C0751291|T191|PM|D008527|MSH|Desmoplastic Medulloblastomas|9471/3
C0751291|T191|ET|D008527|MSH|Medulloblastoma, Desmoplastic|9471/3
C0751291|T191|PM|D008527|MSH|Medulloblastomas, Desmoplastic|9471/3
C0751291|T191|ET|D008527|MSH|Sarcoma, Cerebellar, Circumscribed Arachnoidal|9471/3
C0751291|T191|PN|NOCODE|MTH|Desmoplastic Medulloblastoma|9471/3
C1334970|T191|SY|C5407|NCI|Cerebellar Neuroblastoma|9471/3
C0751291|T191|SY|C4956|NCI|Desmoplastic Medulloblastoma|9471/3
C0751291|T191|SY|C4956|NCI|Desmoplastic Nodular Medulloblastoma|9471/3
C0751291|T191|PT|C4956|NCI|Desmoplastic/Nodular Medulloblastoma|9471/3
C0751291|T191|SY|TCGA|NCI|Desmoplastic/Nodular Medulloblastoma|9471/3
C1334970|T191|PT|C5407|NCI|Medulloblastoma with Extensive Nodularity|9471/3
C1334970|T191|SY|C5407|NCI|Medulloblastoma with Extensive Nodularity and Advanced Neuronal Differentiation|9471/3
C1334970|T191|SY|C5407|NCI|Nodular Medulloblastoma|9471/3
C0751291|T191|PT|BBbU.|RCD|Desmoplastic medulloblastoma|9471/3
C0751291|T191|SY|32456001|SNOMEDCT_US|Circumscribed arachnoidal cerebellar sarcoma|9471/3
C0751291|T191|PT|32456001|SNOMEDCT_US|Desmoplastic medulloblastoma|9471/3
C0751291|T191|SY|32456001|SNOMEDCT_US|Desmoplastic nodular medulloblastoma|9471/3
C1334970|T191|PT|733902001|SNOMEDCT_US|Medulloblastoma with extensive nodularity|9471/3
C0751291|T191|IS|32456001|SNOMEDCT_US|Medulloblastoma with extensive nodularity and advanced neuronal differentiation.|9471/3
C4518213|T191|PT|733874000|SNOMEDCT_US|Sonic hedgehog pathway activated and tumor protein p53 wild-type medulloblastoma|9471/3
C4518213|T191|PTGB|733874000|SNOMEDCT_US|Sonic hedgehog pathway activated and tumour protein p53 wild-type medulloblastoma|9471/3
C0205833|T191|PEP|D008527|MSH|Medullomyoblastoma|9472/3
C0205833|T191|PM|D008527|MSH|Medullomyoblastomas|9472/3
C0205833|T191|PN|NOCODE|MTH|Medullomyoblastoma|9472/3
C0205833|T191|SY|C3706|NCI|Medullomyoblastoma|9472/3
C0205833|T191|PT|C3706|NCI|Medullomyoblastoma with Myogenic Differentiation|9472/3
C0205833|T191|PT|BBbV.|RCD|Medullomyoblastoma|9472/3
C0431114|T191|PT|X77pc|RCD|Melanocytic medullomyoblastoma|9472/3
C0205833|T191|PT|24604009|SNOMEDCT_US|Medullomyoblastoma|9472/3
C0431114|T191|PT|253077009|SNOMEDCT_US|Melanocytic medullomyoblastoma|9472/3
C0206663|T191|SY|0000042698|CHV|neuroectodermal primitive tumors|9473/3
C0206663|T191|SY|0000021005|CHV|pnet|9473/3
C0206663|T191|SY|0000021005|CHV|primitive neuroectodermal tumor|9473/3
C0206663|T191|PT|0000042698|CHV|primitive neuroectodermal tumors|9473/3
C0206663|T191|SY|0000021005|CHV|primitive neuroectodermal tumors|9473/3
C0206663|T191|SY|0000021005|CHV|primitive neuroectodermal tumour|9473/3
C0206663|T191|PT|HP:0030065|HPO|Primitive neuroectodermal tumor|9473/3
C0206663|T191|PT|MTHU052504|ICPC2ICD10ENG|neuroectodermal; tumor, primitive, unspecified site|9473/3
C0206663|T191|PT|MTHU061687|ICPC2ICD10ENG|primitive; neuroectodermal tumor, unspecified site|9473/3
C0206663|T191|PT|MTHU077105|ICPC2ICD10ENG|tumor; neuroectodermal, primitive, unspecified site|9473/3
C0206663|T191|LLT|10057849|MDR|Primitive neuroectodermal tumor|9473/3
C0206663|T191|MTH_PT|10057846|MDR|Primitive neuroectodermal tumor|9473/3
C0206663|T191|LLT|10057846|MDR|Primitive neuroectodermal tumour|9473/3
C0206663|T191|PT|10057846|MDR|Primitive neuroectodermal tumour|9473/3
C0206663|T191|PT|271567|MEDCIN|neuroepithelioma|9473/3
C0206663|T191|DEV|D018242|MSH|NEOPL PRIMITIVE NEUROEPITHELIAL|9473/3
C0206663|T191|PM|D018242|MSH|Neoplasm, Primitive Neuroepithelial|9473/3
C0206663|T191|ET|D018242|MSH|Neoplasms, Primitive Neuroepithelial|9473/3
C0206663|T191|ET|D018242|MSH|Neuroectodermal Tumor, Primitive|9473/3
C0206663|T191|MH|D018242|MSH|Neuroectodermal Tumors, Primitive|9473/3
C0206663|T191|DEV|D018242|MSH|NEUROEPITHELIAL NEOPL PRIMITIVE|9473/3
C0206663|T191|PM|D018242|MSH|Neuroepithelial Neoplasm, Primitive|9473/3
C0206663|T191|ET|D018242|MSH|Neuroepithelial Neoplasms, Primitive|9473/3
C0206663|T191|PM|D018242|MSH|Neuroepithelial Tumor, Primitive|9473/3
C0206663|T191|ET|D018242|MSH|Neuroepithelial Tumors, Primitive|9473/3
C0206663|T191|ET|D018242|MSH|PNET|9473/3
C0206663|T191|PM|D018242|MSH|PNETs|9473/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroectodermal Tumor|9473/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroectodermal Tumors|9473/3
C0206663|T191|DEV|D018242|MSH|PRIMITIVE NEUROEPITHELIAL NEOPL|9473/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroepithelial Neoplasm|9473/3
C0206663|T191|ET|D018242|MSH|Primitive Neuroepithelial Neoplasms|9473/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroepithelial Tumor|9473/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroepithelial Tumors|9473/3
C0206663|T191|PM|D018242|MSH|Tumor, Primitive Neuroectodermal|9473/3
C0206663|T191|PM|D018242|MSH|Tumor, Primitive Neuroepithelial|9473/3
C0206663|T191|PM|D018242|MSH|Tumors, Primitive Neuroectodermal|9473/3
C0206663|T191|PM|D018242|MSH|Tumors, Primitive Neuroepithelial|9473/3
C0206663|T191|PN|NOCODE|MTH|Neuroectodermal Tumor, Primitive|9473/3
C0206663|T191|SY|C3716|NCI|Neuroectodermal Neoplasm|9473/3
C0206663|T191|SY|C3716|NCI|Neuroectodermal Tumor|9473/3
C0206663|T191|SY|C3716|NCI|Neuroepithelioma|9473/3
C0206663|T191|AB|C3716|NCI|PNET|9473/3
C0206663|T191|SY|C3716|NCI|Primitive Neuroectodermal Neoplasm|9473/3
C0206663|T191|SY|TCGA|NCI|Primitive Neuroectodermal Tumor|9473/3
C0206663|T191|PT|C3716|NCI|Primitive Neuroectodermal Tumor|9473/3
C0206663|T191|PT|C3716|NCI_CPTAC|Primitive Neuroectodermal Tumor|9473/3
C0206663|T191|PT|C3716|NCI_CTRP|Primitive Neuroectodermal Tumor|9473/3
C0206663|T191|PT|CDR0000045952|NCI_NCI-GLOSS|neuroectodermal tumor|9473/3
C0206663|T191|PT|CDR0000383924|NCI_NCI-GLOSS|PNET|9473/3
C0206663|T191|PT|CDR0000383920|NCI_NCI-GLOSS|primitive neuroectodermal tumor|9473/3
C0206663|T191|SY|CDR0000039466|PDQ|PNET|9473/3
C0206663|T191|PT|Xa99H|RCD|Neuroepithelioma|9473/3
C0206663|T191|AB|X77pa|RCD|PNET - Primit neuroect tumour|9473/3
C0206663|T191|SY|X77pa|RCD|PNET - Primitive neuroectodermal tumour|9473/3
C0206663|T191|AB|X77pa|RCD|Primitive neuroectodermal tum|9473/3
C0206663|T191|PT|X77pa|RCD|Primitive neuroectodermal tumour|9473/3
C0206663|T191|AB|X77pa|RCDAE|PNET - Primit neuroect tumor|9473/3
C0206663|T191|SY|X77pa|RCDAE|PNET - Primitive neuroectodermal tumor|9473/3
C0206663|T191|PT|X77pa|RCDAE|Primitive neuroectodermal tumor|9473/3
C0206663|T191|OP|BBc4.|RCDSY|Neuroepithelioma NOS|9473/3
C0206663|T191|AB|X77pa|RCDSY|Primit neuroectodermal tumr|9473/3
C0206663|T191|PT|55045006|SNOMEDCT_US|Neuroepithelioma|9473/3
C0206663|T191|IS|55045006|SNOMEDCT_US|Neuroepithelioma, NOS|9473/3
C0206663|T191|SY|39781001|SNOMEDCT_US|PNET|9473/3
C0206663|T191|SY|39781001|SNOMEDCT_US|PNET - Primitive neuroectodermal tumor|9473/3
C0206663|T191|SYGB|39781001|SNOMEDCT_US|PNET - Primitive neuroectodermal tumour|9473/3
C0206663|T191|PT|699028006|SNOMEDCT_US|Primitive neuroectodermal tumor|9473/3
C0206663|T191|PT|39781001|SNOMEDCT_US|Primitive neuroectodermal tumor|9473/3
C0206663|T191|OAP|189925001|SNOMEDCT_US|Primitive neuroectodermal tumor|9473/3
C0206663|T191|OAP|189925001|SNOMEDCT_US|Primitive neuroectodermal tumour|9473/3
C0206663|T191|OF|189925001|SNOMEDCT_US|Primitive neuroectodermal tumour|9473/3
C0206663|T191|PTGB|699028006|SNOMEDCT_US|Primitive neuroectodermal tumour|9473/3
C0206663|T191|PTGB|39781001|SNOMEDCT_US|Primitive neuroectodermal tumour|9473/3
C1266180|T191|PN|NOCODE|MTH|Large cell medulloblastoma|9474/3
C2985220|T191|PT|C92625|NCI|Anaplastic Medulloblastoma|9474/3
C1266180|T191|PT|C6904|NCI|Large Cell Medulloblastoma|9474/3
C1266180|T191|SY|TCGA|NCI|Large Cell Medulloblastoma|9474/3
C1266180|T191|PT|128790006|SNOMEDCT_US|Large cell medulloblastoma|9474/3
C0334592|T191|PT|MTHU015510|ICPC2ICD10ENG|cerebellar; sarcoma|9480/3
C0334592|T191|PT|MTHU065890|ICPC2ICD10ENG|sarcoma; cerebellar|9480/3
C0334592|T191|PT|213034|MEDCIN|cerebellar sarcoma|9480/3
C0334592|T191|PT|236019|MEDCIN|sarcoma of cerebellum|9480/3
C0334592|T191|OP|C66803|NCI|Cerebellar Sarcoma|9480/3
C0334592|T191|PT|C66803|NCI|Cerebellar Sarcoma|9480/3
C0334592|T191|PT|Xa99A|RCD|Cerebellar sarcoma|9480/3
C0334592|T191|OP|BBbW.|RCDSY|Cerebellar sarcoma NOS|9480/3
C0334592|T191|PT|17302008|SNOMEDCT_US|Cerebellar sarcoma|9480/3
C0334592|T191|IS|17302008|SNOMEDCT_US|Cerebellar sarcoma, NOS|9480/3
C0017075|T191|ET|0000004647|AOD|ganglioneuroma|9490/0
C0017075|T191|SY|0000005343|CHV|gangliocytoma|9490/0
C0017075|T191|SY|0000005343|CHV|gangliocytomas|9490/0
C0017075|T191|PT|0000005343|CHV|ganglioneuroma|9490/0
C0017075|T191|SY|0000005343|CHV|ganglioneuromas|9490/0
C0017075|T191|SY|NOCODE|DXP|GANGLIONEUROFIBROMA|9490/0
C0017075|T191|DI|U000693|DXP|GANGLIONEUROMA|9490/0
C0017075|T191|PT|HP:0003005|HPO|Ganglioneuroma|9490/0
C0017075|T191|PT|MTHU030261|ICPC2ICD10ENG|gangliocytoma|9490/0
C0017075|T191|PT|MTHU030278|ICPC2ICD10ENG|ganglioneuroma|9490/0
C0017075|T191|LA|LA26521-7|LNC|Ganglioneuroma|9490/0
C0017075|T191|LLT|10017700|MDR|Gangliocytoma|9490/0
C0017075|T191|PT|10017709|MDR|Ganglioneuroma|9490/0
C0017075|T191|LLT|10017709|MDR|Ganglioneuroma|9490/0
C0017075|T191|ET|D005729|MSH|Gangliocytoma|9490/0
C0017075|T191|PM|D005729|MSH|Gangliocytomas|9490/0
C0017075|T191|MH|D005729|MSH|Ganglioneuroma|9490/0
C0017075|T191|PM|D005729|MSH|Ganglioneuromas|9490/0
C0017075|T191|PN|NOCODE|MTH|Ganglioneuroma|9490/0
C0017075|T191|PT|C6934|NCI|Gangliocytoma|9490/0
C0017075|T191|SY|TCGA|NCI|Gangliocytoma|9490/0
C0017075|T191|PT|C3049|NCI|Ganglioneuroma|9490/0
C0017075|T191|PT|C3049|NCI_CDISC|GANGLIONEUROMA, BENIGN|9490/0
C0017075|T191|SY|C3049|NCI_CDISC|Neural Crest Tumor, Benign|9490/0
C0017075|T191|DN|C3049|NCI_CTRP|Ganglioneuroma|9490/0
C0017075|T191|PT|X77pU|RCD|Gangliocytoma|9490/0
C0017075|T191|PT|BBc00|RCD|Ganglioneuroma|9490/0
C0017075|T191|PT|128919000|SNOMEDCT_US|Gangliocytoma|9490/0
C0017075|T191|IS|53801007|SNOMEDCT_US|Gangliocytoma|9490/0
C0017075|T191|PT|116371000119107|SNOMEDCT_US|Ganglioneuroma|9490/0
C0017075|T191|OAP|189929007|SNOMEDCT_US|Ganglioneuroma|9490/0
C0017075|T191|PT|53801007|SNOMEDCT_US|Ganglioneuroma|9490/0
C0206718|T191|PT|0000021044|CHV|ganglioneuroblastoma|9490/3
C0206718|T191|SY|0000021044|CHV|ganglioneuroblastomas|9490/3
C0206718|T191|PT|HP:0006747|HPO|Ganglioneuroblastoma|9490/3
C0206718|T191|PT|10017708|MDR|Ganglioneuroblastoma|9490/3
C0206718|T191|LLT|10017708|MDR|Ganglioneuroblastoma|9490/3
C0206718|T191|PT|271564|MEDCIN|ganglioneuroblastoma|9490/3
C0206718|T191|MH|D018305|MSH|Ganglioneuroblastoma|9490/3
C0206718|T191|PM|D018305|MSH|Ganglioneuroblastomas|9490/3
C0206718|T191|PN|NOCODE|MTH|Ganglioneuroblastoma|9490/3
C0206718|T191|PT|C3790|NCI|Ganglioneuroblastoma|9490/3
C1517444|T191|PT|C42057|NCI|Ganglioneuroblastoma, Intermixed|9490/3
C1517445|T191|PT|C42058|NCI|Ganglioneuroblastoma, Nodular|9490/3
C0206718|T191|PT|C3790|NCI_CDISC|GANGLIONEUROBLASTOMA, MALIGNANT|9490/3
C0206718|T191|PT|C3790|NCI_CPTAC|Ganglioneuroblastoma|9490/3
C0206718|T191|DN|C3790|NCI_CTRP|Ganglioneuroblastoma|9490/3
C0206718|T191|PT|CDR0000761751|PDQ|ganglioneuroblastoma|9490/3
C0206718|T191|SY|CDR0000761751|PDQ|ganglioneuroblastoma, malignant|9490/3
C0206718|T191|PT|BBc01|RCD|Ganglioneuroblastoma|9490/3
C0206718|T191|PT|116381000119105|SNOMEDCT_US|Ganglioneuroblastoma|9490/3
C0206718|T191|PT|69515008|SNOMEDCT_US|Ganglioneuroblastoma|9490/3
C1517444|T191|SY|822951003|SNOMEDCT_US|Ganglioneuroblastoma, intermixed|9490/3
C1517445|T191|SY|822950002|SNOMEDCT_US|Ganglioneuroblastoma, nodular|9490/3
C1517444|T191|PT|822951003|SNOMEDCT_US|Intermixed ganglioneuroblastoma|9490/3
C1517445|T191|PT|822950002|SNOMEDCT_US|Nodular ganglioneuroblastoma|9490/3
C0334595|T191|PT|HP:0025151|HPO|Ganglioneuromatosis|9491/0
C0334595|T191|PT|MTHU030277|ICPC2ICD10ENG|ganglioneuromatosis|9491/0
C0334595|T191|PT|C66804|NCI|Ganglioneuromatosis|9491/0
C0334595|T191|PT|BBc02|RCD|Ganglioneuromatosis|9491/0
C0334595|T191|PT|12060004|SNOMEDCT_US|Ganglioneuromatosis|9491/0
C0017075|T191|ET|0000004647|AOD|ganglioneuroma|9492/0
C0017075|T191|SY|0000005343|CHV|gangliocytoma|9492/0
C0017075|T191|SY|0000005343|CHV|gangliocytomas|9492/0
C0017075|T191|PT|0000005343|CHV|ganglioneuroma|9492/0
C0017075|T191|SY|0000005343|CHV|ganglioneuromas|9492/0
C0017075|T191|SY|NOCODE|DXP|GANGLIONEUROFIBROMA|9492/0
C0017075|T191|DI|U000693|DXP|GANGLIONEUROMA|9492/0
C0017075|T191|PT|HP:0003005|HPO|Ganglioneuroma|9492/0
C0017075|T191|PT|MTHU030261|ICPC2ICD10ENG|gangliocytoma|9492/0
C0017075|T191|PT|MTHU030278|ICPC2ICD10ENG|ganglioneuroma|9492/0
C0017075|T191|LA|LA26521-7|LNC|Ganglioneuroma|9492/0
C0017075|T191|LLT|10017700|MDR|Gangliocytoma|9492/0
C0017075|T191|LLT|10017709|MDR|Ganglioneuroma|9492/0
C0017075|T191|PT|10017709|MDR|Ganglioneuroma|9492/0
C0017075|T191|ET|D005729|MSH|Gangliocytoma|9492/0
C0017075|T191|PM|D005729|MSH|Gangliocytomas|9492/0
C0017075|T191|MH|D005729|MSH|Ganglioneuroma|9492/0
C0017075|T191|PM|D005729|MSH|Ganglioneuromas|9492/0
C0017075|T191|PN|NOCODE|MTH|Ganglioneuroma|9492/0
C0017075|T191|SY|TCGA|NCI|Gangliocytoma|9492/0
C0017075|T191|PT|C6934|NCI|Gangliocytoma|9492/0
C0017075|T191|PT|C3049|NCI|Ganglioneuroma|9492/0
C0017075|T191|PT|C3049|NCI_CDISC|GANGLIONEUROMA, BENIGN|9492/0
C0017075|T191|SY|C3049|NCI_CDISC|Neural Crest Tumor, Benign|9492/0
C0017075|T191|DN|C3049|NCI_CTRP|Ganglioneuroma|9492/0
C0017075|T191|PT|X77pU|RCD|Gangliocytoma|9492/0
C0017075|T191|PT|BBc00|RCD|Ganglioneuroma|9492/0
C0017075|T191|IS|53801007|SNOMEDCT_US|Gangliocytoma|9492/0
C0017075|T191|PT|128919000|SNOMEDCT_US|Gangliocytoma|9492/0
C0017075|T191|PT|116371000119107|SNOMEDCT_US|Ganglioneuroma|9492/0
C0017075|T191|OAP|189929007|SNOMEDCT_US|Ganglioneuroma|9492/0
C0017075|T191|PT|53801007|SNOMEDCT_US|Ganglioneuroma|9492/0
C0391826|T191|PT|HP:0500009|HPO|Dysplastic gangliocytoma of the cerebellum|9493/0
C0391826|T191|ET|HP:0500009|HPO|LDD|9493/0
C0391826|T191|ET|HP:0500009|HPO|Lhermitte-Duclos disease|9493/0
C0391826|T191|PT|355033|MEDCIN|Lhermitte-Duclos disease|9493/0
C0391826|T191|SY|355033|MEDCIN|neoplasm of head intracranial tumor lhermitte-duclos disease|9493/0
C0391826|T191|PM|D006223|MSH|Cerebellum Dysplastic Gangliocytoma|9493/0
C0391826|T191|PM|D006223|MSH|Cerebellum Dysplastic Gangliocytomas|9493/0
C0391826|T191|ET|D006223|MSH|Dysplastic Gangliocytoma of Cerebellum|9493/0
C0391826|T191|ET|D006223|MSH|Dysplastic Gangliocytoma of the Cerebellum|9493/0
C0391826|T191|PM|D006223|MSH|Lhermitte Duclos Disease|9493/0
C0391826|T191|PEP|D006223|MSH|Lhermitte-Duclos Disease|9493/0
C0391826|T191|PN|NOCODE|MTH|Lhermitte-Duclos disease|9493/0
C0391826|T191|PT|C8419|NCI|Dysplastic Cerebellar Gangliocytoma|9493/0
C0391826|T191|SY|C8419|NCI|Dysplastic Gangliocytoma of Cerebellum|9493/0
C0391826|T191|SY|C8419|NCI|Dysplastic Gangliocytoma of the Cerebellum|9493/0
C0391826|T191|SY|C8419|NCI|Lhermitte-Duclos Disease|9493/0
C0391826|T191|SY|67944007|SNOMEDCT_US|Dysplastic cerebellar gangliocytoma|9493/0
C0391826|T191|PT|67944007|SNOMEDCT_US|Lhermitte-Duclos disease|9493/0
C0027819|T191|ET|0000004648|AOD|neuroblastoma|9500/3
C0027819|T191|PT|0000008628|CHV|neuroblastoma|9500/3
C0027819|T191|SY|0000008628|CHV|neuroblastomas|9500/3
C0027819|T191|PT|NOCODE|COSTAR|Neuroblastoma|9500/3
C0027819|T191|PT|2012-7126|CSP|neuroblastoma|9500/3
C0027819|T191|GT|NEOPL|CST|NEUROBLASTOMA|9500/3
C0027819|T191|DI|U001281|DXP|NEUROBLASTOMA|9500/3
C2239230|T191|SY|NOCODE|DXP|NEUROBLASTOMA SYMPATHICUM|9500/3
C2239230|T191|SY|NOCODE|DXP|SYMPATHICOBLASTOMA|9500/3
C2239230|T191|SY|NOCODE|DXP|SYMPATHICOGONIOMA|9500/3
C0027819|T191|SY|HP:0003006|HPO|Cancer of early nerve cells|9500/3
C0027819|T191|PT|HP:0003006|HPO|Neuroblastoma|9500/3
C0027819|T191|PT|MTHU052494|ICPC2ICD10ENG|neuroblastoma; unspecified site|9500/3
C0027819|T191|PT|U003183|LCH|Neuroblastoma|9500/3
C0027819|T191|PT|sh85091115|LCH_NW|Neuroblastoma|9500/3
C0027819|T191|LLT|10029260|MDR|Neuroblastoma|9500/3
C0027819|T191|PT|10029260|MDR|Neuroblastoma|9500/3
C0027819|T191|LLT|10029261|MDR|Neuroblastoma NOS|9500/3
C0027819|T191|PT|36085|MEDCIN|neuroblastoma|9500/3
C0027819|T191|PT|1240|MEDLINEPLUS|Neuroblastoma|9500/3
C0027819|T191|MH|D009447|MSH|Neuroblastoma|9500/3
C0027819|T191|PM|D009447|MSH|Neuroblastomas|9500/3
C0027819|T191|PN|NOCODE|MTH|Neuroblastoma|9500/3
C0027819|T191|PT|C3270|NCI|Neuroblastoma|9500/3
C0027819|T191|SY|TCGA|NCI|Neuroblastoma|9500/3
C0027819|T191|SY|C3270|NCI_CDISC|Neural Crest Tumor, Malignant|9500/3
C0027819|T191|PT|C3270|NCI_CDISC|NEUROBLASTOMA, MALIGNANT|9500/3
C0027819|T191|PT|C3270|NCI_CPTAC|Neuroblastoma|9500/3
C0027819|T191|PT|10029261|NCI_CTEP-SDC|Neuroblastoma|9500/3
C0027819|T191|PT|C3270|NCI_CTRP|Neuroblastoma|9500/3
C0027819|T191|DN|C3270|NCI_CTRP|Neuroblastoma|9500/3
C0027819|T191|PT|CDR0000045418|NCI_NCI-GLOSS|neuroblastoma|9500/3
C0027819|T191|PT|C3270|NCI_NICHD|Neuroblastoma|9500/3
C0027819|T191|PSC|CDR0000042067|PDQ|neuroblastoma|9500/3
C0027819|T191|ET|CDR0000042067|PDQ|Neuroblastoma|9500/3
C2239230|T191|OP|X77pZ|RCD|Sympathicoblastoma|9500/3
C0027819|T191|OP|XE1wc|RCDSY|Neuroblastoma NOS|9500/3
C2239230|T191|IS|X77pZ|RCDSY|Sympathicogonioma|9500/3
C2239230|T191|IS|X77pZ|RCDSY|Sympathogonioma|9500/3
C0027819|T191|SY|87364003|SNOMEDCT_US|NB - Neuroblastoma|9500/3
C0027819|T191|PT|432328008|SNOMEDCT_US|Neuroblastoma|9500/3
C0027819|T191|PT|87364003|SNOMEDCT_US|Neuroblastoma|9500/3
C0027819|T191|IS|87364003|SNOMEDCT_US|Neuroblastoma, NOS|9500/3
C2239230|T191|PT|253075001|SNOMEDCT_US|Sympathicoblastoma|9500/3
C2239230|T191|SY|87364003|SNOMEDCT_US|Sympathicoblastoma|9500/3
C2239230|T191|SY|253075001|SNOMEDCT_US|Sympathicogonioma|9500/3
C2239230|T191|SY|253075001|SNOMEDCT_US|Sympathogonioma|9500/3
C0027819|T191|PT|1130|WHO|NEUROBLASTOMA|9500/3
C1879808|T191|PT|C66807|NCI|Benign Intraocular Medulloepithelioma|9501/0
C1266182|T191|SY|128910001|SNOMEDCT_US|Diktyoma, benign|9501/0
C1266182|T191|PT|128910001|SNOMEDCT_US|Medulloepithelioma, benign|9501/0
C0334596|T191|PT|0000030012|CHV|medulloepithelioma|9501/3
C0334596|T191|SY|0000030012|CHV|medulloepitheliomas|9501/3
C0334596|T191|PT|HP:0030071|HPO|Medulloepithelioma|9501/3
C0334596|T191|PT|271565|MEDCIN|malignant medulloepithelioma|9501/3
C0334596|T191|SY|271565|MEDCIN|medulloepithelioma|9501/3
C0334596|T191|PEP|D018242|MSH|Medulloepithelioma|9501/3
C0334596|T191|PM|D018242|MSH|Medulloepitheliomas|9501/3
C0334596|T191|PN|NOCODE|MTH|Medulloepithelioma|9501/3
C0334596|T191|SY|C4327|NCI|Central Nervous System Medulloepithelioma|9501/3
C0334596|T191|PT|C4327|NCI|Medulloepithelioma|9501/3
C0334596|T191|OP|C66808|NCI|Medulloepithelioma Not Otherwise Specified|9501/3
C0334596|T191|PT|C66808|NCI|Medulloepithelioma Not Otherwise Specified|9501/3
C0334596|T191|SY|C4327|NCI|Medulloepithelioma, Central Nervous System|9501/3
C0334596|T191|OP|C66808|NCI|Medulloepithelioma, NOS|9501/3
C0334596|T191|DN|C4327|NCI_CTRP|Medulloepithelioma|9501/3
C0334596|T191|PT|C4327|NCI_NICHD|Medulloepithelioma|9501/3
C0334596|T191|PT|Xa99F|RCD|Medulloepithelioma|9501/3
C0457180|T191|PT|Xa0aG|RCD|Nonteratoid medulloepithelioma|9501/3
C0334596|T191|OP|BBc2.|RCDSY|Medulloepithelioma NOS|9501/3
C0334596|T191|SY|39005004|SNOMEDCT_US|Diktyoma|9501/3
C0334596|T191|SY|39005004|SNOMEDCT_US|Diktyoma, malignant|9501/3
C0334596|T191|PT|715903004|SNOMEDCT_US|Medulloepithelioma|9501/3
C0334596|T191|PT|39005004|SNOMEDCT_US|Medulloepithelioma|9501/3
C0334596|T191|IS|39005004|SNOMEDCT_US|Medulloepithelioma, NOS|9501/3
C0457180|T191|PT|277985001|SNOMEDCT_US|Nonteratoid medulloepithelioma|9501/3
C1879809|T191|PT|C66809|NCI|Benign Intraocular Teratoid Medulloepithelioma|9502/0
C1266183|T191|PT|128911002|SNOMEDCT_US|Teratoid medulloepithelioma, benign|9502/0
C0334597|T191|PT|271566|MEDCIN|teratoid medulloepithelioma|9502/3
C1881244|T191|PT|C66810|NCI|Intraocular Teratoid Medulloepithelioma|9502/3
C0334597|T191|PT|BBc3.|RCD|Teratoid medulloepithelioma|9502/3
C0334597|T191|PT|88591002|SNOMEDCT_US|Teratoid medulloepithelioma|9502/3
C0206663|T191|SY|0000042698|CHV|neuroectodermal primitive tumors|9503/3
C0206663|T191|SY|0000021005|CHV|pnet|9503/3
C0206663|T191|SY|0000021005|CHV|primitive neuroectodermal tumor|9503/3
C0206663|T191|PT|0000042698|CHV|primitive neuroectodermal tumors|9503/3
C0206663|T191|SY|0000021005|CHV|primitive neuroectodermal tumors|9503/3
C0206663|T191|SY|0000021005|CHV|primitive neuroectodermal tumour|9503/3
C0206663|T191|PT|HP:0030065|HPO|Primitive neuroectodermal tumor|9503/3
C0206663|T191|PT|MTHU052504|ICPC2ICD10ENG|neuroectodermal; tumor, primitive, unspecified site|9503/3
C0206663|T191|PT|MTHU061687|ICPC2ICD10ENG|primitive; neuroectodermal tumor, unspecified site|9503/3
C0206663|T191|PT|MTHU077105|ICPC2ICD10ENG|tumor; neuroectodermal, primitive, unspecified site|9503/3
C0206663|T191|LLT|10057849|MDR|Primitive neuroectodermal tumor|9503/3
C0206663|T191|MTH_PT|10057846|MDR|Primitive neuroectodermal tumor|9503/3
C0206663|T191|PT|10057846|MDR|Primitive neuroectodermal tumour|9503/3
C0206663|T191|LLT|10057846|MDR|Primitive neuroectodermal tumour|9503/3
C0206663|T191|PT|271567|MEDCIN|neuroepithelioma|9503/3
C0206663|T191|DEV|D018242|MSH|NEOPL PRIMITIVE NEUROEPITHELIAL|9503/3
C0206663|T191|PM|D018242|MSH|Neoplasm, Primitive Neuroepithelial|9503/3
C0206663|T191|ET|D018242|MSH|Neoplasms, Primitive Neuroepithelial|9503/3
C0206663|T191|ET|D018242|MSH|Neuroectodermal Tumor, Primitive|9503/3
C0206663|T191|MH|D018242|MSH|Neuroectodermal Tumors, Primitive|9503/3
C0206663|T191|DEV|D018242|MSH|NEUROEPITHELIAL NEOPL PRIMITIVE|9503/3
C0206663|T191|PM|D018242|MSH|Neuroepithelial Neoplasm, Primitive|9503/3
C0206663|T191|ET|D018242|MSH|Neuroepithelial Neoplasms, Primitive|9503/3
C0206663|T191|PM|D018242|MSH|Neuroepithelial Tumor, Primitive|9503/3
C0206663|T191|ET|D018242|MSH|Neuroepithelial Tumors, Primitive|9503/3
C0206663|T191|ET|D018242|MSH|PNET|9503/3
C0206663|T191|PM|D018242|MSH|PNETs|9503/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroectodermal Tumor|9503/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroectodermal Tumors|9503/3
C0206663|T191|DEV|D018242|MSH|PRIMITIVE NEUROEPITHELIAL NEOPL|9503/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroepithelial Neoplasm|9503/3
C0206663|T191|ET|D018242|MSH|Primitive Neuroepithelial Neoplasms|9503/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroepithelial Tumor|9503/3
C0206663|T191|PM|D018242|MSH|Primitive Neuroepithelial Tumors|9503/3
C0206663|T191|PM|D018242|MSH|Tumor, Primitive Neuroectodermal|9503/3
C0206663|T191|PM|D018242|MSH|Tumor, Primitive Neuroepithelial|9503/3
C0206663|T191|PM|D018242|MSH|Tumors, Primitive Neuroectodermal|9503/3
C0206663|T191|PM|D018242|MSH|Tumors, Primitive Neuroepithelial|9503/3
C0206663|T191|PN|NOCODE|MTH|Neuroectodermal Tumor, Primitive|9503/3
C0206663|T191|SY|C3716|NCI|Neuroectodermal Neoplasm|9503/3
C0206663|T191|SY|C3716|NCI|Neuroectodermal Tumor|9503/3
C0206663|T191|SY|C3716|NCI|Neuroepithelioma|9503/3
C0206663|T191|AB|C3716|NCI|PNET|9503/3
C0206663|T191|SY|C3716|NCI|Primitive Neuroectodermal Neoplasm|9503/3
C0206663|T191|PT|C3716|NCI|Primitive Neuroectodermal Tumor|9503/3
C0206663|T191|SY|TCGA|NCI|Primitive Neuroectodermal Tumor|9503/3
C0206663|T191|PT|C3716|NCI_CPTAC|Primitive Neuroectodermal Tumor|9503/3
C0206663|T191|PT|C3716|NCI_CTRP|Primitive Neuroectodermal Tumor|9503/3
C0206663|T191|PT|CDR0000045952|NCI_NCI-GLOSS|neuroectodermal tumor|9503/3
C0206663|T191|PT|CDR0000383924|NCI_NCI-GLOSS|PNET|9503/3
C0206663|T191|PT|CDR0000383920|NCI_NCI-GLOSS|primitive neuroectodermal tumor|9503/3
C0206663|T191|SY|CDR0000039466|PDQ|PNET|9503/3
C0206663|T191|PT|Xa99H|RCD|Neuroepithelioma|9503/3
C0206663|T191|AB|X77pa|RCD|PNET - Primit neuroect tumour|9503/3
C0206663|T191|SY|X77pa|RCD|PNET - Primitive neuroectodermal tumour|9503/3
C0206663|T191|AB|X77pa|RCD|Primitive neuroectodermal tum|9503/3
C0206663|T191|PT|X77pa|RCD|Primitive neuroectodermal tumour|9503/3
C0206663|T191|AB|X77pa|RCDAE|PNET - Primit neuroect tumor|9503/3
C0206663|T191|SY|X77pa|RCDAE|PNET - Primitive neuroectodermal tumor|9503/3
C0206663|T191|PT|X77pa|RCDAE|Primitive neuroectodermal tumor|9503/3
C0206663|T191|OP|BBc4.|RCDSY|Neuroepithelioma NOS|9503/3
C0206663|T191|AB|X77pa|RCDSY|Primit neuroectodermal tumr|9503/3
C0206663|T191|PT|55045006|SNOMEDCT_US|Neuroepithelioma|9503/3
C0206663|T191|IS|55045006|SNOMEDCT_US|Neuroepithelioma, NOS|9503/3
C0206663|T191|SY|39781001|SNOMEDCT_US|PNET|9503/3
C0206663|T191|SY|39781001|SNOMEDCT_US|PNET - Primitive neuroectodermal tumor|9503/3
C0206663|T191|SYGB|39781001|SNOMEDCT_US|PNET - Primitive neuroectodermal tumour|9503/3
C0206663|T191|OAP|189925001|SNOMEDCT_US|Primitive neuroectodermal tumor|9503/3
C0206663|T191|PT|699028006|SNOMEDCT_US|Primitive neuroectodermal tumor|9503/3
C0206663|T191|PT|39781001|SNOMEDCT_US|Primitive neuroectodermal tumor|9503/3
C0206663|T191|PTGB|699028006|SNOMEDCT_US|Primitive neuroectodermal tumour|9503/3
C0206663|T191|PTGB|39781001|SNOMEDCT_US|Primitive neuroectodermal tumour|9503/3
C0206663|T191|OAP|189925001|SNOMEDCT_US|Primitive neuroectodermal tumour|9503/3
C0206663|T191|OF|189925001|SNOMEDCT_US|Primitive neuroectodermal tumour|9503/3
C0334598|T191|PT|271568|MEDCIN|spongioneuroblastoma|9504/3
C0334598|T191|OP|C66811|NCI|Spongioneuroblastoma|9504/3
C0334598|T191|PT|C66811|NCI|Spongioneuroblastoma|9504/3
C0334598|T191|OP|BBc5.|RCD|Spongioneuroblastoma|9504/3
C0334598|T191|PT|64059005|SNOMEDCT_US|Spongioneuroblastoma|9504/3
C0206716|T191|PT|0000021042|CHV|ganglioglioma|9505/1
C0206716|T191|SY|0000021042|CHV|gangliogliomas|9505/1
C0206716|T191|SY|0000021042|CHV|glioneuroma|9505/1
C0206716|T191|SY|0000021042|CHV|neuroastrocytoma|9505/1
C0206716|T191|ET|2012-6589|CSP|ganglioglioma|9505/1
C0206716|T191|PT|10017701|MDR|Ganglioglioma|9505/1
C0206716|T191|LLT|10017701|MDR|Ganglioglioma|9505/1
C0206716|T191|MH|D018303|MSH|Ganglioglioma|9505/1
C0206716|T191|PM|D018303|MSH|Gangliogliomas|9505/1
C0206716|T191|PN|NOCODE|MTH|Ganglioglioma|9505/1
C0206716|T191|PT|C3788|NCI|Ganglioglioma|9505/1
C0206716|T191|SY|TCGA|NCI|Ganglioglioma|9505/1
C0206716|T191|PT|BBc6.|RCD|Ganglioglioma|9505/1
C0206716|T191|SY|89880005|SNOMEDCT_US|Ganglioglioma|9505/1
C0206716|T191|PT|87191000119100|SNOMEDCT_US|Ganglioglioma|9505/1
C0206716|T191|PT|89880005|SNOMEDCT_US|Ganglioglioma, no ICD-O subtype|9505/1
C0206716|T191|SY|89880005|SNOMEDCT_US|Ganglioglioma, no International Classification of Diseases for Oncology subtype|9505/1
C0206716|T191|SY|89880005|SNOMEDCT_US|Glioneuroma|9505/1
C0206716|T191|SY|89880005|SNOMEDCT_US|Neuroastrocytoma|9505/1
C0431112|T191|PT|271569|MEDCIN|anaplastic ganglioglioma|9505/3
C0431112|T191|PN|NOCODE|MTH|Anaplastic ganglioglioma|9505/3
C0431112|T191|PT|C4717|NCI|Anaplastic Ganglioglioma|9505/3
C0431112|T191|PT|X77pX|RCD|Anaplastic ganglioglioma|9505/3
C0431112|T191|OAP|134212004|SNOMEDCT_US|Anaplastic ganglioglioma|9505/3
C0431112|T191|PT|128912009|SNOMEDCT_US|Ganglioglioma, anaplastic|9505/3
C0206719|T191|SY|0000021045|CHV|central neurocytoma|9506/1
C1370507|T191|SY|0000021045|CHV|cerebellar liponeurocytoma|9506/1
C0206719|T191|PM|D018306|MSH|Central Neurocytoma|9506/1
C0206719|T191|PM|D018306|MSH|Central Neurocytomas|9506/1
C0206719|T191|PEP|D018306|MSH|Neurocytoma, Central|9506/1
C0206719|T191|PM|D018306|MSH|Neurocytomas, Central|9506/1
C0206719|T191|PN|NOCODE|MTH|Central Neurocytoma|9506/1
C1370507|T191|PN|NOCODE|MTH|Cerebellar Liponeurocytoma|9506/1
C0206719|T191|PT|C3791|NCI|Central Neurocytoma|9506/1
C1370507|T191|PT|C6905|NCI|Cerebellar Liponeurocytoma|9506/1
C2985175|T191|PT|C92555|NCI|Extraventricular Neurocytoma|9506/1
C1370507|T191|SY|C6905|NCI|Lipomatous Medulloblastoma|9506/1
C0206719|T191|PT|Xa99I|RCD|Central neurocytoma|9506/1
C0206719|T191|OAP|302832007|SNOMEDCT_US|Central neurocytoma|9506/1
C0206719|T191|PT|128858006|SNOMEDCT_US|Central neurocytoma|9506/1
C0206719|T191|SY|128858006|SNOMEDCT_US|Central neurocytoma - histology|9506/1
C1370507|T191|IS|128858006|SNOMEDCT_US|Cerebellar liponeurocytoma|9506/1
C1370507|T191|PT|734134003|SNOMEDCT_US|Cerebellar liponeurocytoma|9506/1
C1370507|T191|PT|716592003|SNOMEDCT_US|Cerebellar liponeurocytoma|9506/1
C2985175|T191|PT|716787002|SNOMEDCT_US|Extraventricular neurocytoma|9506/1
C2985175|T191|PT|716179006|SNOMEDCT_US|Extraventricular neurocytoma|9506/1
C0206719|T191|SY|128858006|SNOMEDCT_US|Lipomatous medulloblastoma|9506/1
C1370507|T191|SY|716592003|SNOMEDCT_US|Liponeurocytoma of cerebellum|9506/1
C0206719|T191|SY|128858006|SNOMEDCT_US|Medullocytoma|9506/1
C0206719|T191|SY|128858006|SNOMEDCT_US|Neurolipocytoma|9506/1
C0334599|T191|PT|C4328|NCI|Pacinian Neurofibroma|9507/0
C0334599|T191|SY|BBc8.|RCD|Pacinian neurofibroma|9507/0
C0334599|T191|PT|BBc8.|RCD|Pacinian tumour|9507/0
C0334599|T191|PT|BBc8.|RCDAE|Pacinian tumor|9507/0
C0334599|T191|SY|4230004|SNOMEDCT_US|Pacinian neurofibroma|9507/0
C0334599|T191|PT|404033003|SNOMEDCT_US|Pacinian neurofibroma|9507/0
C0334599|T191|PT|4230004|SNOMEDCT_US|Pacinian tumor|9507/0
C0334599|T191|PTGB|4230004|SNOMEDCT_US|Pacinian tumour|9507/0
C1266184|T191|PN|NOCODE|MTH|Atypical Teratoid Rhabdoid Tumor|9508/3
C1266184|T191|AB|C6906|NCI|AT/RT|9508/3
C1266184|T191|PT|C6906|NCI|Atypical Teratoid/Rhabdoid Tumor|9508/3
C1266184|T191|SY|TCGA|NCI|Atypical Teratoid/Rhabdoid Tumor|9508/3
C1266184|T191|SY|C6906|NCI|Central Nervous System Rhabdoid Neoplasm|9508/3
C1266184|T191|SY|C6906|NCI|Central Nervous System Rhabdoid Tumor|9508/3
C1266184|T191|SY|C6906|NCI|CNS Rhabdoid Neoplasm|9508/3
C1266184|T191|SY|C6906|NCI|CNS Rhabdoid Tumor|9508/3
C1266184|T191|SY|C6906|NCI|Malignant Brain Rhabdoid Neoplasm|9508/3
C1266184|T191|SY|C6906|NCI|Malignant Brain Rhabdoid Tumor|9508/3
C1266184|T191|SY|C6906|NCI|Malignant Rhabdoid Neoplasm of Brain|9508/3
C1266184|T191|SY|C6906|NCI|Malignant Rhabdoid Neoplasm of the Brain|9508/3
C1266184|T191|SY|C6906|NCI|Malignant Rhabdoid Tumor of Brain|9508/3
C1266184|T191|SY|C6906|NCI|Malignant Rhabdoid Tumor of the Brain|9508/3
C1266184|T191|SY|C6906|NCI|Primary Malignant Brain Rhabdoid Neoplasm|9508/3
C1266184|T191|SY|C6906|NCI|Primary Malignant Brain Rhabdoid Tumor|9508/3
C1266184|T191|SY|C6906|NCI|Primary Malignant Rhabdoid Neoplasm of Brain|9508/3
C1266184|T191|SY|C6906|NCI|Primary Malignant Rhabdoid Neoplasm of the Brain|9508/3
C1266184|T191|SY|C6906|NCI|Primary Malignant Rhabdoid Tumor of Brain|9508/3
C1266184|T191|SY|C6906|NCI|Primary Malignant Rhabdoid Tumor of the Brain|9508/3
C1266184|T191|SY|C6906|NCI|Rhabdoid Neoplasm of Central Nervous System|9508/3
C1266184|T191|SY|C6906|NCI|Rhabdoid Neoplasm of CNS|9508/3
C1266184|T191|SY|C6906|NCI|Rhabdoid Neoplasm of the Central Nervous System|9508/3
C1266184|T191|SY|C6906|NCI|Rhabdoid Neoplasm of the CNS|9508/3
C1266184|T191|SY|C6906|NCI|Rhabdoid Tumor of Central Nervous System|9508/3
C1266184|T191|SY|C6906|NCI|Rhabdoid Tumor of CNS|9508/3
C1266184|T191|SY|C6906|NCI|Rhabdoid Tumor of the Central Nervous System|9508/3
C1266184|T191|SY|C6906|NCI|Rhabdoid Tumor of the CNS|9508/3
C1266184|T191|PT|C6906|NCI_CPTAC|Atypical Teratoid/Rhabdoid Tumor|9508/3
C1266184|T191|PT|10065870|NCI_CTEP-SDC|Atypical teratoid/rhabdoid tumor|9508/3
C1266184|T191|PT|CDR0000584380|NCI_NCI-GLOSS|AT/RT|9508/3
C1266184|T191|PT|CDR0000584379|NCI_NCI-GLOSS|ATT/RHT|9508/3
C1266184|T191|PT|CDR0000285639|NCI_NCI-GLOSS|atypical teratoid/rhabdoid tumor|9508/3
C1266184|T191|PT|128792003|SNOMEDCT_US|Atypical teratoid/rhabdoid tumor|9508/3
C1266184|T191|PTGB|128792003|SNOMEDCT_US|Atypical teratoid/rhabdoid tumour|9508/3
C4518368|T191|PT|734068006|SNOMEDCT_US|Embryonal central nervous system neoplasm with rhabdoid feature|9508/3
C4331262|T191|SY|HP:0025171|HPO|Rosette-forming glioneuronal neoplasm|9509/1
C4331262|T191|PT|HP:0025171|HPO|Rosette-forming glioneuronal tumor|9509/1
C2347979|T191|ET|HP:0025171|HPO|Rosette-forming glioneuronal tumor of the fourth ventricle|9509/1
C4331262|T191|SY|HP:0025171|HPO|Rosette-forming glioneuronal tumour|9509/1
C2985174|T191|PT|C92554|NCI|Papillary Glioneuronal Tumor|9509/1
C4331262|T191|AB|C129431|NCI|RGNT|9509/1
C4331262|T191|PT|C129431|NCI|Rosette-Forming Glioneuronal Tumor|9509/1
C2347979|T191|PT|C67559|NCI|Rosette-Forming Glioneuronal Tumor of the Fourth Ventricle|9509/1
C2985174|T191|PT|450902001|SNOMEDCT_US|Papillary glioneuronal tumor|9509/1
C2985174|T191|PTGB|450902001|SNOMEDCT_US|Papillary glioneuronal tumour|9509/1
C4331262|T191|PT|733906003|SNOMEDCT_US|Rosette-forming glioneuronal neoplasm|9509/1
C4331262|T191|PT|770682007|SNOMEDCT_US|Rosette-forming glioneuronal neoplasm|9509/1
C4331262|T191|SY|770682007|SNOMEDCT_US|Rosette-forming glioneuronal tumor|9509/1
C4331262|T191|SY|733906003|SNOMEDCT_US|Rosette-forming glioneuronal tumor|9509/1
C4331262|T191|SYGB|770682007|SNOMEDCT_US|Rosette-forming glioneuronal tumour|9509/1
C4331262|T191|SYGB|733906003|SNOMEDCT_US|Rosette-forming glioneuronal tumour|9509/1
C0346396|T191|SY|365990|MEDCIN|eye neoplasm benign retinocytoma|9510/0
C0346396|T191|PT|365990|MEDCIN|Retinocytoma|9510/0
C0346396|T191|PN|NOCODE|MTH|Retinoma|9510/0
C0346396|T191|PT|C66812|NCI|Retinocytoma|9510/0
C0346396|T191|SY|X78c9|RCD|Adenoma of retinal pigment epithelium|9510/0
C0346396|T191|AB|X78c9|RCD|Adenoma ret pigment epithelium|9510/0
C0346396|T191|SY|X78c8|RCD|Retinocytoma|9510/0
C0346396|T191|PT|X78c9|RCD|Retinoma|9510/0
C0346396|T191|SY|255027009|SNOMEDCT_US|Adenoma of retinal pigment epithelium|9510/0
C0346396|T191|PT|416864007|SNOMEDCT_US|Retinocytoma|9510/0
C0346396|T191|PT|128913004|SNOMEDCT_US|Retinocytoma|9510/0
C0346396|T191|IS|255026000|SNOMEDCT_US|Retinocytoma|9510/0
C0346396|T191|PT|255027009|SNOMEDCT_US|Retinoma|9510/0
C0346396|T191|IS|416864007|SNOMEDCT_US|Retinoma|9510/0
C0035335|T191|ET|0000004646|AOD|retinoblastoma|9510/3
C0035335|T191|PT|0041900|CCPSS|RETINOBLASTOMA|9510/3
C0035335|T191|SY|0000010813|CHV|disorders retinoblastoma|9510/3
C0035335|T191|PT|0000010813|CHV|retinoblastoma|9510/3
C0035335|T191|SY|0000010813|CHV|retinoblastomas|9510/3
C0035335|T191|PT|2018-3452|CSP|retinoblastoma|9510/3
C0035335|T191|SY|NOCODE|DXP|RETINA, GLIOMA|9510/3
C0035335|T191|DI|U001674|DXP|RETINOBLASTOMA|9510/3
C0035335|T191|PT|HP:0009919|HPO|Retinoblastoma|9510/3
C0035335|T191|PT|MTHU064505|ICPC2ICD10ENG|retinoblastoma|9510/3
C0035335|T191|PTN|F74006|ICPC2P|retinoblastoma|9510/3
C0035335|T191|PT|F74006|ICPC2P|Retinoblastoma|9510/3
C0035335|T191|PT|U004110|LCH|Retinoblastoma|9510/3
C0035335|T191|PT|sh85113337|LCH_NW|Retinoblastoma|9510/3
C0035335|T191|LA|LA16305-7|LNC|Retinoblastoma|9510/3
C0035335|T191|LLT|10038916|MDR|Retinoblastoma|9510/3
C0035335|T191|PT|10038916|MDR|Retinoblastoma|9510/3
C0035335|T191|LLT|10038918|MDR|Retinoblastoma NOS|9510/3
C0035335|T191|PT|235049|MEDCIN|malignant retinoblastoma of eye|9510/3
C0035335|T191|PT|38366|MEDCIN|retinoblastoma|9510/3
C0035335|T191|ET|491|MEDLINEPLUS|Retinoblastoma|9510/3
C0035335|T191|PM|D012175|MSH|Cancer, Retinoblastoma Eye|9510/3
C0035335|T191|PM|D012175|MSH|Cancers, Retinoblastoma Eye|9510/3
C0035335|T191|ET|D012175|MSH|Eye Cancer, Retinoblastoma|9510/3
C0035335|T191|PM|D012175|MSH|Eye Cancers, Retinoblastoma|9510/3
C0035335|T191|ET|D012175|MSH|Glioblastoma, Retinal|9510/3
C0035335|T191|PM|D012175|MSH|Glioblastomas, Retinal|9510/3
C0035335|T191|ET|D012175|MSH|Glioma, Retinal|9510/3
C0035335|T191|PM|D012175|MSH|Gliomas, Retinal|9510/3
C0035335|T191|ET|D012175|MSH|Neuroblastoma, Retinal|9510/3
C0035335|T191|PM|D012175|MSH|Neuroblastomas, Retinal|9510/3
C0035335|T191|PM|D012175|MSH|Retinal Glioblastoma|9510/3
C0035335|T191|PM|D012175|MSH|Retinal Glioblastomas|9510/3
C0035335|T191|PM|D012175|MSH|Retinal Glioma|9510/3
C0035335|T191|PM|D012175|MSH|Retinal Gliomas|9510/3
C0035335|T191|PM|D012175|MSH|Retinal Neuroblastoma|9510/3
C0035335|T191|PM|D012175|MSH|Retinal Neuroblastomas|9510/3
C0035335|T191|MH|D012175|MSH|Retinoblastoma|9510/3
C0035335|T191|PM|D012175|MSH|Retinoblastoma Eye Cancer|9510/3
C0035335|T191|PM|D012175|MSH|Retinoblastoma Eye Cancers|9510/3
C0035335|T191|PM|D012175|MSH|Retinoblastomas|9510/3
C0035335|T191|PN|NOCODE|MTH|Retinoblastoma|9510/3
C0035335|T191|SY|C6956|NCI|Neuroblastoma of Retina|9510/3
C0035335|T191|SY|C6956|NCI|Neuroblastoma of the Retina|9510/3
C0035335|T191|AB|C7541|NCI|RB|9510/3
C0035335|T191|PT|C6956|NCI|Retinal Neuroblastoma|9510/3
C0035335|T191|PT|C7541|NCI|Retinoblastoma|9510/3
C0035335|T191|SY|C7541|NCI_CDISC|RB|9510/3
C0035335|T191|PT|C7541|NCI_CDISC|RETINOBLASTOMA, MALIGNANT|9510/3
C0035335|T191|PT|C7541|NCI_CPTAC|Retinoblastoma|9510/3
C0035335|T191|PT|10038918|NCI_CTEP-SDC|Retinoblastoma|9510/3
C0035335|T191|PT|C7541|NCI_CTRP|Retinoblastoma|9510/3
C0035335|T191|DN|C7541|NCI_CTRP|Retinoblastoma|9510/3
C0035335|T191|PT|CDR0000046774|NCI_NCI-GLOSS|retinoblastoma|9510/3
C0035335|T191|PT|C7541|NCI_NICHD|Retinoblastoma|9510/3
C0035335|T191|PSC|CDR0000043733|PDQ|retinoblastoma|9510/3
C0035335|T191|ET|CDR0000043733|PDQ|Retinoblastoma|9510/3
C0035335|T191|SY|X00eS|RCD|RB - Retinoblastoma|9510/3
C0035335|T191|PT|X00eS|RCD|Retinoblastoma|9510/3
C0035335|T191|PT|XaBB5|RCD|Retinoblastoma - morphology|9510/3
C0035335|T191|OP|BBc9z|RCDSY|Retinoblastoma NOS|9510/3
C0035335|T191|OP|BBc9.|RCDSY|Retinoblastomas|9510/3
C0035335|T191|OAS|134191003|SNOMEDCT_US|RB - Retinoblastoma|9510/3
C0035335|T191|OAS|269614001|SNOMEDCT_US|Retinoblastoma|9510/3
C0035335|T191|OAP|134191003|SNOMEDCT_US|Retinoblastoma|9510/3
C0035335|T191|OAS|154553002|SNOMEDCT_US|Retinoblastoma|9510/3
C0035335|T191|PT|370967009|SNOMEDCT_US|Retinoblastoma|9510/3
C0035335|T191|OF|134191003|SNOMEDCT_US|Retinoblastoma|9510/3
C0035335|T191|PT|19906005|SNOMEDCT_US|Retinoblastoma|9510/3
C0035335|T191|SY|19906005|SNOMEDCT_US|Retinoblastoma - morphology|9510/3
C0035335|T191|IS|19906005|SNOMEDCT_US|Retinoblastoma, NOS|9510/3
C0035335|T191|PT|1682|WHO|RETINOBLASTOMA|9510/3
C0334600|T191|PT|MTHU030788|ICPC2ICD10ENG|differentiated; retinoblastoma|9511/3
C0334600|T191|PT|MTHU064506|ICPC2ICD10ENG|retinoblastoma; differentiated|9511/3
C0334600|T191|PT|235050|MEDCIN|differentiated retinoblastoma|9511/3
C0334600|T191|PT|C66813|NCI|Differentiated Retinoblastoma|9511/3
C0334600|T191|PT|BBc90|RCD|Retinoblastoma - differentiated|9511/3
C0334600|T191|AB|BBc90|RCD|Retinoblastoma-differentiated|9511/3
C0334600|T191|SY|26019009|SNOMEDCT_US|Retinoblastoma - differentiated|9511/3
C0334600|T191|PT|26019009|SNOMEDCT_US|Retinoblastoma, differentiated|9511/3
C0334601|T191|PT|MTHU064507|ICPC2ICD10ENG|retinoblastoma; undifferentiated|9512/3
C0334601|T191|PT|MTHU054663|ICPC2ICD10ENG|undifferentiated; retinoblastoma|9512/3
C0334601|T191|PT|235051|MEDCIN|undifferentiated retinoblastoma|9512/3
C0334601|T191|PT|C66814|NCI|Undifferentiated Retinoblastoma|9512/3
C0334601|T191|AB|BBc91|RCD|Retinoblastoma - undifferent|9512/3
C0334601|T191|PT|BBc91|RCD|Retinoblastoma - undifferentiated|9512/3
C0334601|T191|SY|12354007|SNOMEDCT_US|Retinoblastoma - undifferentiated|9512/3
C0334601|T191|PT|12354007|SNOMEDCT_US|Retinoblastoma, undifferentiated|9512/3
C1266185|T191|PT|235052|MEDCIN|diffuse retinoblastoma|9513/3
C1266185|T191|PT|C66815|NCI|Diffuse Retinoblastoma|9513/3
C1266185|T191|PT|128793008|SNOMEDCT_US|Retinoblastoma, diffuse|9513/3
C1266186|T191|PN|NOCODE|MTH|Retinoblastoma, spontaneously regressed|9514/1
C1266186|T191|SY|C66816|NCI|Retinoma|9514/1
C1266186|T191|PT|C66816|NCI|Spontaneously Regressing Retinoblastoma|9514/1
C1266186|T191|PT|128794002|SNOMEDCT_US|Retinoblastoma, spontaneously regressed|9514/1
C0334602|T191|PT|MTHU052519|ICPC2ICD10ENG|neurogenic olfactory; tumor|9520/3
C0334602|T191|PT|MTHU077106|ICPC2ICD10ENG|tumor; neurogenic olfactory|9520/3
C0334602|T191|PT|271570|MEDCIN|olfactory neurogenic tumor|9520/3
C0334602|T191|PT|C67155|NCI|Olfactory Neurogenic Tumor|9520/3
C0334602|T191|PT|BBcA.|RCD|Olfactory neurogenic tumour|9520/3
C0334602|T191|PT|BBcA.|RCDAE|Olfactory neurogenic tumor|9520/3
C0334602|T191|PT|53968002|SNOMEDCT_US|Olfactory neurogenic tumor|9520/3
C0334602|T191|PTGB|53968002|SNOMEDCT_US|Olfactory neurogenic tumour|9520/3
C0555201|T191|PT|MTHU027103|ICPC2ICD10ENG|esthesioneurocytoma|9521/3
C0555201|T191|PT|C67156|NCI|Olfactory Neurocytoma|9521/3
C0555201|T191|OP|BBcB.|RCD|Asthesioneurocytoma|9521/3
C0555201|T191|PTGB|46710009|SNOMEDCT_US|Aesthesioneurocytoma|9521/3
C0555201|T191|IS|46710009|SNOMEDCT_US|Asthesioneurocytoma|9521/3
C0555201|T191|PT|46710009|SNOMEDCT_US|Esthesioneurocytoma|9521/3
C0555201|T191|SY|46710009|SNOMEDCT_US|Olfactory neurocytoma|9521/3
C0206717|T191|PT|0000021043|CHV|esthesioneuroblastoma|9522/3
C0206717|T191|SY|0000021043|CHV|esthesioneuroblastoma olfactory|9522/3
C0206717|T191|SY|0000021043|CHV|esthesioneuroblastomas|9522/3
C0206717|T191|SY|0000021043|CHV|olfactory neuroblastoma|9522/3
C0206717|T191|PT|HP:0030068|HPO|Olfactory esthesioneuroblastoma|9522/3
C0206717|T191|PT|MTHU027102|ICPC2ICD10ENG|esthesioneuroblastoma|9522/3
C0206717|T191|PT|MTHU027104|ICPC2ICD10ENG|esthesioneuroepithelioma|9522/3
C0206717|T191|LLT|10001433|MDR|Aesthesioneuroblastoma|9522/3
C0206717|T191|PT|10001433|MDR|Aesthesioneuroblastoma|9522/3
C0206717|T191|LLT|10015498|MDR|Esthesioneuroblastoma|9522/3
C0206717|T191|LLT|10028732|MDR|Nasal cavity esthesioneuroblastoma|9522/3
C0206717|T191|LLT|10033863|MDR|Paranasal sinus esthesioneuroblastoma|9522/3
C0206717|T191|SY|351911|MEDCIN|malignant neoplasm neuroblastoma olfactory|9522/3
C0206717|T191|PT|351911|MEDCIN|Olfactory neuroblastoma|9522/3
C0206717|T191|ET|D018304|MSH|Aesthesioneuroblastoma|9522/3
C0206717|T191|PM|D018304|MSH|Aesthesioneuroblastomas|9522/3
C0206717|T191|ET|D018304|MSH|Esthesioneuroblastoma|9522/3
C0206717|T191|MH|D018304|MSH|Esthesioneuroblastoma, Olfactory|9522/3
C0206717|T191|PM|D018304|MSH|Esthesioneuroblastoma, Paranasal Sinus Nasal Cavity|9522/3
C0206717|T191|ET|D018304|MSH|Esthesioneuroblastoma, Paranasal Sinus-Nasal Cavity|9522/3
C0206717|T191|PM|D018304|MSH|Esthesioneuroblastomas|9522/3
C0206717|T191|PM|D018304|MSH|Esthesioneuroblastomas, Olfactory|9522/3
C0206717|T191|ET|D018304|MSH|Neuroblastoma, Olfactory|9522/3
C0206717|T191|PM|D018304|MSH|Neuroblastomas, Olfactory|9522/3
C0206717|T191|PM|D018304|MSH|Olfactory Esthesioneuroblastoma|9522/3
C0206717|T191|PM|D018304|MSH|Olfactory Esthesioneuroblastomas|9522/3
C0206717|T191|ET|D018304|MSH|Olfactory Neuroblastoma|9522/3
C0206717|T191|PM|D018304|MSH|Olfactory Neuroblastomas|9522/3
C0206717|T191|PM|D018304|MSH|Paranasal Sinus Nasal Cavity Esthesioneuroblastoma|9522/3
C0206717|T191|ET|D018304|MSH|Paranasal Sinus-Nasal Cavity Esthesioneuroblastoma|9522/3
C0206717|T191|PN|NOCODE|MTH|Olfactory Neuroblastoma|9522/3
C0206717|T191|SY|C6016|NCI|Accessory Sinus Esthesioneuroblastoma|9522/3
C0206717|T191|SY|C3789|NCI|Esthesioneuroblastoma|9522/3
C0206717|T191|SY|C6016|NCI|Esthesioneuroblastoma of Accessory Sinus|9522/3
C0206717|T191|SY|C6016|NCI|Esthesioneuroblastoma of Paranasal Sinus|9522/3
C0206717|T191|SY|C6016|NCI|Esthesioneuroblastoma of the Accessory Sinus|9522/3
C0206717|T191|SY|C6016|NCI|Esthesioneuroblastoma of the Paranasal Sinus|9522/3
C0206717|T191|SY|C3789|NCI|Esthesioneuroepithelioma|9522/3
C0206717|T191|SY|C3789|NCI|Olfactory Esthesioneuroblastoma|9522/3
C0206717|T191|PT|C3789|NCI|Olfactory Neuroblastoma|9522/3
C0206717|T191|SY|C3789|NCI|Olfactory Neuroepithelioma|9522/3
C0206717|T191|SY|C6016|NCI|Paranasal Sinus Esthesioneuroblastoma|9522/3
C0206717|T191|PT|C6016|NCI|Paranasal Sinus Olfactory Neuroblastoma|9522/3
C0206717|T191|DN|C3789|NCI_CTRP|Olfactory Neuroblastoma|9522/3
C0206717|T191|SY|CDR0000040691|PDQ|Esthesioneuroblastoma|9522/3
C0206717|T191|SY|CDR0000040691|PDQ|esthesioneuroblastoma, paranasal sinus and nasal cavity|9522/3
C0206717|T191|SY|CDR0000040691|PDQ|Esthesioneuroepithelioma|9522/3
C0206717|T191|SY|CDR0000040691|PDQ|nasal cavity and paranasal sinus esthesioneuroblastoma|9522/3
C0206717|T191|SY|CDR0000040691|PDQ|Olfactory Esthesioneuroblastoma|9522/3
C0206717|T191|SY|CDR0000040691|PDQ|Olfactory Neuroblastoma|9522/3
C0206717|T191|SY|CDR0000040691|PDQ|Olfactory Neuroepithelioma|9522/3
C0206717|T191|PT|CDR0000040691|PDQ|paranasal sinus and nasal cavity esthesioneuroblastoma|9522/3
C0206717|T191|OP|BBcD.|RCD|Aesthesioneuroepithelioma|9522/3
C0206717|T191|OP|BBcC.|RCD|Asthesioneuroblastoma|9522/3
C0206717|T191|PT|Xa99K|RCD|Olfactory neuroblastoma|9522/3
C0206717|T191|PT|Xa99L|RCD|Olfactory neuroepithelioma|9522/3
C0206717|T191|PTGB|76060004|SNOMEDCT_US|Aesthesioneuroblastoma|9522/3
C0206717|T191|SYGB|422886007|SNOMEDCT_US|Aesthesioneuroblastoma|9522/3
C0206717|T191|OAP|189938009|SNOMEDCT_US|Aesthesioneuroepithelioma|9522/3
C0206717|T191|PTGB|68614005|SNOMEDCT_US|Aesthesioneuroepithelioma|9522/3
C0206717|T191|OAP|189937004|SNOMEDCT_US|Asthesioneuroblastoma|9522/3
C0206717|T191|SY|76060004|SNOMEDCT_US|Asthesioneuroblastoma|9522/3
C0206717|T191|PT|76060004|SNOMEDCT_US|Esthesioneuroblastoma|9522/3
C0206717|T191|SY|422886007|SNOMEDCT_US|Esthesioneuroblastoma|9522/3
C0206717|T191|OAP|189938009|SNOMEDCT_US|Esthesioneuroepithelioma|9522/3
C0206717|T191|PT|68614005|SNOMEDCT_US|Esthesioneuroepithelioma|9522/3
C0206717|T191|PT|422886007|SNOMEDCT_US|Olfactory neuroblastoma|9522/3
C0206717|T191|SY|76060004|SNOMEDCT_US|Olfactory neuroblastoma|9522/3
C0206717|T191|SY|68614005|SNOMEDCT_US|Olfactory neuroepithelioma|9522/3
C0206717|T191|PT|0000021043|CHV|esthesioneuroblastoma|9523/3
C0206717|T191|SY|0000021043|CHV|esthesioneuroblastoma olfactory|9523/3
C0206717|T191|SY|0000021043|CHV|esthesioneuroblastomas|9523/3
C0206717|T191|SY|0000021043|CHV|olfactory neuroblastoma|9523/3
C0206717|T191|PT|HP:0030068|HPO|Olfactory esthesioneuroblastoma|9523/3
C0206717|T191|PT|MTHU027102|ICPC2ICD10ENG|esthesioneuroblastoma|9523/3
C0206717|T191|PT|MTHU027104|ICPC2ICD10ENG|esthesioneuroepithelioma|9523/3
C0206717|T191|PT|10001433|MDR|Aesthesioneuroblastoma|9523/3
C0206717|T191|LLT|10001433|MDR|Aesthesioneuroblastoma|9523/3
C0206717|T191|LLT|10015498|MDR|Esthesioneuroblastoma|9523/3
C0206717|T191|LLT|10028732|MDR|Nasal cavity esthesioneuroblastoma|9523/3
C0206717|T191|LLT|10033863|MDR|Paranasal sinus esthesioneuroblastoma|9523/3
C0206717|T191|SY|351911|MEDCIN|malignant neoplasm neuroblastoma olfactory|9523/3
C0206717|T191|PT|351911|MEDCIN|Olfactory neuroblastoma|9523/3
C0206717|T191|ET|D018304|MSH|Aesthesioneuroblastoma|9523/3
C0206717|T191|PM|D018304|MSH|Aesthesioneuroblastomas|9523/3
C0206717|T191|ET|D018304|MSH|Esthesioneuroblastoma|9523/3
C0206717|T191|MH|D018304|MSH|Esthesioneuroblastoma, Olfactory|9523/3
C0206717|T191|PM|D018304|MSH|Esthesioneuroblastoma, Paranasal Sinus Nasal Cavity|9523/3
C0206717|T191|ET|D018304|MSH|Esthesioneuroblastoma, Paranasal Sinus-Nasal Cavity|9523/3
C0206717|T191|PM|D018304|MSH|Esthesioneuroblastomas|9523/3
C0206717|T191|PM|D018304|MSH|Esthesioneuroblastomas, Olfactory|9523/3
C0206717|T191|ET|D018304|MSH|Neuroblastoma, Olfactory|9523/3
C0206717|T191|PM|D018304|MSH|Neuroblastomas, Olfactory|9523/3
C0206717|T191|PM|D018304|MSH|Olfactory Esthesioneuroblastoma|9523/3
C0206717|T191|PM|D018304|MSH|Olfactory Esthesioneuroblastomas|9523/3
C0206717|T191|ET|D018304|MSH|Olfactory Neuroblastoma|9523/3
C0206717|T191|PM|D018304|MSH|Olfactory Neuroblastomas|9523/3
C0206717|T191|PM|D018304|MSH|Paranasal Sinus Nasal Cavity Esthesioneuroblastoma|9523/3
C0206717|T191|ET|D018304|MSH|Paranasal Sinus-Nasal Cavity Esthesioneuroblastoma|9523/3
C0206717|T191|PN|NOCODE|MTH|Olfactory Neuroblastoma|9523/3
C0206717|T191|SY|C6016|NCI|Accessory Sinus Esthesioneuroblastoma|9523/3
C0206717|T191|SY|C3789|NCI|Esthesioneuroblastoma|9523/3
C0206717|T191|SY|C6016|NCI|Esthesioneuroblastoma of Accessory Sinus|9523/3
C0206717|T191|SY|C6016|NCI|Esthesioneuroblastoma of Paranasal Sinus|9523/3
C0206717|T191|SY|C6016|NCI|Esthesioneuroblastoma of the Accessory Sinus|9523/3
C0206717|T191|SY|C6016|NCI|Esthesioneuroblastoma of the Paranasal Sinus|9523/3
C0206717|T191|SY|C3789|NCI|Esthesioneuroepithelioma|9523/3
C0206717|T191|SY|C3789|NCI|Olfactory Esthesioneuroblastoma|9523/3
C0206717|T191|PT|C3789|NCI|Olfactory Neuroblastoma|9523/3
C0206717|T191|SY|C3789|NCI|Olfactory Neuroepithelioma|9523/3
C0206717|T191|SY|C6016|NCI|Paranasal Sinus Esthesioneuroblastoma|9523/3
C0206717|T191|PT|C6016|NCI|Paranasal Sinus Olfactory Neuroblastoma|9523/3
C0206717|T191|DN|C3789|NCI_CTRP|Olfactory Neuroblastoma|9523/3
C0206717|T191|SY|CDR0000040691|PDQ|Esthesioneuroblastoma|9523/3
C0206717|T191|SY|CDR0000040691|PDQ|esthesioneuroblastoma, paranasal sinus and nasal cavity|9523/3
C0206717|T191|SY|CDR0000040691|PDQ|Esthesioneuroepithelioma|9523/3
C0206717|T191|SY|CDR0000040691|PDQ|nasal cavity and paranasal sinus esthesioneuroblastoma|9523/3
C0206717|T191|SY|CDR0000040691|PDQ|Olfactory Esthesioneuroblastoma|9523/3
C0206717|T191|SY|CDR0000040691|PDQ|Olfactory Neuroblastoma|9523/3
C0206717|T191|SY|CDR0000040691|PDQ|Olfactory Neuroepithelioma|9523/3
C0206717|T191|PT|CDR0000040691|PDQ|paranasal sinus and nasal cavity esthesioneuroblastoma|9523/3
C0206717|T191|OP|BBcD.|RCD|Aesthesioneuroepithelioma|9523/3
C0206717|T191|OP|BBcC.|RCD|Asthesioneuroblastoma|9523/3
C0206717|T191|PT|Xa99K|RCD|Olfactory neuroblastoma|9523/3
C0206717|T191|PT|Xa99L|RCD|Olfactory neuroepithelioma|9523/3
C0206717|T191|PTGB|76060004|SNOMEDCT_US|Aesthesioneuroblastoma|9523/3
C0206717|T191|SYGB|422886007|SNOMEDCT_US|Aesthesioneuroblastoma|9523/3
C0206717|T191|OAP|189938009|SNOMEDCT_US|Aesthesioneuroepithelioma|9523/3
C0206717|T191|PTGB|68614005|SNOMEDCT_US|Aesthesioneuroepithelioma|9523/3
C0206717|T191|SY|76060004|SNOMEDCT_US|Asthesioneuroblastoma|9523/3
C0206717|T191|OAP|189937004|SNOMEDCT_US|Asthesioneuroblastoma|9523/3
C0206717|T191|SY|422886007|SNOMEDCT_US|Esthesioneuroblastoma|9523/3
C0206717|T191|PT|76060004|SNOMEDCT_US|Esthesioneuroblastoma|9523/3
C0206717|T191|OAP|189938009|SNOMEDCT_US|Esthesioneuroepithelioma|9523/3
C0206717|T191|PT|68614005|SNOMEDCT_US|Esthesioneuroepithelioma|9523/3
C0206717|T191|PT|422886007|SNOMEDCT_US|Olfactory neuroblastoma|9523/3
C0206717|T191|SY|76060004|SNOMEDCT_US|Olfactory neuroblastoma|9523/3
C0206717|T191|SY|68614005|SNOMEDCT_US|Olfactory neuroepithelioma|9523/3
C0025286|T191|ET|0000004656|AOD|meningioma|9530/0
C0025286|T191|SY|0000007930|CHV|brain meningioma tumors|9530/0
C0025286|T191|SY|0000007930|CHV|leptomeningioma|9530/0
C0025286|T191|SY|0000007930|CHV|lymphoplasmacyte-rich meningioma|9530/0
C0025286|T191|PT|0000007930|CHV|meningioma|9530/0
C0025286|T191|SY|0000007930|CHV|meningioma brain tumor|9530/0
C0025286|T191|SY|0000007930|CHV|meningiomas|9530/0
C0025286|T191|SY|0000007930|CHV|secretory meningioma|9530/0
C0025286|T191|PT|U000440|COSTAR|MENINGIOMA|9530/0
C0025286|T191|PT|2012-5515|CSP|meningioma|9530/0
C0025286|T191|SY|NOCODE|DXP|BRAIN TUMOR, MENINGIOMA|9530/0
C0025286|T191|SY|NOCODE|DXP|ENDOTHELIOMA, DURAL|9530/0
C0025286|T191|SY|NOCODE|DXP|FIBROBLASTOMA, ARACHNOIDAL|9530/0
C0025286|T191|SY|NOCODE|DXP|FIBROBLASTOMA, MENINGEAL|9530/0
C0025286|T191|SY|NOCODE|DXP|INTRACRANIAL NEOPLASM, MENINGIOMA|9530/0
C0025286|T191|SY|NOCODE|DXP|LEPTOMENINGIOMA|9530/0
C0025286|T191|DI|U001156|DXP|MENINGIOMA|9530/0
C0025286|T191|PT|HP:0002858|HPO|Meningioma|9530/0
C0348426|T191|HT|D32|ICD10|Benign neoplasm of meninges|9530/0
C0348426|T191|PX|D32.9|ICD10|Benign neoplasm of meninges, unspecified|9530/0
C0348426|T191|PS|D32.9|ICD10|Meninges, unspecified|9530/0
C0348426|T191|AB|D32|ICD10CM|Benign neoplasm of meninges|9530/0
C0348426|T191|HT|D32|ICD10CM|Benign neoplasm of meninges|9530/0
C0348426|T191|PT|D32.9|ICD10CM|Benign neoplasm of meninges, unspecified|9530/0
C0348426|T191|AB|D32.9|ICD10CM|Benign neoplasm of meninges, unspecified|9530/0
C0025286|T191|ET|D32.9|ICD10CM|Meningioma NOS|9530/0
C0348426|T191|PTN|N75005|ICPC2P|benign neoplasm of the meninges|9530/0
C0025286|T191|PTN|N75001|ICPC2P|meningioma|9530/0
C0025286|T191|PT|N75001|ICPC2P|Meningioma|9530/0
C0348426|T191|PT|N75005|ICPC2P|Neoplasm benign;meninges|9530/0
C0025286|T191|PT|U002900|LCH|Meningioma|9530/0
C0025286|T191|PT|sh85083561|LCH_NW|Meningioma|9530/0
C0025286|T191|PT|10027191|MDR|Meningioma|9530/0
C0025286|T191|LLT|10027191|MDR|Meningioma|9530/0
C0348426|T191|PT|272433|MEDCIN|benign neoplasm of meninges|9530/0
C0348426|T191|SY|272433|MEDCIN|benign tumor of meninges|9530/0
C0025286|T191|PT|31913|MEDCIN|meningioma|9530/0
C0025286|T191|ET|173|MEDLINEPLUS|Meningioma|9530/0
C0348426|T191|DEV|D008577|MSH|BENIGN MENINGEAL NEOPL|9530/0
C0348426|T191|PM|D008577|MSH|Benign Meningeal Neoplasm|9530/0
C0348426|T191|PEP|D008577|MSH|Benign Meningeal Neoplasms|9530/0
C0348426|T191|DEV|D008577|MSH|MENINGEAL NEOPL BENIGN|9530/0
C0348426|T191|PM|D008577|MSH|Meningeal Neoplasm, Benign|9530/0
C0348426|T191|ET|D008577|MSH|Meningeal Neoplasms, Benign|9530/0
C0025286|T191|MH|D008579|MSH|Meningioma|9530/0
C1384408|T191|PM|D008579|MSH|Meningioma, Microcystic|9530/0
C1384406|T191|PM|D008579|MSH|Meningioma, Secretory|9530/0
C0457190|T191|PM|D008579|MSH|Meningioma, Xanthomatous|9530/0
C0025286|T191|PM|D008579|MSH|Meningiomas|9530/0
C1384408|T191|PM|D008579|MSH|Meningiomas, Microcystic|9530/0
C1384406|T191|PM|D008579|MSH|Meningiomas, Secretory|9530/0
C0457190|T191|PM|D008579|MSH|Meningiomas, Xanthomatous|9530/0
C1384408|T191|PEP|D008579|MSH|Microcystic Meningioma|9530/0
C1384408|T191|PM|D008579|MSH|Microcystic Meningiomas|9530/0
C0348426|T191|PM|D008577|MSH|Neoplasm, Benign Meningeal|9530/0
C0348426|T191|PM|D008577|MSH|Neoplasms, Benign Meningeal|9530/0
C1384406|T191|PEP|D008579|MSH|Secretory Meningioma|9530/0
C1384406|T191|PM|D008579|MSH|Secretory Meningiomas|9530/0
C0457190|T191|PEP|D008579|MSH|Xanthomatous Meningioma|9530/0
C0457190|T191|PM|D008579|MSH|Xanthomatous Meningiomas|9530/0
C0348426|T191|PN|U001079|MTH|Benign neoplasm of meninges|9530/0
C0431119|T191|PN|NOCODE|MTH|Lymphoplasmacyte-rich meningioma|9530/0
C0025286|T191|PN|NOCODE|MTH|Meningioma|9530/0
C1762616|T191|PN|NOCODE|MTH|Meningioma, benign, no ICD-O subtype|9530/0
C1384408|T191|PN|NOCODE|MTH|Microcystic meningioma|9530/0
C1384406|T191|PN|NOCODE|MTH|Secretory meningioma|9530/0
C0348426|T191|ET|225.2|MTHICD9|Benign neoplasm of meninges NOS|9530/0
C0025286|T191|ET|225.2|MTHICD9|Meningioma|9530/0
C0348426|T191|SY|C4957|NCI|Benign Meningeal Neoplasm|9530/0
C0348426|T191|SY|C4957|NCI|Benign Meningeal Neoplasms|9530/0
C0348426|T191|SY|C4957|NCI|Benign Meningeal Tumor|9530/0
C0348426|T191|SY|C4957|NCI|Benign Meningeal Tumors|9530/0
C0348426|T191|SY|C4957|NCI|Benign Meninges Neoplasm|9530/0
C0348426|T191|SY|C4957|NCI|Benign Meninges Tumor|9530/0
C0348426|T191|SY|C4957|NCI|Benign Neoplasm of Meninges|9530/0
C0348426|T191|PT|C4957|NCI|Benign Neoplasm of the Meninges|9530/0
C0348426|T191|SY|C4957|NCI|Benign Neoplasms of Meninges|9530/0
C0348426|T191|SY|C4957|NCI|Benign Neoplasms of the Meninges|9530/0
C0348426|T191|SY|C4957|NCI|Benign Tumor of Meninges|9530/0
C0348426|T191|SY|C4957|NCI|Benign Tumor of the Meninges|9530/0
C0431119|T191|PT|C4720|NCI|Lymphoplasmacyte-Rich Meningioma|9530/0
C0348426|T191|SY|C4957|NCI|Meningeal Tumors, Benign|9530/0
C0025286|T191|SY|TCGA|NCI|Meningioma|9530/0
C0025286|T191|PT|C3230|NCI|Meningioma|9530/0
C1384408|T191|PT|C4721|NCI|Microcystic Meningioma|9530/0
C1384406|T191|PT|C4718|NCI|Secretory Meningioma|9530/0
C0348426|T191|PT|C4957|NCI_CPTAC|Benign Neoplasm of the Meninges|9530/0
C0025286|T191|PT|C3230|NCI_CPTAC|Meningioma|9530/0
C0025286|T191|PT|10027189|NCI_CTEP-SDC|Meningioma, NOS|9530/0
C0025286|T191|DN|C3230|NCI_CTRP|Meningioma|9530/0
C0025286|T191|PT|C3230|NCI_CTRP|Meningioma|9530/0
C0025286|T191|PT|CDR0000045783|NCI_NCI-GLOSS|meningioma|9530/0
C0025286|T191|PT|C3230|NCI_NICHD|Meningioma|9530/0
C0025286|T191|ET|CDR0000580900|PDQ|Meningioma|9530/0
C0025286|T191|PT|CDR0000580900|PDQ|meningioma|9530/0
C0025286|T191|PT|R0121679|QMR|MENINGIOMA|9530/0
C0348426|T191|PT|X78aZ|RCD|Benign tumour of meninges|9530/0
C0431119|T191|AB|X77pi|RCD|Lymphoplasmocyte-rich meningio|9530/0
C0431119|T191|PT|X77pi|RCD|Lymphoplasmocyte-rich meningioma|9530/0
C0025286|T191|PT|XM0C9|RCD|Meningioma|9530/0
C0025286|T191|SY|XM0C9|RCD|MGM - Meningioma|9530/0
C1384408|T191|PT|X77pj|RCD|Microcystic meningioma|9530/0
C1384406|T191|PT|X77pg|RCD|Secretory meningioma|9530/0
C0457190|T191|PT|Xa0aV|RCD|Xanthomatous meningioma|9530/0
C0348426|T191|PT|X78aZ|RCDAE|Benign tumor of meninges|9530/0
C0348426|T191|OA|ByuGP|RCDSY|Ben neop meninges, unspecif|9530/0
C0348426|T191|OP|ByuGP|RCDSY|Benign neoplasm of meninges, unspecified|9530/0
C0025286|T191|OP|BBdz.|RCDSY|Meningioma NOS|9530/0
C0025286|T191|OP|BBd..|RCDSY|Meningiomas|9530/0
C0348426|T191|PT|409659004|SNOMEDCT_US|Benign meningeal neoplasm|9530/0
C1762616|T191|PT|19453003|SNOMEDCT_US|Benign meningioma|9530/0
C0348426|T191|PT|109913001|SNOMEDCT_US|Benign neoplasm of meninges|9530/0
C0348426|T191|SY|109913001|SNOMEDCT_US|Benign tumor of meninges|9530/0
C0348426|T191|SYGB|109913001|SNOMEDCT_US|Benign tumour of meninges|9530/0
C0431119|T191|IS|19453003|SNOMEDCT_US|Lymphoplasmacyte-rich meningioma|9530/0
C0431119|T191|PT|253083007|SNOMEDCT_US|Lymphoplasmocyte-rich meningioma|9530/0
C0431119|T191|SY|19453003|SNOMEDCT_US|Lymphoplasmocyte-rich meningioma|9530/0
C0025286|T191|OAP|393566004|SNOMEDCT_US|Meningioma|9530/0
C0025286|T191|OAS|269643009|SNOMEDCT_US|Meningioma|9530/0
C0025286|T191|OAS|154621002|SNOMEDCT_US|Meningioma|9530/0
C0025286|T191|OF|393566004|SNOMEDCT_US|Meningioma|9530/0
C1762616|T191|OP|19453003|SNOMEDCT_US|Meningioma|9530/0
C1762616|T191|SY|19453003|SNOMEDCT_US|Meningioma, benign, no ICD-O subtype|9530/0
C1762616|T191|SY|19453003|SNOMEDCT_US|Meningioma, benign, no International Classification of Diseases for Oncology subtype|9530/0
C1762616|T191|IS|19453003|SNOMEDCT_US|Meningioma, NOS|9530/0
C1762616|T191|IS|19453003|SNOMEDCT_US|MGM - Meningioma|9530/0
C1384408|T191|SY|19453003|SNOMEDCT_US|Microcystic meningioma|9530/0
C1384408|T191|PT|253084001|SNOMEDCT_US|Microcystic meningioma|9530/0
C1384406|T191|PT|253081009|SNOMEDCT_US|Secretory meningioma|9530/0
C1384406|T191|SY|19453003|SNOMEDCT_US|Secretory meningioma|9530/0
C0457190|T191|PT|277999002|SNOMEDCT_US|Xanthomatous meningioma|9530/0
C0205834|T191|PT|0000020728|CHV|meningiomatosis|9530/1
C0205834|T191|SY|0000020728|CHV|multiple meningioma|9530/1
C0205834|T191|SY|0000020728|CHV|multiple meningiomas|9530/1
C0205834|T191|LLT|10065014|MDR|Multiple meningioma|9530/1
C0205834|T191|PM|D008579|MSH|Meningioma, Multiple|9530/1
C0205834|T191|PEP|D008579|MSH|Meningiomas, Multiple|9530/1
C0205834|T191|PM|D008579|MSH|Meningiomatoses|9530/1
C0205834|T191|ET|D008579|MSH|Meningiomatosis|9530/1
C0205834|T191|PM|D008579|MSH|Multiple Meningioma|9530/1
C0205834|T191|PM|D008579|MSH|Multiple Meningiomas|9530/1
C0205834|T191|SY|C3707|NCI|Meningiomas, Multiple|9530/1
C0205834|T191|PT|C3707|NCI|Meningiomatosis|9530/1
C0205834|T191|SY|Xa99N|RCD|Diffuse meningiomatosis|9530/1
C0205834|T191|PT|Xa99N|RCD|Meningiomatosis|9530/1
C0205834|T191|SY|Xa99N|RCD|Multiple meningiomas|9530/1
C0205834|T191|OP|BBd1.|RCDSY|Meningiomatosis NOS|9530/1
C0205834|T191|SY|40935003|SNOMEDCT_US|Diffuse meningiomatosis|9530/1
C0205834|T191|PT|40935003|SNOMEDCT_US|Meningiomatosis|9530/1
C0205834|T191|IS|40935003|SNOMEDCT_US|Meningiomatosis, NOS|9530/1
C0205834|T191|SY|40935003|SNOMEDCT_US|Multiple meningiomas|9530/1
C0259785|T191|PT|0000025234|CHV|malignant meningioma|9530/3
C0259785|T191|PT|U000397|COSTAR|MALIGNANT MENINGIOMA|9530/3
C0259785|T191|LLT|10073127|MDR|Anaplastic meningioma|9530/3
C0259785|T191|PT|10073127|MDR|Anaplastic meningioma|9530/3
C0259785|T191|LLT|10025672|MDR|Malignant meningioma|9530/3
C0259785|T191|LLT|10027193|MDR|Meningioma malignant|9530/3
C0259785|T191|PT|10027193|MDR|Meningioma malignant|9530/3
C0259785|T191|LLT|10027194|MDR|Meningioma malignant NOS|9530/3
C0259785|T191|HT|10027196|MDR|Meningiomas malignant|9530/3
C0259785|T191|PT|34998|MEDCIN|malignant meningioma|9530/3
C0259785|T191|PEP|D008579|MSH|Malignant Meningioma|9530/3
C0259785|T191|PM|D008579|MSH|Malignant Meningiomas|9530/3
C0259785|T191|PM|D008579|MSH|Meningioma, Malignant|9530/3
C0259785|T191|PM|D008579|MSH|Meningiomas, Malignant|9530/3
C0259785|T191|PN|NOCODE|MTH|Malignant Meningioma|9530/3
C0259785|T191|SY|C4051|NCI|Anaplastic Meningioma|9530/3
C0259785|T191|SY|C4051|NCI|Malignant Meningioma|9530/3
C0259785|T191|SY|C4051|NCI|Meningioma, Malignant|9530/3
C0259785|T191|PT|CDR0000045773|NCI_NCI-GLOSS|malignant meningioma|9530/3
C0259785|T191|SY|BBd2.|RCD|Anaplastic meningioma|9530/3
C0259785|T191|PT|BBd2.|RCD|Malignant meningioma|9530/3
C0259785|T191|OAS|134174002|SNOMEDCT_US|Anaplastic meningioma|9530/3
C0259785|T191|OAP|134174002|SNOMEDCT_US|Malignant meningioma|9530/3
C0259785|T191|SY|78303004|SNOMEDCT_US|Meningioma, anaplastic|9530/3
C0259785|T191|PT|78303004|SNOMEDCT_US|Meningioma, malignant|9530/3
C0334605|T191|PT|MTHU026177|ICPC2ICD10ENG|endotheliomatous; meningioma|9531/0
C0334605|T191|PT|MTHU048419|ICPC2ICD10ENG|meningioma; endotheliomatous|9531/0
C0334605|T191|PT|MTHU048426|ICPC2ICD10ENG|meningioma; meningotheliomatous|9531/0
C0334605|T191|PT|MTHU048429|ICPC2ICD10ENG|meningioma; syncytial|9531/0
C0334605|T191|PT|MTHU048749|ICPC2ICD10ENG|meningotheliomatous; meningioma|9531/0
C0334605|T191|PT|MTHU072532|ICPC2ICD10ENG|syncytial; meningioma|9531/0
C0334605|T191|PM|D008579|MSH|Meningioma, Meningotheliomatous|9531/0
C0334605|T191|PM|D008579|MSH|Meningiomas, Meningotheliomatous|9531/0
C0334605|T191|PEP|D008579|MSH|Meningotheliomatous Meningioma|9531/0
C0334605|T191|PM|D008579|MSH|Meningotheliomatous Meningiomas|9531/0
C0334605|T191|PN|NOCODE|MTH|Meningothelial meningioma|9531/0
C0334605|T191|PT|C4329|NCI|Meningothelial Meningioma|9531/0
C0334605|T191|SY|C4329|NCI|Meningotheliomatous Meningioma|9531/0
C0334605|T191|PT|BBd3.|RCD|Meningotheliomatous meningioma|9531/0
C0334605|T191|SY|BBd3.|RCD|Syncytial meningioma|9531/0
C0334605|T191|SY|68944005|SNOMEDCT_US|Endotheliomatous meningioma|9531/0
C0334605|T191|PT|68944005|SNOMEDCT_US|Meningothelial meningioma|9531/0
C0334605|T191|IS|68944005|SNOMEDCT_US|Meningotheliomatous meningioma|9531/0
C0334605|T191|SY|68944005|SNOMEDCT_US|Syncytial meningioma|9531/0
C0334606|T191|PT|MTHU028173|ICPC2ICD10ENG|fibroblastic; meningioma|9532/0
C0334606|T191|PT|MTHU028114|ICPC2ICD10ENG|fibrous; meningioma|9532/0
C0334606|T191|PT|MTHU048421|ICPC2ICD10ENG|meningioma; fibroblastic|9532/0
C0334606|T191|PT|MTHU048420|ICPC2ICD10ENG|meningioma; fibrous|9532/0
C0334606|T191|PEP|D008579|MSH|Fibrous Meningioma|9532/0
C0334606|T191|PM|D008579|MSH|Fibrous Meningiomas|9532/0
C0334606|T191|PM|D008579|MSH|Meningioma, Fibrous|9532/0
C0334606|T191|PM|D008579|MSH|Meningiomas, Fibrous|9532/0
C0334606|T191|SY|C4330|NCI|Fibroblastic Meningioma|9532/0
C0334606|T191|PT|C4330|NCI|Fibrous Meningioma|9532/0
C0334606|T191|SY|BBd4.|RCD|Fibroblastic meningioma|9532/0
C0334606|T191|PT|BBd4.|RCD|Fibrous meningioma|9532/0
C0334606|T191|SY|511008|SNOMEDCT_US|Fibroblastic meningioma|9532/0
C0334606|T191|PT|511008|SNOMEDCT_US|Fibrous meningioma|9532/0
C0334607|T191|SY|0000030013|CHV|meningioma psammomatous|9533/0
C0334607|T191|PT|0000030013|CHV|psammoma|9533/0
C0334607|T191|SY|0000030013|CHV|psammomas|9533/0
C0334607|T191|PT|MTHU048428|ICPC2ICD10ENG|meningioma; psammomatous|9533/0
C0334607|T191|PT|MTHU062229|ICPC2ICD10ENG|psammomatous; meningioma|9533/0
C0334607|T191|PM|D008579|MSH|Meningioma, Psammomatous|9533/0
C0334607|T191|PM|D008579|MSH|Meningiomas, Psammomatous|9533/0
C0334607|T191|PEP|D008579|MSH|Psammomatous Meningioma|9533/0
C0334607|T191|PM|D008579|MSH|Psammomatous Meningiomas|9533/0
C0334607|T191|PN|NOCODE|MTH|Psammomatous Meningioma|9533/0
C0334607|T191|PT|C4331|NCI|Psammomatous Meningioma|9533/0
C0334607|T191|PT|BBd5.|RCD|Psammomatous meningioma|9533/0
C0334607|T191|SY|38431002|SNOMEDCT_US|Psammoma|9533/0
C0334607|T191|PT|38431002|SNOMEDCT_US|Psammomatous meningioma|9533/0
C0334608|T191|PT|MTHU006371|ICPC2ICD10ENG|angiomatous; meningioma|9534/0
C0334608|T191|PT|MTHU048418|ICPC2ICD10ENG|meningioma; angiomatous|9534/0
C0334608|T191|PEP|D008579|MSH|Angiomatous Meningioma|9534/0
C0334608|T191|PM|D008579|MSH|Angiomatous Meningiomas|9534/0
C0334608|T191|PM|D008579|MSH|Meningioma, Angiomatous|9534/0
C0334608|T191|PM|D008579|MSH|Meningiomas, Angiomatous|9534/0
C0334608|T191|PN|NOCODE|MTH|Angiomatous Meningioma|9534/0
C0334608|T191|PT|C4332|NCI|Angiomatous Meningioma|9534/0
C0334608|T191|PT|BBd6.|RCD|Angiomatous meningioma|9534/0
C0334608|T191|PT|73918009|SNOMEDCT_US|Angiomatous meningioma|9534/0
C0334609|T191|PT|MTHU033754|ICPC2ICD10ENG|hemangioblastic; meningioma|9535/0
C0334609|T191|PT|MTHU048423|ICPC2ICD10ENG|meningioma; hemangioblastic|9535/0
C0334609|T191|PEP|D008579|MSH|Hemangioblastic Meningioma|9535/0
C0334609|T191|PM|D008579|MSH|Hemangioblastic Meningiomas|9535/0
C0334609|T191|PM|D008579|MSH|Meningioma, Hemangioblastic|9535/0
C0334609|T191|PM|D008579|MSH|Meningiomas, Hemangioblastic|9535/0
C0334609|T191|PN|NOCODE|MTH|Hemangioblastic Meningioma|9535/0
C0334609|T191|OP|C66817|NCI|Hemangioblastic Meningioma|9535/0
C0334609|T191|PT|C66817|NCI|Hemangioblastic Meningioma|9535/0
C0334609|T191|OP|BBd7.|RCD|Haemangioblastic meningioma|9535/0
C0334609|T191|OAP|189943002|SNOMEDCT_US|Haemangioblastic meningioma|9535/0
C0334609|T191|PTGB|35701008|SNOMEDCT_US|Haemangioblastic meningioma|9535/0
C0334609|T191|PT|35701008|SNOMEDCT_US|Hemangioblastic meningioma|9535/0
C0334609|T191|OAP|189943002|SNOMEDCT_US|Hemangioblastic meningioma|9535/0
C0334611|T191|PT|MTHU048422|ICPC2ICD10ENG|meningioma; mixed|9537/0
C0334611|T191|PT|MTHU048427|ICPC2ICD10ENG|meningioma; transitional|9537/0
C0334611|T191|PT|MTHU031216|ICPC2ICD10ENG|mixed; meningioma|9537/0
C0334611|T191|PT|MTHU056837|ICPC2ICD10ENG|transitional; meningioma|9537/0
C0334611|T191|PM|D008579|MSH|Meningioma, Transitional|9537/0
C0334611|T191|PM|D008579|MSH|Meningiomas, Transitional|9537/0
C0334611|T191|PEP|D008579|MSH|Transitional Meningioma|9537/0
C0334611|T191|PM|D008579|MSH|Transitional Meningiomas|9537/0
C0334611|T191|SY|C4333|NCI|Mixed Meningioma|9537/0
C0334611|T191|PT|C4333|NCI|Transitional Meningioma|9537/0
C0334611|T191|SY|BBd9.|RCD|Mixed meningioma|9537/0
C0334611|T191|PT|BBd9.|RCD|Transitional meningioma|9537/0
C0334611|T191|SY|64967004|SNOMEDCT_US|Mixed meningioma|9537/0
C0334611|T191|PT|64967004|SNOMEDCT_US|Transitional meningioma|9537/0
C0431121|T191|PEP|D008579|MSH|Clear Cell Meningioma|9538/1
C0431121|T191|PM|D008579|MSH|Clear Cell Meningiomas|9538/1
C0431121|T191|PM|D008579|MSH|Meningioma, Clear Cell|9538/1
C0431121|T191|PM|D008579|MSH|Meningiomas, Clear Cell|9538/1
C1370510|T191|PN|NOCODE|MTH|Chordoid meningioma|9538/1
C0431121|T191|PN|NOCODE|MTH|Clear Cell Meningioma|9538/1
C1370510|T191|PT|C6908|NCI|Chordoid Meningioma|9538/1
C1370510|T191|SY|TCGA|NCI|Chordoid Meningioma|9538/1
C0431121|T191|PT|C4722|NCI|Clear Cell Meningioma|9538/1
C0431121|T191|SY|TCGA|NCI|Clear Cell Meningioma|9538/1
C0431121|T191|PT|X77pk|RCD|Clear cell meningioma|9538/1
C1370510|T191|SY|399709001|SNOMEDCT_US|Chordoid meningioma|9538/1
C1370510|T191|IS|57606003|SNOMEDCT_US|Chordoid meningioma|9538/1
C0431121|T191|PT|57606003|SNOMEDCT_US|Clear cell meningioma|9538/1
C0431121|T191|OAP|134213009|SNOMEDCT_US|Clear cell meningioma|9538/1
C0431121|T191|OF|134213009|SNOMEDCT_US|Clear cell meningioma|9538/1
C1370510|T191|PT|399709001|SNOMEDCT_US|Meningioma, chordoid|9538/1
C0259786|T191|LLT|10069511|MDR|Rhabdoid meningioma|9538/3
C3163622|T191|PT|34997|MEDCIN|papillary meningioma|9538/3
C3163622|T191|PM|D008579|MSH|Meningioma, Papillary|9538/3
C3163622|T191|PM|D008579|MSH|Meningiomas, Papillary|9538/3
C3163622|T191|PEP|D008579|MSH|Papillary Meningioma|9538/3
C3163622|T191|PM|D008579|MSH|Papillary Meningiomas|9538/3
C3163622|T191|PN|NOCODE|MTH|Papillary Meningioma|9538/3
C0259786|T191|PN|NOCODE|MTH|Rhabdoid meningioma|9538/3
C3163622|T191|PT|C3904|NCI|Papillary Meningioma|9538/3
C3163622|T191|SY|TCGA|NCI|Papillary Meningioma|9538/3
C0259786|T191|PT|C6909|NCI|Rhabdoid Meningioma|9538/3
C0259786|T191|SY|TCGA|NCI|Rhabdoid Meningioma|9538/3
C3163622|T191|PT|BBdA.|RCD|Papillary meningioma|9538/3
C0259786|T191|PT|399469000|SNOMEDCT_US|Meningioma, rhabdoid|9538/3
C3163622|T191|IS|57606003|SNOMEDCT_US|Papillary meningioma|9538/3
C3163622|T191|PT|128840000|SNOMEDCT_US|Papillary meningioma|9538/3
C3163622|T191|SY|128840000|SNOMEDCT_US|Rhabdoid meningioma|9538/3
C0259786|T191|SY|399469000|SNOMEDCT_US|Rhabdoid meningioma|9538/3
C0431122|T191|PT|0000034149|CHV|atypical meningioma|9539/1
C0431122|T191|SY|0000034149|CHV|meningioma atypical|9539/1
C0431122|T191|PN|NOCODE|MTH|Atypical meningioma|9539/1
C0431122|T191|SY|TCGA|NCI|Atypical Meningioma|9539/1
C0431122|T191|PT|C4723|NCI|Atypical Meningioma|9539/1
C0431122|T191|PT|X77pl|RCD|Atypical meningioma|9539/1
C0431122|T191|PT|128914005|SNOMEDCT_US|Atypical meningioma|9539/1
C0334612|T191|PT|C4334|NCI|Meningeal Sarcomatosis|9539/3
C0334612|T191|SY|C4334|NCI|Meninges Sarcomatosis|9539/3
C0334612|T191|SY|C4334|NCI|Sarcomatosis of Meninges|9539/3
C0334612|T191|SY|C4334|NCI|Sarcomatosis of the Meninges|9539/3
C0334612|T191|PT|BBdB.|RCD|Meningeal sarcomatosis|9539/3
C0334612|T191|PT|14494009|SNOMEDCT_US|Meningeal sarcomatosis|9539/3
C0027830|T191|PT|0000008633|CHV|neurofibroma|9540/0
C0027830|T191|SY|0000008633|CHV|neurofibromas|9540/0
C0027830|T191|PT|2012-7305|CSP|neurofibroma|9540/0
C0027830|T191|PT|U003187|LCH|Neurofibroma|9540/0
C0027830|T191|PT|sh85091120|LCH_NW|Neurofibroma|9540/0
C0027830|T191|PT|10029267|MDR|Neurofibroma|9540/0
C0027830|T191|LLT|10029267|MDR|Neurofibroma|9540/0
C0027830|T191|MH|D009455|MSH|Neurofibroma|9540/0
C0027830|T191|PM|D009455|MSH|Neurofibromas|9540/0
C0027830|T191|PN|NOCODE|MTH|neurofibroma|9540/0
C1510961|T191|PT|C41426|NCI|Atypical Neurofibroma|9540/0
C0027830|T191|PT|C3272|NCI|Neurofibroma|9540/0
C0027830|T191|SY|TCGA|NCI|Neurofibroma|9540/0
C0027830|T191|PT|C3272|NCI_CDISC|NEUROFIBROMA, BENIGN|9540/0
C0027830|T191|PT|CDR0000045095|NCI_NCI-GLOSS|neurofibroma|9540/0
C0431123|T191|PT|X77pn|RCD|Circumscribed neurofibroma|9540/0
C0027830|T191|PT|Xa99R|RCD|Neurofibroma|9540/0
C0431123|T191|SY|X77pn|RCD|Solitary neurofibroma|9540/0
C0027830|T191|OP|BBe0.|RCDSY|Neurofibroma NOS|9540/0
C0027830|T191|SY|X77pm|RCDSY|Neurofibromas|9540/0
C1510961|T191|PT|734083001|SNOMEDCT_US|Atypical neurofibroma|9540/0
C0431123|T191|PT|253085000|SNOMEDCT_US|Circumscribed neurofibroma|9540/0
C0027830|T191|PT|89084002|SNOMEDCT_US|Neurofibroma|9540/0
C0027830|T191|PT|404029005|SNOMEDCT_US|Neurofibroma|9540/0
C0027830|T191|SY|89084002|SNOMEDCT_US|Neurofibroma, no ICD-O subtype|9540/0
C0027830|T191|SY|89084002|SNOMEDCT_US|Neurofibroma, no International Classification of Diseases for Oncology subtype|9540/0
C0027830|T191|IS|89084002|SNOMEDCT_US|Neurofibroma, NOS|9540/0
C0431123|T191|SY|253085000|SNOMEDCT_US|Solitary neurofibroma|9540/0
C0431123|T191|PT|404030000|SNOMEDCT_US|Solitary neurofibroma|9540/0
C0162678|T191|PT|1014171|CCPSS|NEUROFIBROMATOSIS|9540/1
C0162678|T191|SY|0000017943|CHV|multiple neurofibromatosis|9540/1
C0162678|T191|SY|0000017943|CHV|neurofibromatoses|9540/1
C0162678|T191|PT|0000017943|CHV|neurofibromatosis|9540/1
C0162678|T191|PT|U000475|COSTAR|NEUROFIBROMATOSIS|9540/1
C0162678|T191|ET|2012-7338|CSP|neurofibromatoses|9540/1
C0162678|T191|PT|2012-7338|CSP|neurofibromatosis|9540/1
C0162678|T191|SY|NOCODE|DXP|NEUROFIBROMA, MULTIPLE|9540/1
C0162678|T191|DI|U001284|DXP|NEUROFIBROMATOSIS|9540/1
C0162678|T191|ET|HP:0001067|HPO|multiple neurofibromas|9540/1
C0162678|T191|PT|HP:0001067|HPO|Neurofibromas|9540/1
C0162678|T191|SY|HP:0001067|HPO|Neurofibromata|9540/1
C0162678|T191|SY|HP:0001067|HPO|Neurofibromatosis|9540/1
C0162678|T191|PT|Q85.00|ICD10CM|Neurofibromatosis, unspecified|9540/1
C0162678|T191|AB|Q85.00|ICD10CM|Neurofibromatosis, unspecified|9540/1
C0162678|T191|HT|237.7|ICD9CM|Neurofibromatosis|9540/1
C0162678|T191|AB|237.70|ICD9CM|Neurofibromatosis NOS|9540/1
C0162678|T191|PT|237.70|ICD9CM|Neurofibromatosis, unspecified|9540/1
C0162678|T191|PT|MTHU052508|ICPC2ICD10ENG|neurofibromatosis|9540/1
C0162678|T191|PTN|A90012|ICPC2P|neurofibromatosis|9540/1
C0162678|T191|OP|N76001|ICPC2P|Neurofibromatosis|9540/1
C0162678|T191|PT|A90012|ICPC2P|Neurofibromatosis|9540/1
C0162678|T191|PT|U003188|LCH|Neurofibromatosis|9540/1
C0162678|T191|PT|sh85091121|LCH_NW|Neurofibromatosis|9540/1
C0162678|T191|PT|10029268|MDR|Neurofibromatosis|9540/1
C0162678|T191|LLT|10029268|MDR|Neurofibromatosis|9540/1
C0162678|T191|LLT|10029272|MDR|Neurofibromatosis, unspecified|9540/1
C0162678|T191|PT|99819|MEDCIN|neurofibromatosis|9540/1
C0162678|T191|PT|1387|MEDLINEPLUS|Neurofibromatosis|9540/1
C0162678|T191|PM|D017253|MSH|Multiple Neurofibroma|9540/1
C0162678|T191|ET|D017253|MSH|Multiple Neurofibromas|9540/1
C0162678|T191|PM|D017253|MSH|Neurofibroma, Multiple|9540/1
C0162678|T191|PM|D017253|MSH|Neurofibromas, Multiple|9540/1
C0162678|T191|MH|D017253|MSH|Neurofibromatoses|9540/1
C0162678|T191|ET|D017253|MSH|Neurofibromatosis|9540/1
C0162678|T191|ET|D017253|MSH|Neurofibromatosis Syndrome|9540/1
C0162678|T191|PM|D017253|MSH|Neurofibromatosis Syndromes|9540/1
C0162678|T191|PM|D017253|MSH|Syndrome, Neurofibromatosis|9540/1
C0162678|T191|PM|D017253|MSH|Syndromes, Neurofibromatosis|9540/1
C0162678|T191|PN|NOCODE|MTH|Neurofibromatoses|9540/1
C0162678|T191|PT|C6727|NCI|Neurofibromatosis|9540/1
C0162678|T191|PT|C6727|NCI_CPTAC|Neurofibromatosis|9540/1
C0162678|T191|PT|10029268|NCI_CTEP-SDC|Neurofibromatosis|9540/1
C0162678|T191|PT|C6727|NCI_NICHD|Neurofibromatosis|9540/1
C0162678|T191|SY|C6727|NCI_NICHD|Neurofibromatosis Syndrome|9540/1
C0162678|T191|PT|Xa99T|RCD|Neurofibromatosis|9540/1
C0162678|T191|SY|Xa99T|RCD|NF - Neurofibromatosis|9540/1
C0162678|T191|IS|BBe1.|RCDSY|Multiple neurofibromatosis|9540/1
C0162678|T191|OP|BBe1.|RCDSY|Neurofibromatosis NOS|9540/1
C0162678|T191|SY|19133005|SNOMEDCT_US|Clinical neurofibromatosis|9540/1
C0162678|T191|SY|81669005|SNOMEDCT_US|Multiple neurofibromatosis|9540/1
C0162678|T191|OAP|154642000|SNOMEDCT_US|Neurofibromatosis|9540/1
C0162678|T191|OF|154642000|SNOMEDCT_US|Neurofibromatosis|9540/1
C0162678|T191|PT|81669005|SNOMEDCT_US|Neurofibromatosis|9540/1
C0162678|T191|PT|19133005|SNOMEDCT_US|Neurofibromatosis syndrome|9540/1
C0162678|T191|IS|81669005|SNOMEDCT_US|Neurofibromatosis, NOS|9540/1
C0162678|T191|SY|19133005|SNOMEDCT_US|NF - Neurofibromatosis|9540/1
C0474847|T191|PT|0000037072|CHV|malignant melanotic schwannoma|9540/3
C0751690|T191|PT|0000048479|CHV|malignant schwannoma|9540/3
C0751690|T191|PT|0000045030|CHV|malignant schwannoma|9540/3
C0751690|T191|SY|0000048479|CHV|mpnst|9540/3
C0751690|T191|SY|HP:0100697|HPO|Malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|SY|HP:0100697|HPO|Malignant schwannoma|9540/3
C0751690|T191|LLT|10026667|MDR|Malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|LLT|10073836|MDR|Malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|LLT|10029236|MDR|Neurilemmoma malignant|9540/3
C0751690|T191|LLT|10029239|MDR|Neurilemoma malignant|9540/3
C0751690|T191|LLT|10034589|MDR|Peripheral nerve sheath tumor malignant|9540/3
C0751690|T191|LLT|10034590|MDR|Peripheral nerve sheath tumour malignant|9540/3
C0751690|T191|LLT|10058387|MDR|Schwannoma malignant|9540/3
C0474847|T191|PT|355154|MEDCIN|malignant melanotic nerve sheath tumor|9540/3
C0751690|T191|PT|271574|MEDCIN|malignant neurilemoma|9540/3
C1266188|T191|PT|271573|MEDCIN|malignant perineurioma|9540/3
C0751690|T191|SY|271571|MEDCIN|malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|SY|271571|MEDCIN|MPNST|9540/3
C0751690|T191|ET|D018319|MSH|Malignant Neurilemmoma|9540/3
C0751690|T191|PM|D018319|MSH|Malignant Neurilemmomas|9540/3
C0751690|T191|ET|D018319|MSH|Malignant Neurilemoma|9540/3
C0751690|T191|PM|D018319|MSH|Malignant Neurilemomas|9540/3
C0751690|T191|ET|D018319|MSH|Malignant Peripheral Nerve Sheath Tumor|9540/3
C0751690|T191|PEP|D018319|MSH|Malignant Peripheral Nerve Sheath Tumors|9540/3
C0751690|T191|PM|D018319|MSH|Malignant Schwannoma|9540/3
C0751690|T191|PM|D018319|MSH|Malignant Schwannomas|9540/3
C0751690|T191|ET|D018319|MSH|MPNST|9540/3
C0751690|T191|PM|D018319|MSH|Neurilemmoma, Malignant|9540/3
C0751690|T191|ET|D018319|MSH|Neurilemmosarcoma|9540/3
C0751690|T191|PM|D018319|MSH|Neurilemmosarcomas|9540/3
C0751690|T191|PM|D018319|MSH|Neurilemoma, Malignant|9540/3
C0751690|T191|ET|D018319|MSH|Peripheral Nerve Sheath Tumors, Malignant|9540/3
C0751690|T191|ET|D018319|MSH|Schwannoma, Malignant|9540/3
C0751690|T191|PN|NOCODE|MTH|Malignant Peripheral Nerve Sheath Tumor|9540/3
C1333821|T191|PT|C6560|NCI|Glandular Malignant Peripheral Nerve Sheath Tumor|9540/3
C1333821|T191|SY|C6560|NCI|Glandular MPNST|9540/3
C1333821|T191|SY|C6560|NCI|Malignant Glandular Neoplasm of Peripheral Nerve Sheath|9540/3
C1333821|T191|SY|C6560|NCI|Malignant Glandular Neoplasm of the Peripheral Nerve Sheath|9540/3
C1333821|T191|SY|C6560|NCI|Malignant Glandular Peripheral Nerve Sheath Neoplasm|9540/3
C1333821|T191|SY|C6560|NCI|Malignant Glandular Peripheral Nerve Sheath Tumor|9540/3
C1333821|T191|SY|C6560|NCI|Malignant Glandular Schwannoma|9540/3
C1333821|T191|SY|C6560|NCI|Malignant Glandular Tumor of Peripheral Nerve Sheath|9540/3
C1333821|T191|SY|C6560|NCI|Malignant Glandular Tumor of the Peripheral Nerve Sheath|9540/3
C0474847|T191|SY|C4748|NCI|Malignant Melanocytic Neoplasm of Peripheral Nerve Sheath|9540/3
C0474847|T191|SY|C4748|NCI|Malignant Melanocytic Neoplasm of the Peripheral Nerve Sheath|9540/3
C0474847|T191|SY|C4748|NCI|Malignant Melanocytic Peripheral Nerve Sheath Tumor|9540/3
C0474847|T191|PT|C4748|NCI|Malignant Melanotic Peripheral Nerve Sheath Tumor|9540/3
C0474847|T191|SY|TCGA|NCI|Malignant Melanotic Peripheral Nerve Sheath Tumor|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Neoplasm of Peripheral Nerve Sheath|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Neoplasm of the Peripheral Nerve Sheath|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Neurilemmoma|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Neurilemoma|9540/3
C1266188|T191|SY|C66845|NCI|Malignant Perineurioma|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Peripheral Nerve Sheath Neoplasm|9540/3
C0751690|T191|PT|C3798|NCI|Malignant Peripheral Nerve Sheath Tumor|9540/3
C0751690|T191|SY|TCGA|NCI|Malignant Peripheral Nerve Sheath Tumor|9540/3
C1266188|T191|PT|C66845|NCI|Malignant Peripheral Nerve Sheath Tumor with Perineurial Differentiation|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Peripheral Nerve Sheath Tumour|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Schwannoma|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Tumor of Peripheral Nerve Sheath|9540/3
C0751690|T191|SY|C3798|NCI|Malignant Tumor of the Peripheral Nerve Sheath|9540/3
C0474847|T191|SY|C4748|NCI|Melanocytic MPNST|9540/3
C0751690|T191|AB|C3798|NCI|MPNST|9540/3
C0751690|T191|SY|C3798|NCI|Neurofibrosarcoma|9540/3
C0751690|T191|SY|C3798|NCI|Neurogenic Sarcoma|9540/3
C1266188|T191|SY|C66845|NCI|Perineurial Malignant Peripheral Nerve Sheath Tumor|9540/3
C0751690|T191|SY|C3798|NCI_CDISC|Malignant Neurilemmoma|9540/3
C0751690|T191|SY|C3798|NCI_CDISC|Malignant Peripheral Nerve Sheath Tumour|9540/3
C0751690|T191|SY|C3798|NCI_CDISC|Neurofibrosarcoma, Malignant|9540/3
C0751690|T191|PT|C3798|NCI_CDISC|SCHWANNOMA, MALIGNANT|9540/3
C0751690|T191|PT|C3798|NCI_CPTAC|Malignant Peripheral Nerve Sheath Tumor|9540/3
C0751690|T191|SY|10026667|NCI_CTEP-SDC|Malig. periph. nerve sheath tum.|9540/3
C0751690|T191|PT|10026667|NCI_CTEP-SDC|Malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|PT|CDR0000335496|NCI_NCI-GLOSS|malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|PT|CDR0000335498|NCI_NCI-GLOSS|MPNST|9540/3
C0431127|T191|OA|X77pv|RCD|Mal Schwann+mesench+epith diff|9540/3
C0751690|T191|AB|Xa99V|RCD|Malig periph nerve sheath tum|9540/3
C0431127|T191|OA|X77pv|RCD|Malig Schwan+div mesench diff|9540/3
C0431127|T191|OA|X77pv|RCD|Malig Schwann+div epithel diff|9540/3
C0431127|T191|OA|X77pv|RCD|Malig Schwannoma + divergent mesenchymal & epithelial diff|9540/3
C0431127|T191|OA|X77pv|RCD|Malig Schwannoma with divergent epithelial differentiation|9540/3
C0431127|T191|OA|X77pv|RCD|Malig Schwannoma with divergent mesenchymal differentiation|9540/3
C0474847|T191|SY|X77py|RCD|Malignant melanotic Schwannoma|9540/3
C0751690|T191|OP|BBe7.|RCD|Malignant neurilemmoma|9540/3
C0751690|T191|PT|Xa99V|RCD|Malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|SY|Xa99V|RCD|Malignant Schwannoma|9540/3
C0431127|T191|IS|X77pv|RCD|Malignant Schwannoma with divergent epithelial differentiation|9540/3
C0431127|T191|OP|X77pv|RCD|Malignant Schwannoma with divergent mesenchymal and epithelial differentiation|9540/3
C0431127|T191|IS|X77pv|RCD|Malignant Schwannoma with divergent mesenchymal differentiation|9540/3
C0474847|T191|AB|X77py|RCD|Melan mal perip nerv sheat tum|9540/3
C0474847|T191|PT|X77py|RCD|Melanotic malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|SY|Xa99V|RCD|MPNST - Malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|AB|Xa99V|RCD|MPNST-Mal perip ner sheath tum|9540/3
C0751690|T191|SY|Xa99V|RCD|Neurilemmosarcoma|9540/3
C0751690|T191|OP|BBe7.|RCDAE|Malignant neurilemoma|9540/3
C0751690|T191|PT|Xa99V|RCDAE|Malignant peripheral nerve sheath tumor|9540/3
C0474847|T191|PT|X77py|RCDAE|Melanotic malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|SY|Xa99V|RCDAE|MPNST - Malignant peripheral nerve sheath tumor|9540/3
C1333821|T191|PT|699659007|SNOMEDCT_US|Glandular malignant peripheral nerve sheath tumor|9540/3
C1333821|T191|PT|699658004|SNOMEDCT_US|Glandular malignant peripheral nerve sheath tumor|9540/3
C1333821|T191|PTGB|699659007|SNOMEDCT_US|Glandular malignant peripheral nerve sheath tumour|9540/3
C1333821|T191|PTGB|699658004|SNOMEDCT_US|Glandular malignant peripheral nerve sheath tumour|9540/3
C0474847|T191|SY|253094006|SNOMEDCT_US|Malignant melanotic neurilemmoma|9540/3
C0474847|T191|SY|404039004|SNOMEDCT_US|Malignant melanotic neurilemmoma|9540/3
C0474847|T191|IS|253094006|SNOMEDCT_US|Malignant melanotic Schwannoma|9540/3
C0474847|T191|SY|253094006|SNOMEDCT_US|Malignant melanotic schwannoma|9540/3
C0474847|T191|SY|404039004|SNOMEDCT_US|Malignant melanotic schwannoma|9540/3
C0751690|T191|SYGB|404037002|SNOMEDCT_US|Malignant neurilemmoma|9540/3
C0751690|T191|OAP|189949003|SNOMEDCT_US|Malignant neurilemmoma|9540/3
C0751690|T191|OF|189949003|SNOMEDCT_US|Malignant neurilemmoma|9540/3
C0431127|T191|SY|253092005|SNOMEDCT_US|Malignant neurilemmoma with divergent mesenchymal and epithelial differentiation|9540/3
C0751690|T191|SY|404037002|SNOMEDCT_US|Malignant neurilemoma|9540/3
C1266188|T191|PT|761958009|SNOMEDCT_US|Malignant perineurioma|9540/3
C1266188|T191|OAP|734069003|SNOMEDCT_US|Malignant peripheral nerve sheath neoplasm with perineurial differentiation|9540/3
C1266188|T191|SY|761958009|SNOMEDCT_US|Malignant peripheral nerve sheath neoplasm with perineurial differentiation|9540/3
C1266188|T191|SY|128796000|SNOMEDCT_US|Malignant peripheral nerve sheath neoplasm with perineurial differentiation|9540/3
C0751690|T191|PT|404037002|SNOMEDCT_US|Malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|PT|19897006|SNOMEDCT_US|Malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|OAP|134324009|SNOMEDCT_US|Malignant peripheral nerve sheath tumor|9540/3
C0431127|T191|PT|253092005|SNOMEDCT_US|Malignant peripheral nerve sheath tumor with divergent mesenchymal and epithelial differentiation|9540/3
C1266188|T191|SY|761958009|SNOMEDCT_US|Malignant peripheral nerve sheath tumor with perineurial differentiation|9540/3
C0751690|T191|OAP|134324009|SNOMEDCT_US|Malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|PTGB|404037002|SNOMEDCT_US|Malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|PTGB|19897006|SNOMEDCT_US|Malignant peripheral nerve sheath tumour|9540/3
C0431127|T191|PTGB|253092005|SNOMEDCT_US|Malignant peripheral nerve sheath tumour with divergent mesenchymal and epithelial differentiation|9540/3
C1266188|T191|SYGB|761958009|SNOMEDCT_US|Malignant peripheral nerve sheath tumour with perineurial differentiation|9540/3
C0751690|T191|OAS|77418004|SNOMEDCT_US|Malignant Schwannoma|9540/3
C0751690|T191|SY|404037002|SNOMEDCT_US|Malignant schwannoma|9540/3
C0431127|T191|IS|253092005|SNOMEDCT_US|Malignant Schwannoma with divergent epithelial differentiation|9540/3
C0431127|T191|SY|253092005|SNOMEDCT_US|Malignant schwannoma with divergent epithelial differentiation|9540/3
C0431127|T191|SY|253092005|SNOMEDCT_US|Malignant schwannoma with divergent mesenchymal and epithelial differentiation|9540/3
C0431127|T191|OP|253092005|SNOMEDCT_US|Malignant Schwannoma with divergent mesenchymal and epithelial differentiation|9540/3
C0431127|T191|IS|253092005|SNOMEDCT_US|Malignant Schwannoma with divergent mesenchymal differentiation|9540/3
C0431127|T191|SY|253092005|SNOMEDCT_US|Malignant schwannoma with divergent mesenchymal differentiation|9540/3
C0751690|T191|IS|77418004|SNOMEDCT_US|Malignant Schwannoma, NOS|9540/3
C0474847|T191|PT|404039004|SNOMEDCT_US|Melanotic malignant nerve sheath tumor|9540/3
C0474847|T191|PTGB|404039004|SNOMEDCT_US|Melanotic malignant nerve sheath tumour|9540/3
C0474847|T191|OAP|253095007|SNOMEDCT_US|Melanotic malignant peripheral nerve sheath tumor|9540/3
C0474847|T191|PT|253094006|SNOMEDCT_US|Melanotic malignant peripheral nerve sheath tumor|9540/3
C0474847|T191|OAP|253095007|SNOMEDCT_US|Melanotic malignant peripheral nerve sheath tumour|9540/3
C0474847|T191|OF|253095007|SNOMEDCT_US|Melanotic malignant peripheral nerve sheath tumour|9540/3
C0474847|T191|PTGB|253094006|SNOMEDCT_US|Melanotic malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|IS|19897006|SNOMEDCT_US|MPNST|9540/3
C0751690|T191|OAS|134324009|SNOMEDCT_US|MPNST - Malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|SY|19897006|SNOMEDCT_US|MPNST - Malignant peripheral nerve sheath tumor|9540/3
C0751690|T191|OAS|134324009|SNOMEDCT_US|MPNST - Malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|SYGB|19897006|SNOMEDCT_US|MPNST - Malignant peripheral nerve sheath tumour|9540/3
C0751690|T191|OAS|77418004|SNOMEDCT_US|Neurilemmoma, malignant|9540/3
C0751690|T191|OAS|77418004|SNOMEDCT_US|Neurilemmosarcoma|9540/3
C0751690|T191|OAP|77418004|SNOMEDCT_US|Neurilemoma, malignant|9540/3
C1266188|T191|IS|128796000|SNOMEDCT_US|Perineural MPNST|9540/3
C1266188|T191|PT|128796000|SNOMEDCT_US|Perineurioma, malignant|9540/3
C0334613|T191|PT|C66841|NCI|Melanotic Neurofibroma|9541/0
C0334613|T191|SY|C66841|NCI|Pigmented Neurofibroma|9541/0
C0334613|T191|PT|BBe3.|RCD|Melanotic neurofibroma|9541/0
C0334613|T191|PT|28237007|SNOMEDCT_US|Melanotic neurofibroma|9541/0
C0334613|T191|PT|703088001|SNOMEDCT_US|Pigmented neurofibroma|9541/0
C1321427|T191|PT|355153|MEDCIN|malignant epithelioid nerve sheath tumor|9542/3
C1321427|T191|SY|355153|MEDCIN|malignant peripheral nerve sheath tumor epithelioid|9542/3
C1321427|T191|PN|NOCODE|MTH|Epithelioid Malignant Peripheral Nerve Sheath Tumor|9542/3
C1321427|T191|PT|C6561|NCI|Epithelioid Malignant Peripheral Nerve Sheath Tumor|9542/3
C1321427|T191|SY|TCGA|NCI|Epithelioid Malignant Peripheral Nerve Sheath Tumor|9542/3
C1321427|T191|SY|C6561|NCI|Epithelioid MPNST|9542/3
C1321427|T191|SY|C6561|NCI|Malignant Epithelioid Neoplasm of Peripheral Nerve Sheath|9542/3
C1321427|T191|SY|C6561|NCI|Malignant Epithelioid Neoplasm of the Peripheral Nerve Sheath|9542/3
C1321427|T191|SY|C6561|NCI|Malignant Epithelioid Peripheral Nerve Sheath Neoplasm|9542/3
C1321427|T191|SY|C6561|NCI|Malignant Epithelioid Peripheral Nerve Sheath Tumor|9542/3
C1321427|T191|SY|C6561|NCI|Malignant Epithelioid Tumor of Peripheral Nerve Sheath|9542/3
C1321427|T191|SY|C6561|NCI|Malignant Epithelioid Tumor of the Peripheral Nerve Sheath|9542/3
C1321427|T191|AB|X77px|RCD|Epithelioid malig nerve sh tum|9542/3
C1321427|T191|PT|X77px|RCD|Epithelioid malignant nerve sheath tumour|9542/3
C1321427|T191|PT|X77px|RCDAE|Epithelioid malignant nerve sheath tumor|9542/3
C1321427|T191|PT|404038007|SNOMEDCT_US|Epithelioid malignant nerve sheath tumor|9542/3
C1321427|T191|PT|253093000|SNOMEDCT_US|Epithelioid malignant nerve sheath tumor|9542/3
C1321427|T191|PTGB|253093000|SNOMEDCT_US|Epithelioid malignant nerve sheath tumour|9542/3
C1321427|T191|PTGB|404038007|SNOMEDCT_US|Epithelioid malignant nerve sheath tumour|9542/3
C1321427|T191|IS|19897006|SNOMEDCT_US|Epithelioid MPNST|9542/3
C1321427|T191|SY|253093000|SNOMEDCT_US|Epithelioid MPNST|9542/3
C1321427|T191|SY|253093000|SNOMEDCT_US|Malignant peripheral nerve sheath tumor, epithelioid|9542/3
C1321427|T191|SYGB|253093000|SNOMEDCT_US|Malignant peripheral nerve sheath tumour, epithelioid|9542/3
C0206728|T191|SY|0000021052|CHV|neurofibroma plexiform|9550/0
C0206728|T191|PT|0000021052|CHV|plexiform neurofibroma|9550/0
C0206728|T191|SY|0000021052|CHV|plexiform neuromas|9550/0
C0206728|T191|PT|HP:0009732|HPO|Plexiform neurofibroma|9550/0
C0206728|T191|PT|MTHU057010|ICPC2ICD10ENG|pachydermatocele|9550/0
C0206728|T191|LLT|10065866|MDR|Plexiform neurofibroma|9550/0
C0206728|T191|PM|D018318|MSH|Elephantiasis Neuromatoses|9550/0
C0206728|T191|ET|D018318|MSH|Elephantiasis Neuromatosis|9550/0
C0206728|T191|MH|D018318|MSH|Neurofibroma, Plexiform|9550/0
C0206728|T191|PM|D018318|MSH|Neurofibromas, Plexiform|9550/0
C0206728|T191|PM|D018318|MSH|Neuroma, Plexiform|9550/0
C0206728|T191|ET|D018318|MSH|Neuromas, Plexiform|9550/0
C0206728|T191|ET|D018318|MSH|Pachydermatocele|9550/0
C0206728|T191|PM|D018318|MSH|Pachydermatoceles|9550/0
C0206728|T191|PM|D018318|MSH|Plexiform Neurofibroma|9550/0
C0206728|T191|PM|D018318|MSH|Plexiform Neurofibromas|9550/0
C0206728|T191|PM|D018318|MSH|Plexiform Neuroma|9550/0
C0206728|T191|PM|D018318|MSH|Plexiform Neuromas|9550/0
C0206728|T191|ET|D018318|MSH|Tumor Royale|9550/0
C0206728|T191|PN|NOCODE|MTH|Plexiform Neurofibroma|9550/0
C0206728|T191|PT|C3797|NCI|Plexiform Neurofibroma|9550/0
C0206728|T191|SY|TCGA|NCI|Plexiform Neurofibroma|9550/0
C0206728|T191|PT|10065866|NCI_CTEP-SDC|Plexiform neurofibroma|9550/0
C0206728|T191|DN|C3797|NCI_CTRP|Plexiform Neurofibroma|9550/0
C0206728|T191|PT|CDR0000045094|NCI_NCI-GLOSS|plexiform neurofibroma|9550/0
C0206728|T191|PT|CDR0000472003|PDQ|plexiform neurofibroma|9550/0
C0206728|T191|PT|BBe4.|RCD|Plexiform neurofibroma|9550/0
C0206728|T191|SY|BBe4.|RCD|Plexiform neuroma|9550/0
C0206728|T191|PT|41252002|SNOMEDCT_US|Plexiform neurofibroma|9550/0
C0206728|T191|PT|403818001|SNOMEDCT_US|Plexiform neurofibroma|9550/0
C0206728|T191|SY|41252002|SNOMEDCT_US|Plexiform neuroma|9550/0
C0027809|T191|PT|0020072|CCPSS|SCHWANNOMA|9560/0
C0027809|T191|SY|0000008624|CHV|ancient schwannoma|9560/0
C0027809|T191|PT|0000008624|CHV|neurilemmoma|9560/0
C0027809|T191|SY|0000008624|CHV|neurilemmomas|9560/0
C0027809|T191|SY|0000008624|CHV|neurilemoma|9560/0
C0027809|T191|SY|0000008624|CHV|neurinoma|9560/0
C0027809|T191|SY|0000008624|CHV|neurinomas|9560/0
C0027809|T191|SY|0000008624|CHV|schwannoma|9560/0
C0027809|T191|SY|0000008624|CHV|schwannomas|9560/0
C0027809|T191|ET|2012-6947|CSP|neurilemmoma|9560/0
C0027809|T191|ET|2012-6947|CSP|neurinoma|9560/0
C0027809|T191|ET|2012-6947|CSP|schwannoma|9560/0
C0027809|T191|SY|HP:0100008|HPO|Neurilemmoma|9560/0
C0027809|T191|SY|HP:0100008|HPO|Neurinoma|9560/0
C0027809|T191|SY|HP:0100008|HPO|Neurolemmoma|9560/0
C0027809|T191|SY|HP:0100008|HPO|Schwann cell tumor|9560/0
C0027809|T191|SY|HP:0100008|HPO|Schwann cell tumour|9560/0
C0027809|T191|PT|HP:0100008|HPO|Schwannoma|9560/0
C0027809|T191|ET|HP:0100008|HPO|Schwannomas|9560/0
C0027809|T191|LA|LA26519-1|LNC|Schwannoma, NOS|9560/0
C0027809|T191|LLT|10029234|MDR|Neurilemmoma|9560/0
C0027809|T191|LLT|10029237|MDR|Neurilemoma|9560/0
C0027809|T191|LLT|10039667|MDR|Schwannoma|9560/0
C0027809|T191|PT|10039667|MDR|Schwannoma|9560/0
C0027809|T191|MH|D009442|MSH|Neurilemmoma|9560/0
C0027809|T191|PM|D009442|MSH|Neurilemmomas|9560/0
C0027809|T191|ET|D009442|MSH|Neurilemoma|9560/0
C0027809|T191|PM|D009442|MSH|Neurilemomas|9560/0
C0027809|T191|ET|D009442|MSH|Neurinoma|9560/0
C0027809|T191|PM|D009442|MSH|Neurinomas|9560/0
C0027809|T191|ET|D009442|MSH|Schwannoma|9560/0
C0027809|T191|PM|D009442|MSH|Schwannomas|9560/0
C0431124|T191|PN|NOCODE|MTH|Cellular Schwannoma|9560/0
C1536561|T191|PN|NOCODE|MTH|Degenerated Schwannoma|9560/0
C0027809|T191|PN|NOCODE|MTH|Neurilemmoma|9560/0
C1370659|T191|PN|NOCODE|MTH|Plexiform Schwannoma|9560/0
C1536561|T191|SY|C6556|NCI|Ancient Neurilemmoma|9560/0
C1536561|T191|SY|C6556|NCI|Ancient Schwannoma|9560/0
C0027809|T191|SY|C3269|NCI|Benign Neurilemmoma|9560/0
C0027809|T191|SY|C3269|NCI|Benign Schwannoma|9560/0
C0431124|T191|SY|C4724|NCI|Cellular Neurilemmoma|9560/0
C0431124|T191|SY|C4724|NCI|Cellular Neurinoma|9560/0
C0431124|T191|PT|C4724|NCI|Cellular Schwannoma|9560/0
C0431124|T191|SY|TCGA|NCI|Cellular Schwannoma|9560/0
C1536561|T191|SY|C6556|NCI|Degenerated Neurilemmoma|9560/0
C1536561|T191|PT|C6556|NCI|Degenerated Schwannoma|9560/0
C0027809|T191|SY|C3269|NCI|Neurilemmoma|9560/0
C0027809|T191|OP|C3269|NCI|Neurinoma|9560/0
C1370659|T191|SY|C6969|NCI|Plexiform Neurilemmoma|9560/0
C1370659|T191|SY|C6969|NCI|Plexiform Neurinoma|9560/0
C1370659|T191|SY|TCGA|NCI|Plexiform Schwannoma|9560/0
C1370659|T191|PT|C6969|NCI|Plexiform Schwannoma|9560/0
C0027809|T191|PT|C3269|NCI|Schwannoma|9560/0
C0027809|T191|SY|TCGA|NCI|Schwannoma|9560/0
C0027809|T191|SY|C3269|NCI_CDISC|Neurilemmoma|9560/0
C0027809|T191|SY|C3269|NCI_CDISC|Neurinoma|9560/0
C0027809|T191|SY|C3269|NCI_CDISC|Schwannoma|9560/0
C0027809|T191|PT|C3269|NCI_CDISC|SCHWANNOMA, BENIGN|9560/0
C0027809|T191|PT|CDR0000046572|NCI_NCI-GLOSS|schwannoma|9560/0
C0431124|T191|PT|X77po|RCD|Cellular Schwannoma|9560/0
C0027809|T191|SY|Xa99U|RCD|Neurilemmoma|9560/0
C0027809|T191|SY|Xa99U|RCD|Neurinoma|9560/0
C1370659|T191|PT|X77pp|RCD|Plexiform Schwannoma|9560/0
C0027809|T191|PT|Xa99U|RCD|Schwannoma|9560/0
C0027809|T191|SY|Xa99U|RCDAE|Neurilemoma|9560/0
C1536561|T191|SY|404023006|SNOMEDCT_US|Ancient neurilemmoma|9560/0
C1536561|T191|SYGB|409704009|SNOMEDCT_US|Ancient neurilemmoma|9560/0
C1536561|T191|SY|409704009|SNOMEDCT_US|Ancient neurilemoma|9560/0
C1536561|T191|IS|985004|SNOMEDCT_US|Ancient schwannoma|9560/0
C1536561|T191|IS|404023006|SNOMEDCT_US|Ancient Schwannoma|9560/0
C1536561|T191|PT|404023006|SNOMEDCT_US|Ancient schwannoma|9560/0
C1536561|T191|PT|409704009|SNOMEDCT_US|Ancient schwannoma|9560/0
C0431124|T191|SY|253086004|SNOMEDCT_US|Cellular neurilemmoma|9560/0
C0431124|T191|SY|404026003|SNOMEDCT_US|Cellular neurilemmoma|9560/0
C0431124|T191|OP|253086004|SNOMEDCT_US|Cellular Schwannoma|9560/0
C0431124|T191|PT|404026003|SNOMEDCT_US|Cellular schwannoma|9560/0
C0431124|T191|PT|253086004|SNOMEDCT_US|Cellular schwannoma|9560/0
C0431124|T191|IS|985004|SNOMEDCT_US|Cellular schwannoma|9560/0
C1536561|T191|IS|985004|SNOMEDCT_US|Degenerated schwannoma|9560/0
C0027809|T191|SY|985004|SNOMEDCT_US|Neurilemmoma|9560/0
C0027809|T191|SY|189948006|SNOMEDCT_US|Neurilemmoma|9560/0
C0027809|T191|OAP|404022001|SNOMEDCT_US|Neurilemmoma|9560/0
C0027809|T191|IS|985004|SNOMEDCT_US|Neurilemmoma, NOS|9560/0
C0027809|T191|OAS|404022001|SNOMEDCT_US|Neurilemoma|9560/0
C0027809|T191|SY|985004|SNOMEDCT_US|Neurilemoma|9560/0
C0027809|T191|SY|985004|SNOMEDCT_US|Neurinoma|9560/0
C1370659|T191|SY|404025004|SNOMEDCT_US|Plexiform neurilemmoma|9560/0
C1370659|T191|SY|253087008|SNOMEDCT_US|Plexiform neurilemmoma|9560/0
C1370659|T191|PT|404025004|SNOMEDCT_US|Plexiform schwannoma|9560/0
C1370659|T191|PT|253087008|SNOMEDCT_US|Plexiform schwannoma|9560/0
C1370659|T191|IS|404025004|SNOMEDCT_US|Plexiform Schwannoma|9560/0
C1370659|T191|IS|985004|SNOMEDCT_US|Plexiform schwannoma|9560/0
C1370659|T191|OP|253087008|SNOMEDCT_US|Plexiform Schwannoma|9560/0
C0027809|T191|SY|985004|SNOMEDCT_US|Psammomatous schwannoma|9560/0
C0027809|T191|PT|189948006|SNOMEDCT_US|Schwannoma|9560/0
C0027809|T191|PT|985004|SNOMEDCT_US|Schwannoma|9560/0
C0027809|T191|OAS|404022001|SNOMEDCT_US|Schwannoma|9560/0
C0027809|T191|OF|189948006|SNOMEDCT_US|Schwannoma|9560/0
C0027809|T191|IS|985004|SNOMEDCT_US|Schwannoma, NOS|9560/0
C1265858|T191|PT|125351005|SNOMEDCT_US|Verocay body|9560/0
C1306247|T191|SY|0000057856|CHV|melanocytic schwannoma|9560/1
C1306247|T191|PT|0000057856|CHV|melanotic schwannoma|9560/1
C1335929|T191|AB|Q85.03|ICD10CM|Schwannomatosis|9560/1
C1335929|T191|PT|Q85.03|ICD10CM|Schwannomatosis|9560/1
C1335929|T191|AB|237.73|ICD9CM|Schwannomatosis|9560/1
C1335929|T191|PT|237.73|ICD9CM|Schwannomatosis|9560/1
C1335929|T191|PT|314591|MEDCIN|schwannomatosis|9560/1
C1335929|T191|NM|C536641|MSH|Schwannomatosis|9560/1
C1335929|T191|PN|NOCODE|MTH|Schwannomatosis|9560/1
C1306247|T191|SY|C6970|NCI|Melanocytic Neurilemmoma|9560/1
C1306247|T191|SY|C6970|NCI|Melanocytic Schwannoma|9560/1
C1306247|T191|SY|C6970|NCI|Melanotic Neurilemmoma|9560/1
C1306247|T191|SY|C6970|NCI|Melanotic Neurinoma|9560/1
C1306247|T191|PT|C6970|NCI|Melanotic Schwannoma|9560/1
C1306247|T191|SY|TCGA|NCI|Melanotic Schwannoma|9560/1
C1335929|T191|SY|C6557|NCI|Neurilemmomatosis|9560/1
C1335929|T191|SY|C6557|NCI|Neurinomatosis|9560/1
C1306247|T191|SY|C6970|NCI|Pigmented Neurilemmoma|9560/1
C1306247|T191|SY|C6970|NCI|Pigmented Schwannoma|9560/1
C1335929|T191|PT|C6557|NCI|Schwannomatosis|9560/1
C1335929|T191|PT|C6557|NCI_CPTAC|Schwannomatosis|9560/1
C1335929|T191|SY|CDR0000751907|PDQ|neurilemmomatosis|9560/1
C1335929|T191|SY|CDR0000751907|PDQ|neurinomatosis|9560/1
C1335929|T191|PT|CDR0000751907|PDQ|schwannomatosis|9560/1
C1306247|T191|PT|X77pq|RCD|Melanotic Schwannoma|9560/1
C1306247|T191|SY|X77pq|RCD|Pigmented Schwannoma|9560/1
C1335929|T191|OP|BBe6.|RCDSY|Neurinomatosis|9560/1
C1306247|T191|IS|985004|SNOMEDCT_US|Melanocytic Schwannoma|9560/1
C1306247|T191|SY|253088003|SNOMEDCT_US|Melanotic neurilemmoma|9560/1
C1306247|T191|SY|404024000|SNOMEDCT_US|Melanotic neurilemmoma|9560/1
C1306247|T191|IS|985004|SNOMEDCT_US|Melanotic schwannoma|9560/1
C1306247|T191|OP|253088003|SNOMEDCT_US|Melanotic Schwannoma|9560/1
C1306247|T191|PT|253088003|SNOMEDCT_US|Melanotic schwannoma|9560/1
C1306247|T191|PT|404024000|SNOMEDCT_US|Melanotic schwannoma|9560/1
C1335929|T191|SY|781641005|SNOMEDCT_US|Neurilemmomatosis|9560/1
C1335929|T191|OAP|72080001|SNOMEDCT_US|Neurinomatosis|9560/1
C1306247|T191|IS|985004|SNOMEDCT_US|Pigmented Schawnnoma|9560/1
C1306247|T191|IS|985004|SNOMEDCT_US|Pigmented schwannoma|9560/1
C1306247|T191|IS|253088003|SNOMEDCT_US|Pigmented Schwannoma|9560/1
C1306247|T191|SY|253088003|SNOMEDCT_US|Pigmented schwannoma|9560/1
C1335929|T191|OAP|142071000119101|SNOMEDCT_US|Schwannomatosis|9560/1
C1335929|T191|PT|781641005|SNOMEDCT_US|Schwannomatosis|9560/1
C0751690|T191|PT|0000048479|CHV|malignant schwannoma|9560/3
C0751690|T191|PT|0000045030|CHV|malignant schwannoma|9560/3
C0751690|T191|SY|0000048479|CHV|mpnst|9560/3
C0751690|T191|SY|HP:0100697|HPO|Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|SY|HP:0100697|HPO|Malignant schwannoma|9560/3
C0751690|T191|LLT|10026667|MDR|Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|LLT|10073836|MDR|Malignant peripheral nerve sheath tumour|9560/3
C0751690|T191|LLT|10029236|MDR|Neurilemmoma malignant|9560/3
C0751690|T191|LLT|10029239|MDR|Neurilemoma malignant|9560/3
C0751690|T191|LLT|10034589|MDR|Peripheral nerve sheath tumor malignant|9560/3
C0751690|T191|LLT|10034590|MDR|Peripheral nerve sheath tumour malignant|9560/3
C0751690|T191|LLT|10058387|MDR|Schwannoma malignant|9560/3
C0751690|T191|PT|271574|MEDCIN|malignant neurilemoma|9560/3
C0751690|T191|SY|271571|MEDCIN|malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|SY|271571|MEDCIN|MPNST|9560/3
C0751690|T191|ET|D018319|MSH|Malignant Neurilemmoma|9560/3
C0751690|T191|PM|D018319|MSH|Malignant Neurilemmomas|9560/3
C0751690|T191|ET|D018319|MSH|Malignant Neurilemoma|9560/3
C0751690|T191|PM|D018319|MSH|Malignant Neurilemomas|9560/3
C0751690|T191|ET|D018319|MSH|Malignant Peripheral Nerve Sheath Tumor|9560/3
C0751690|T191|PEP|D018319|MSH|Malignant Peripheral Nerve Sheath Tumors|9560/3
C0751690|T191|PM|D018319|MSH|Malignant Schwannoma|9560/3
C0751690|T191|PM|D018319|MSH|Malignant Schwannomas|9560/3
C0751690|T191|ET|D018319|MSH|MPNST|9560/3
C0751690|T191|PM|D018319|MSH|Neurilemmoma, Malignant|9560/3
C0751690|T191|ET|D018319|MSH|Neurilemmosarcoma|9560/3
C0751690|T191|PM|D018319|MSH|Neurilemmosarcomas|9560/3
C0751690|T191|PM|D018319|MSH|Neurilemoma, Malignant|9560/3
C0751690|T191|ET|D018319|MSH|Peripheral Nerve Sheath Tumors, Malignant|9560/3
C0751690|T191|ET|D018319|MSH|Schwannoma, Malignant|9560/3
C0751690|T191|PN|NOCODE|MTH|Malignant Peripheral Nerve Sheath Tumor|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Neoplasm of Peripheral Nerve Sheath|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Neoplasm of the Peripheral Nerve Sheath|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Neurilemmoma|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Neurilemoma|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Peripheral Nerve Sheath Neoplasm|9560/3
C0751690|T191|PT|C3798|NCI|Malignant Peripheral Nerve Sheath Tumor|9560/3
C0751690|T191|SY|TCGA|NCI|Malignant Peripheral Nerve Sheath Tumor|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Peripheral Nerve Sheath Tumour|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Schwannoma|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Tumor of Peripheral Nerve Sheath|9560/3
C0751690|T191|SY|C3798|NCI|Malignant Tumor of the Peripheral Nerve Sheath|9560/3
C0751690|T191|AB|C3798|NCI|MPNST|9560/3
C0751690|T191|SY|C3798|NCI|Neurofibrosarcoma|9560/3
C0751690|T191|SY|C3798|NCI|Neurogenic Sarcoma|9560/3
C0751690|T191|SY|C3798|NCI_CDISC|Malignant Neurilemmoma|9560/3
C0751690|T191|SY|C3798|NCI_CDISC|Malignant Peripheral Nerve Sheath Tumour|9560/3
C0751690|T191|SY|C3798|NCI_CDISC|Neurofibrosarcoma, Malignant|9560/3
C0751690|T191|PT|C3798|NCI_CDISC|SCHWANNOMA, MALIGNANT|9560/3
C0751690|T191|PT|C3798|NCI_CPTAC|Malignant Peripheral Nerve Sheath Tumor|9560/3
C0751690|T191|SY|10026667|NCI_CTEP-SDC|Malig. periph. nerve sheath tum.|9560/3
C0751690|T191|PT|10026667|NCI_CTEP-SDC|Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|PT|CDR0000335496|NCI_NCI-GLOSS|malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|PT|CDR0000335498|NCI_NCI-GLOSS|MPNST|9560/3
C0751690|T191|AB|Xa99V|RCD|Malig periph nerve sheath tum|9560/3
C0751690|T191|OP|BBe7.|RCD|Malignant neurilemmoma|9560/3
C0751690|T191|PT|Xa99V|RCD|Malignant peripheral nerve sheath tumour|9560/3
C0751690|T191|SY|Xa99V|RCD|Malignant Schwannoma|9560/3
C0751690|T191|SY|Xa99V|RCD|MPNST - Malignant peripheral nerve sheath tumour|9560/3
C0751690|T191|AB|Xa99V|RCD|MPNST-Mal perip ner sheath tum|9560/3
C0751690|T191|SY|Xa99V|RCD|Neurilemmosarcoma|9560/3
C0751690|T191|OP|BBe7.|RCDAE|Malignant neurilemoma|9560/3
C0751690|T191|PT|Xa99V|RCDAE|Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|SY|Xa99V|RCDAE|MPNST - Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|SYGB|404037002|SNOMEDCT_US|Malignant neurilemmoma|9560/3
C0751690|T191|OAP|189949003|SNOMEDCT_US|Malignant neurilemmoma|9560/3
C0751690|T191|OF|189949003|SNOMEDCT_US|Malignant neurilemmoma|9560/3
C0751690|T191|SY|404037002|SNOMEDCT_US|Malignant neurilemoma|9560/3
C0751690|T191|PT|404037002|SNOMEDCT_US|Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|PT|19897006|SNOMEDCT_US|Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|OAP|134324009|SNOMEDCT_US|Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|OAP|134324009|SNOMEDCT_US|Malignant peripheral nerve sheath tumour|9560/3
C0751690|T191|PTGB|404037002|SNOMEDCT_US|Malignant peripheral nerve sheath tumour|9560/3
C0751690|T191|PTGB|19897006|SNOMEDCT_US|Malignant peripheral nerve sheath tumour|9560/3
C0751690|T191|SY|404037002|SNOMEDCT_US|Malignant schwannoma|9560/3
C0751690|T191|OAS|77418004|SNOMEDCT_US|Malignant Schwannoma|9560/3
C0751690|T191|IS|77418004|SNOMEDCT_US|Malignant Schwannoma, NOS|9560/3
C0751690|T191|IS|19897006|SNOMEDCT_US|MPNST|9560/3
C0751690|T191|OAS|134324009|SNOMEDCT_US|MPNST - Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|SY|19897006|SNOMEDCT_US|MPNST - Malignant peripheral nerve sheath tumor|9560/3
C0751690|T191|OAS|134324009|SNOMEDCT_US|MPNST - Malignant peripheral nerve sheath tumour|9560/3
C0751690|T191|SYGB|19897006|SNOMEDCT_US|MPNST - Malignant peripheral nerve sheath tumour|9560/3
C0751690|T191|OAS|77418004|SNOMEDCT_US|Neurilemmoma, malignant|9560/3
C0751690|T191|OAS|77418004|SNOMEDCT_US|Neurilemmosarcoma|9560/3
C0751690|T191|OAP|77418004|SNOMEDCT_US|Neurilemoma, malignant|9560/3
C0334616|T191|PT|355155|MEDCIN|malignant Triton tumor|9561/3
C0334616|T191|SY|C4335|NCI|Malignant Neoplasm of Peripheral Nerve Sheath with Rhabdomyosarcoma|9561/3
C0334616|T191|SY|C4335|NCI|Malignant Neoplasm of the Peripheral Nerve Sheath with Rhabdomyosarcoma|9561/3
C0334616|T191|SY|C4335|NCI|Malignant Peripheral Nerve Sheath Neoplasm with Rhabdomyosarcoma|9561/3
C0334616|T191|SY|C4335|NCI|Malignant Peripheral Nerve Sheath Tumor with Rhabdomyosarcoma|9561/3
C0334616|T191|PT|C4335|NCI|Malignant Triton Tumor|9561/3
C0334616|T191|SY|C4335|NCI|Malignant Tumor of Peripheral Nerve Sheath with Rhabdomyosarcoma|9561/3
C0334616|T191|SY|C4335|NCI|Malignant Tumor of the Peripheral Nerve Sheath with Rhabdomyosarcoma|9561/3
C0334616|T191|SY|C4335|NCI|MPNST with Rhabdomyosarcoma|9561/3
C0334616|T191|AB|X77pw|RCD|Malig Schwannoma+rhabdomy diff|9561/3
C0334616|T191|SY|X77pw|RCD|Malignant Schwannoma with rhabdomyoblastic differentiation|9561/3
C0334616|T191|PT|X77pw|RCD|Malignant Triton tumour|9561/3
C0334616|T191|PT|X77pw|RCDAE|Malignant Triton tumor|9561/3
C0334616|T191|SY|X77pw|RCDSA|Triton tumor, malignant|9561/3
C0334616|T191|SY|X77pw|RCDSY|Triton tumour, malignant|9561/3
C0334616|T191|SY|354002|SNOMEDCT_US|Malignant neurilemmoma with rhabdomyoblastic differentiation|9561/3
C0334616|T191|PT|354002|SNOMEDCT_US|Malignant peripheral nerve sheath tumor with rhabdomyoblastic differentiation|9561/3
C0334616|T191|PTGB|354002|SNOMEDCT_US|Malignant peripheral nerve sheath tumour with rhabdomyoblastic differentiation|9561/3
C0334616|T191|IS|354002|SNOMEDCT_US|Malignant Schwannoma with rhabdomyoblastic differentiation|9561/3
C0334616|T191|SY|354002|SNOMEDCT_US|Malignant schwannoma with rhabdomyoblastic differentiation|9561/3
C0334616|T191|PT|404040002|SNOMEDCT_US|Malignant Triton tumor|9561/3
C0334616|T191|OAP|189951004|SNOMEDCT_US|Malignant Triton tumor|9561/3
C0334616|T191|PTGB|404040002|SNOMEDCT_US|Malignant Triton tumour|9561/3
C0334616|T191|OAP|189951004|SNOMEDCT_US|Malignant Triton tumour|9561/3
C0334616|T191|OF|189951004|SNOMEDCT_US|Malignant Triton tumour|9561/3
C0334616|T191|SY|354002|SNOMEDCT_US|MPNST with rhabdomyoblastic differentiation|9561/3
C0334616|T191|SY|354002|SNOMEDCT_US|Triton tumor, malignant|9561/3
C0334616|T191|SYGB|354002|SNOMEDCT_US|Triton tumour, malignant|9561/3
C0206730|T191|SY|0000021054|CHV|nerve sheath myxoma|9562/0
C0206730|T191|SY|0000021054|CHV|neurothecoma|9562/0
C0206730|T191|PT|0000021054|CHV|neurothekeoma|9562/0
C0206730|T191|ET|2012-6947|CSP|neurothekeoma|9562/0
C0206730|T191|ET|D018321|MSH|Myxoma, Nerve Sheath|9562/0
C0206730|T191|PM|D018321|MSH|Myxomas, Nerve Sheath|9562/0
C0206730|T191|PM|D018321|MSH|Nerve Sheath Myxoma|9562/0
C0206730|T191|PM|D018321|MSH|Nerve Sheath Myxomas|9562/0
C0206730|T191|ET|D018321|MSH|Neurotheceoma|9562/0
C0206730|T191|PM|D018321|MSH|Neurotheceomas|9562/0
C0206730|T191|ET|D018321|MSH|Neurothecoma|9562/0
C0206730|T191|PM|D018321|MSH|Neurothecomas|9562/0
C0206730|T191|MH|D018321|MSH|Neurothekeoma|9562/0
C0206730|T191|PM|D018321|MSH|Neurothekeomas|9562/0
C1275959|T191|PT|C156278|NCI|Cellular Neurothekeoma|9562/0
C0206730|T191|SY|C7018|NCI|Nerve Sheath Myxoma|9562/0
C0206730|T191|PT|C7018|NCI|Neurothekeoma|9562/0
C0206730|T191|SY|X77ps|RCD|Lobular neuromyxoma|9562/0
C0206730|T191|PT|X77ps|RCD|Nerve sheath myxoma|9562/0
C0206730|T191|PT|X77pr|RCD|Neurothekeoma|9562/0
C1275959|T191|SY|399922004|SNOMEDCT_US|Cellular nerve sheath myxoma|9562/0
C1275959|T191|PT|399922004|SNOMEDCT_US|Cellular neurothekeoma|9562/0
C0206730|T191|OAS|253089006|SNOMEDCT_US|Lobular neuromyxoma|9562/0
C0206730|T191|SY|51836001|SNOMEDCT_US|Nerve sheath myxoma|9562/0
C0206730|T191|OAP|253089006|SNOMEDCT_US|Nerve sheath myxoma|9562/0
C0206730|T191|OF|253089006|SNOMEDCT_US|Nerve sheath myxoma|9562/0
C0206730|T191|PT|51836001|SNOMEDCT_US|Neurothekeoma|9562/0
C0206730|T191|OAP|189952006|SNOMEDCT_US|Neurothekeoma|9562/0
C0206730|T191|OF|189952006|SNOMEDCT_US|Neurothekeoma|9562/0
C3839433|T191|SY|C121686|NCI|Hybrid Nerve Sheath Neoplasm|9563/0
C3839433|T191|PT|C121686|NCI|Hybrid Nerve Sheath Tumor|9563/0
C3839433|T191|SY|C121686|NCI|Hybrid Neurofibroma-Perineurioma|9563/0
C3839433|T191|SY|C121686|NCI|Hybrid Neurofibroma-Schwannoma|9563/0
C3839433|T191|SY|C121686|NCI|Hybrid Schwannoma-Perineurioma|9563/0
C3839433|T191|SY|C121686|NCI|Nerve Sheath Tumor, NOS|9563/0
C3839433|T191|SY|C121686|NCI|Nerve Sheath Tumor, Not Otherwise Specified|9563/0
C3839433|T191|PT|703710008|SNOMEDCT_US|Hybrid nerve sheath tumor|9563/0
C3839433|T191|PTGB|703710008|SNOMEDCT_US|Hybrid nerve sheath tumour|9563/0
C3839008|T191|PT|703709003|SNOMEDCT_US|Nerve sheath tumor, no ICD-O subtype|9563/0
C3839008|T191|SY|703709003|SNOMEDCT_US|Nerve sheath tumor, no International Classification of Diseases for Oncology subtype|9563/0
C3839008|T191|PTGB|703709003|SNOMEDCT_US|Nerve sheath tumour, no ICD-O subtype|9563/0
C0027858|T191|PT|0000008645|CHV|A tumor made up of nerve cells and nerve fibers|9570/0
C0027858|T191|SY|0000008645|CHV|neuroma|9570/0
C0027858|T191|SY|0000008645|CHV|neuromas|9570/0
C0406848|T191|PT|0000032694|CHV|scar neuroma|9570/0
C0027858|T191|PT|U000477|COSTAR|NEUROMA|9570/0
C0027858|T191|ET|2012-5157|CSP|neuroma|9570/0
C0027858|T191|GT|NEOPL CNS|CST|NEUROMA|9570/0
C0027858|T191|SY|HP:0030430|HPO|Nerve tumor|9570/0
C0027858|T191|PT|HP:0030430|HPO|Neuroma|9570/0
C0027858|T191|PT|N75007|ICPC2P|Neuroma|9570/0
C0027858|T191|PTN|N75007|ICPC2P|neuroma|9570/0
C0027858|T191|PT|sh92003433|LCH_NW|Neuromas|9570/0
C0027858|T191|PT|10029308|MDR|Neuroma|9570/0
C0027858|T191|LLT|10029308|MDR|Neuroma|9570/0
C0027858|T191|LLT|10029310|MDR|Neuroma NOS|9570/0
C0027858|T191|HT|10029312|MDR|Neuromas|9570/0
C0027858|T191|MH|D009463|MSH|Neuroma|9570/0
C0027858|T191|PM|D009463|MSH|Neuromas|9570/0
C0027858|T191|PT|C3275|NCI|Neuroma|9570/0
C0431126|T191|SY|C121681|NCI|Palisaded Encapsulated Neuroma|9570/0
C0431126|T191|PT|C121681|NCI|Solitary Circumscribed Neuroma|9570/0
C0027858|T191|PT|CDR0000046268|NCI_NCI-GLOSS|neuroma|9570/0
C0027858|T191|PT|Xa99W|RCD|Neuroma|9570/0
C0406848|T191|PT|X50LC|RCD|Scar neuroma|9570/0
C0431126|T191|PT|X77pu|RCD|Solitary circumscribed neuroma|9570/0
C0027858|T191|OP|BBe8.|RCDSY|Neuroma NOS|9570/0
C0027858|T191|SY|25169009|SNOMEDCT_US|Neuroma|9570/0
C0027858|T191|PT|443892003|SNOMEDCT_US|Neuroma|9570/0
C2732416|T191|PT|443818003|SNOMEDCT_US|Neuroma - category|9570/0
C0027858|T191|PT|25169009|SNOMEDCT_US|Neuroma, no ICD-O subtype|9570/0
C0027858|T191|SY|25169009|SNOMEDCT_US|Neuroma, no International Classification of Diseases for Oncology subtype|9570/0
C0027858|T191|IS|25169009|SNOMEDCT_US|Neuroma, NOS|9570/0
C0431126|T191|PT|404019003|SNOMEDCT_US|Palisaded encapsulated neuroma|9570/0
C0406848|T191|PT|371432009|SNOMEDCT_US|Scar neuroma|9570/0
C0406848|T191|PT|239178001|SNOMEDCT_US|Scar neuroma|9570/0
C0431126|T191|SY|404019003|SNOMEDCT_US|Solitary circumscribed neuroma|9570/0
C0431126|T191|PT|253091003|SNOMEDCT_US|Solitary circumscribed neuroma|9570/0
C0027858|T191|PT|1344|WHO|NEUROMA|9570/0
C0751691|T191|LA|LA26520-9|LNC|Perineurioma, NOS|9571/0
C0751691|T191|PEP|D018317|MSH|Perineurioma|9571/0
C0751691|T191|PM|D018317|MSH|Perineuriomas|9571/0
C0751691|T191|PN|NOCODE|MTH|Perineurioma|9571/0
C0751691|T191|PT|C4973|NCI|Perineurioma|9571/0
C0751691|T191|PT|404036006|SNOMEDCT_US|Perineurioma|9571/0
C0751691|T191|PT|128795001|SNOMEDCT_US|Perineurioma|9571/0
C1266188|T191|PT|271573|MEDCIN|malignant perineurioma|9571/3
C1266188|T191|SY|C66845|NCI|Malignant Perineurioma|9571/3
C1266188|T191|PT|C66845|NCI|Malignant Peripheral Nerve Sheath Tumor with Perineurial Differentiation|9571/3
C1266188|T191|SY|C66845|NCI|Perineurial Malignant Peripheral Nerve Sheath Tumor|9571/3
C1266188|T191|PT|761958009|SNOMEDCT_US|Malignant perineurioma|9571/3
C1266188|T191|OAP|734069003|SNOMEDCT_US|Malignant peripheral nerve sheath neoplasm with perineurial differentiation|9571/3
C1266188|T191|SY|761958009|SNOMEDCT_US|Malignant peripheral nerve sheath neoplasm with perineurial differentiation|9571/3
C1266188|T191|SY|128796000|SNOMEDCT_US|Malignant peripheral nerve sheath neoplasm with perineurial differentiation|9571/3
C1266188|T191|SY|761958009|SNOMEDCT_US|Malignant peripheral nerve sheath tumor with perineurial differentiation|9571/3
C1266188|T191|SYGB|761958009|SNOMEDCT_US|Malignant peripheral nerve sheath tumour with perineurial differentiation|9571/3
C1266188|T191|IS|128796000|SNOMEDCT_US|Perineural MPNST|9571/3
C1266188|T191|PT|128796000|SNOMEDCT_US|Perineurioma, malignant|9571/3
C0085167|T191|PT|0055864|CCPSS|GRANULAR CELL TUMOR|9580/0
C0085167|T191|SY|0000015475|CHV|cells granular tumor|9580/0
C0085167|T191|SY|0000015475|CHV|granular cell myoblastoma|9580/0
C0085167|T191|SY|0000015475|CHV|granular cell myoblastomas|9580/0
C0085167|T191|PT|0000015475|CHV|granular cell tumor|9580/0
C0085167|T191|SY|0000015475|CHV|granular cell tumors|9580/0
C0085167|T191|SY|0000015475|CHV|granular cell tumour|9580/0
C0085167|T191|LA|LA26522-5|LNC|Granular cell tumor, NOS|9580/0
C0085167|T191|MTH_PT|10060980|MDR|Granular cell tumor|9580/0
C0085167|T191|LLT|10060982|MDR|Granular cell tumor|9580/0
C0085167|T191|LLT|10060980|MDR|Granular cell tumour|9580/0
C0085167|T191|PT|10060980|MDR|Granular cell tumour|9580/0
C0085167|T191|PT|271577|MEDCIN|granular cell tumor|9580/0
C0085167|T191|SY|271577|MEDCIN|malignant granular cell tumor|9580/0
C0085167|T191|PM|D016586|MSH|Cell Myoblastoma, Granular|9580/0
C0085167|T191|PM|D016586|MSH|Cell Myoblastomas, Granular|9580/0
C0085167|T191|PM|D016586|MSH|Cell Tumor, Granular|9580/0
C0085167|T191|PM|D016586|MSH|Cell Tumors, Granular|9580/0
C0085167|T191|ET|D016586|MSH|Granular Cell Myoblastoma|9580/0
C0085167|T191|PM|D016586|MSH|Granular Cell Myoblastomas|9580/0
C0085167|T191|MH|D016586|MSH|Granular Cell Tumor|9580/0
C0085167|T191|PM|D016586|MSH|Granular Cell Tumors|9580/0
C0085167|T191|ET|D016586|MSH|Myoblastoma, Granular Cell|9580/0
C0085167|T191|PM|D016586|MSH|Myoblastomas, Granular Cell|9580/0
C0085167|T191|PM|D016586|MSH|Tumor, Granular Cell|9580/0
C0085167|T191|PM|D016586|MSH|Tumors, Granular Cell|9580/0
C0085167|T191|PN|NOCODE|MTH|Granular cell tumor|9580/0
C0085167|T191|SY|C3474|NCI|Abrikossoff Tumor|9580/0
C0085167|T191|SY|C3474|NCI|Abrikossoff's Tumor|9580/0
C0085167|T191|SY|C3474|NCI|Granular Cell Myoblastoma|9580/0
C0085167|T191|SY|C3474|NCI|Granular Cell Neoplasm|9580/0
C0085167|T191|SY|C3474|NCI|Granular Cell Nerve Sheath Tumor|9580/0
C0085167|T191|SY|C3474|NCI|Granular Cell Schwannoma|9580/0
C0085167|T191|PT|C3474|NCI|Granular Cell Tumor|9580/0
C0085167|T191|SY|Xa99d|RCD|Granular cell myoblastoma|9580/0
C0085167|T191|PT|Xa99d|RCD|Granular cell tumour|9580/0
C0085167|T191|PT|Xa99d|RCDAE|Granular cell tumor|9580/0
C0085167|T191|OP|BBf0.|RCDSA|Granular cell tumor NOS|9580/0
C0085167|T191|OP|BBf0.|RCDSY|Granular cell tumour NOS|9580/0
C0085167|T191|SY|404035005|SNOMEDCT_US|Abrikossoff's tumor|9580/0
C0085167|T191|SYGB|404035005|SNOMEDCT_US|Abrikossoff's tumour|9580/0
C0085167|T191|SY|404035005|SNOMEDCT_US|Granular cell myoblastoma|9580/0
C0085167|T191|SY|12169001|SNOMEDCT_US|Granular cell myoblastoma|9580/0
C0085167|T191|IS|12169001|SNOMEDCT_US|Granular cell myoblastoma, NOS|9580/0
C0085167|T191|PT|12169001|SNOMEDCT_US|Granular cell tumor|9580/0
C0085167|T191|PT|404035005|SNOMEDCT_US|Granular cell tumor|9580/0
C0085167|T191|IS|12169001|SNOMEDCT_US|Granular cell tumor, NOS|9580/0
C0085167|T191|PTGB|404035005|SNOMEDCT_US|Granular cell tumour|9580/0
C0085167|T191|PTGB|12169001|SNOMEDCT_US|Granular cell tumour|9580/0
C0334618|T191|PT|355159|MEDCIN|malignant granular cell neoplasm|9580/3
C0334618|T191|SY|355159|MEDCIN|neoplasm of nerve sheath origin malignant granular cell|9580/3
C0334618|T191|PN|NOCODE|MTH|Malignant granular cell tumor|9580/3
C0334618|T191|SY|C4336|NCI|Malignant Granular Cell Myoblastoma|9580/3
C0334618|T191|SY|C4336|NCI|Malignant Granular Cell Neoplasm|9580/3
C0334618|T191|PT|C4336|NCI|Malignant Granular Cell Tumor|9580/3
C0334618|T191|PT|C4336|NCI_CDISC|GRANULAR CELL TUMOR, MALIGNANT|9580/3
C0334618|T191|SY|C4336|NCI_CDISC|Malignant Granular Cell Myoblastoma|9580/3
C0334618|T191|SY|C4336|NCI_CDISC|Malignant Granular Cell Neoplasm|9580/3
C0334618|T191|SY|C4336|NCI_CDISC|Myoblastoma, Malignant|9580/3
C0334618|T191|AB|BBf1.|RCD|Malig granul cell myoblastoma|9580/3
C0334618|T191|SY|BBf1.|RCD|Malignant granular cell myoblastoma|9580/3
C0334618|T191|PT|BBf1.|RCD|Malignant granular cell tumour|9580/3
C0334618|T191|PT|BBf1.|RCDAE|Malignant granular cell tumor|9580/3
C0334618|T191|SY|13238004|SNOMEDCT_US|Granular cell myoblastoma, malignant|9580/3
C0334618|T191|PT|13238004|SNOMEDCT_US|Granular cell tumor, malignant|9580/3
C0334618|T191|PTGB|13238004|SNOMEDCT_US|Granular cell tumour, malignant|9580/3
C0334618|T191|SY|13238004|SNOMEDCT_US|Malignant granular cell myoblastoma|9580/3
C0334618|T191|PT|404041003|SNOMEDCT_US|Malignant granular cell tumor|9580/3
C0334618|T191|SY|13238004|SNOMEDCT_US|Malignant granular cell tumor|9580/3
C0334618|T191|PTGB|404041003|SNOMEDCT_US|Malignant granular cell tumour|9580/3
C0334618|T191|SYGB|13238004|SNOMEDCT_US|Malignant granular cell tumour|9580/3
C0206657|T191|PT|0033728|CCPSS|ALVEOLAR SOFT PART SARCOMA|9581/3
C0206657|T191|PT|HP:0012218|HPO|Alveolar soft part sarcoma|9581/3
C0206657|T191|PT|MTHU005108|ICPC2ICD10ENG|alveolar; soft part sarcoma|9581/3
C0206657|T191|PT|MTHU065885|ICPC2ICD10ENG|sarcoma; alveolar, soft part|9581/3
C0206657|T191|PT|10001882|MDR|Alveolar soft part sarcoma|9581/3
C0206657|T191|LLT|10001882|MDR|Alveolar soft part sarcoma|9581/3
C0206657|T191|LLT|10001886|MDR|Alveolar soft part sarcoma NOS|9581/3
C0206657|T191|HT|10001883|MDR|Alveolar soft part sarcomas|9581/3
C0206657|T191|PT|271502|MEDCIN|alveolar soft part sarcoma|9581/3
C0206657|T191|PT|231896|MEDCIN|alveolar soft part sarcoma of soft tissue|9581/3
C0206657|T191|ET|D018234|MSH|Alveolar Soft Part Sarcoma|9581/3
C0206657|T191|ET|D018234|MSH|Alveolar Soft-Part Sarcoma|9581/3
C0206657|T191|MH|D018234|MSH|Sarcoma, Alveolar Soft Part|9581/3
C0206657|T191|PN|NOCODE|MTH|Alveolar Soft Part Sarcoma|9581/3
C0206657|T191|PT|C3750|NCI|Alveolar Soft Part Sarcoma|9581/3
C0206657|T191|AB|C3750|NCI|ASPS|9581/3
C0206657|T191|PT|10001886|NCI_CTEP-SDC|Alveolar soft part sarcoma|9581/3
C0206657|T191|DN|C3750|NCI_CTRP|Alveolar Soft Part Sarcoma|9581/3
C0206657|T191|PT|CDR0000641933|NCI_NCI-GLOSS|alveolar soft part sarcoma|9581/3
C0206657|T191|PT|CDR0000641934|NCI_NCI-GLOSS|ASPS|9581/3
C0206657|T191|PT|Xa99f|RCD|Alveolar soft tissue sarcoma|9581/3
C0206657|T191|OP|BBf2.|RCDSY|Alveolar soft part sarcoma|9581/3
C0206657|T191|PT|88195001|SNOMEDCT_US|Alveolar soft part sarcoma|9581/3
C0206657|T191|PT|404056007|SNOMEDCT_US|Alveolar soft part sarcoma|9581/3
C0206657|T191|OAP|302839003|SNOMEDCT_US|Alveolar soft tissue sarcoma|9581/3
C1333873|T191|PN|NOCODE|MTH|Granular Cell Tumor of the Neurohypophysis|9582/0
C1266189|T191|PN|NOCODE|MTH|Granular cell tumor of the sellar region|9582/0
C1333873|T191|SY|C7017|NCI|Granular Cell Tumor of Neurohypophysis|9582/0
C1333873|T191|SY|C7017|NCI|Granular Cell Tumor of the Neurohypophysis|9582/0
C1333873|T191|SY|C7017|NCI|Granular Cell Tumor of the Posterior Pituitary Gland|9582/0
C1333873|T191|PT|C7017|NCI|Granular Cell Tumor of the Sellar Region|9582/0
C1333873|T191|PT|699331002|SNOMEDCT_US|Granular cell tumor of neurohypophysis|9582/0
C1333873|T191|SY|699331002|SNOMEDCT_US|Granular cell tumor of posterior pituitary|9582/0
C1266189|T191|PT|128797009|SNOMEDCT_US|Granular cell tumor of the sellar region|9582/0
C1333873|T191|PTGB|699331002|SNOMEDCT_US|Granular cell tumour of neurohypophysis|9582/0
C1333873|T191|SYGB|699331002|SNOMEDCT_US|Granular cell tumour of posterior pituitary|9582/0
C1266189|T191|PTGB|128797009|SNOMEDCT_US|Granular cell tumour of the sellar region|9582/0
C0024299|T191|ET|0000004624|AOD|lymphoma|9590/3
C0024299|T191|SY|BI00323|BI|lymphoma|9590/3
C0024305|T191|AB|BI00323|BI|nhl|9590/3
C0024305|T191|PT|BI00323|BI|non-hodgkin's lymphoma|9590/3
C0024299|T191|PT|1017994|CCPSS|LYMPHOMA|9590/3
C0024305|T191|PT|0001640|CCPSS|LYMPHOMA NON HODGKIN|9590/3
C0024305|T191|SD|38|CCS|Non-Hodgkin`s lymphoma|9590/3
C0024305|T191|MD|2.10.2|CCS|Non-Hodgkins lymphoma|9590/3
C0024305|T191|SD|NEO058|CCSR_10|Non-Hodgkin lymphoma|9590/3
C0024299|T191|PT|0000007617|CHV|lymphoma|9590/3
C0024299|T191|SY|0000007617|CHV|lymphoma malignant|9590/3
C0024299|T191|SY|0000007617|CHV|lymphomas|9590/3
C0024299|T191|SY|0000007617|CHV|lymphomas malignant|9590/3
C0024299|T191|SY|0000007617|CHV|malignant lymphoma|9590/3
C0024299|T191|SY|0000007617|CHV|malignant lymphomas|9590/3
C0024305|T191|SY|0000007621|CHV|nhl|9590/3
C0024305|T191|SY|0000007621|CHV|non hodgkin lymphoma|9590/3
C0024305|T191|SY|0000007621|CHV|non hodgkin's lymphoma|9590/3
C0024305|T191|SY|0000007621|CHV|non hodgkins lymphoma|9590/3
C0024305|T191|SY|0000007621|CHV|non-hodgkin lymphoma|9590/3
C0024305|T191|SY|0000007621|CHV|non-hodgkin's lymphoma|9590/3
C0024305|T191|SY|0000007621|CHV|non-hodgkins lymphoma|9590/3
C0024305|T191|SY|0000007621|CHV|nonhodgkin lymphoma|9590/3
C0024305|T191|SY|0000007621|CHV|nonhodgkin's lymphoma|9590/3
C0024305|T191|SY|0000007621|CHV|nonhodgkins lymphoma|9590/3
C0024299|T191|PT|462|COSTAR|LYMPHOMA|9590/3
C0024305|T191|PT|U000045|COSTAR|NON HODGKINS LYMPHOMA|9590/3
C0024305|T191|PT|525|COSTAR|NONHODGKINS LYMPHOMA|9590/3
C0024299|T191|PT|2004-6589|CSP|lymphoma|9590/3
C0024305|T191|PT|4001-0094|CSP|nonHodgkin's lymphoma|9590/3
C0024299|T191|GT|LYMPHOMA LIKE REACT|CST|LYMPHOMA|9590/3
C0024299|T191|GT|LYMPHOMA LIKE REACT|CST|LYMPHOMA MALIGNANT|9590/3
C0024299|T191|FI|U002475|DXP|LYMPHOMA|9590/3
C0024305|T191|SY|NOCODE|DXP|LYMPHOMA, NON HODGKIN|9590/3
C0024305|T191|SY|NOCODE|DXP|NHL|9590/3
C0024305|T191|FI|U002830|DXP|NON-HODGKIN LYMPHOMA|9590/3
C0024299|T191|SY|HP:0002665|HPO|Cancer of lymphatic system|9590/3
C0024299|T191|PT|HP:0002665|HPO|Lymphoma|9590/3
C0024305|T191|PT|HP:0012539|HPO|Non-Hodgkin lymphoma|9590/3
C0024305|T191|PT|C85.9|ICD10|Non-Hodgkin's lymphoma, unspecified type|9590/3
C0024299|T191|ET|C85.9|ICD10CM|Lymphoma NOS|9590/3
C0024299|T191|ET|C85.9|ICD10CM|Malignant lymphoma NOS|9590/3
C0024305|T191|ET|C85.9|ICD10CM|Non-Hodgkin lymphoma NOS|9590/3
C0024305|T191|PT|MTHU023065|ICPC2ICD10ENG|diffuse; lymphoma, small cell, cleaved|9590/3
C0024299|T191|PT|MTHU031393|ICPC2ICD10ENG|germinoblastoma|9590/3
C0024299|T191|PT|MTHU046733|ICPC2ICD10ENG|lymphoma|9590/3
C0024305|T191|PT|MTHU046759|ICPC2ICD10ENG|lymphoma; diffuse, small cell, cleaved|9590/3
C0024305|T191|PT|MTHU046842|ICPC2ICD10ENG|lymphoma; non-Hodgkin's|9590/3
C0024305|T191|PT|MTHU053464|ICPC2ICD10ENG|non-Hodgkin's lymphoma|9590/3
C0024305|T191|PT|MTHU053462|ICPC2ICD10ENG|non-Hodgkin's; lymphoma|9590/3
C0024299|T191|PT|MTHU064357|ICPC2ICD10ENG|reticulolymphosarcoma|9590/3
C0024299|T191|PT|B72002|ICPC2P|Lymphoma|9590/3
C0024299|T191|PTN|B72002|ICPC2P|lymphoma|9590/3
C0024305|T191|PT|B74002|ICPC2P|Lymphoma;non Hodgkins|9590/3
C0024305|T191|PTN|B74002|ICPC2P|non hodgkins lymphoma|9590/3
C0024299|T191|PT|U002766|LCH|Lymphomas|9590/3
C0024299|T191|PT|sh85079154|LCH_NW|Lymphomas|9590/3
C0024299|T191|LA|LA15685-3|LNC|Lymphoma|9590/3
C0024299|T191|LPN|LP266900-2|LNC|Lymphoma|9590/3
C0024299|T191|LLT|10025310|MDR|Lymphoma|9590/3
C0024299|T191|PT|10025310|MDR|Lymphoma|9590/3
C0024299|T191|LLT|10025315|MDR|Lymphoma malignant|9590/3
C0024299|T191|LLT|10025316|MDR|Lymphoma NOS|9590/3
C0024299|T191|LLT|10025632|MDR|Malignant lymphoma|9590/3
C0024299|T191|LLT|10025633|MDR|Malignant lymphoma NOS|9590/3
C0024305|T191|PT|10029547|MDR|Non-Hodgkin's lymphoma|9590/3
C0024305|T191|LLT|10029547|MDR|Non-Hodgkin's lymphoma|9590/3
C0024305|T191|LLT|10029593|MDR|Non-Hodgkin's lymphoma NOS|9590/3
C0024299|T191|SY|36081|MEDCIN|lymphoma|9590/3
C0024299|T191|PT|36081|MEDCIN|malignant lymphoma|9590/3
C0024305|T191|PT|35839|MEDCIN|non-Hodgkin's lymphoma|9590/3
C0024299|T191|PT|117|MEDLINEPLUS|Lymphoma|9590/3
C0024305|T191|ET|117|MEDLINEPLUS|Non-Hodgkin Lymphoma|9590/3
C0024305|T191|SY|117|MEDLINEPLUS|Non-Hodgkin lymphoma|9590/3
C0024305|T191|PM|D008228|MSH|Diffuse Small Cleaved Cell Lymphoma|9590/3
C0024305|T191|DEV|D008228|MSH|DIFFUSE SMALL CLEAVED LYMPHOMA|9590/3
C0024305|T191|ET|D008228|MSH|Diffuse Small Cleaved-Cell Lymphoma|9590/3
C0024299|T191|PM|D008223|MSH|Germinoblastic Sarcoma|9590/3
C0024299|T191|PM|D008223|MSH|Germinoblastic Sarcomas|9590/3
C0024299|T191|ET|D008223|MSH|Germinoblastoma|9590/3
C0024299|T191|PM|D008223|MSH|Germinoblastomas|9590/3
C0024299|T191|MH|D008223|MSH|Lymphoma|9590/3
C0024305|T191|DEV|D008228|MSH|LYMPHOMA SMALL CLEAVED DIFFUSE|9590/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Atypical Diffuse Small Lymphoid|9590/3
C0024299|T191|ET|D008223|MSH|Lymphoma, Malignant|9590/3
C0024305|T191|PM|D008228|MSH|Lymphoma, Non Hodgkin|9590/3
C0024305|T191|PM|D008228|MSH|Lymphoma, Non Hodgkin's|9590/3
C0024305|T191|PM|D008228|MSH|Lymphoma, Non Hodgkins|9590/3
C0024305|T191|MH|D008228|MSH|Lymphoma, Non-Hodgkin|9590/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Non-Hodgkin's|9590/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Non-Hodgkins|9590/3
C0024305|T191|PM|D008228|MSH|Lymphoma, Nonhodgkin|9590/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Nonhodgkin's|9590/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Nonhodgkins|9590/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Small Cleaved Cell, Diffuse|9590/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Small Cleaved-Cell, Diffuse|9590/3
C0024299|T191|PM|D008223|MSH|Lymphomas|9590/3
C0024299|T191|PM|D008223|MSH|Lymphomas, Malignant|9590/3
C0024299|T191|PM|D008223|MSH|Malignant Lymphoma|9590/3
C0024299|T191|PM|D008223|MSH|Malignant Lymphomas|9590/3
C0024305|T191|PM|D008228|MSH|Non Hodgkin Lymphoma|9590/3
C0024305|T191|PM|D008228|MSH|Non Hodgkin's Lymphoma|9590/3
C0024305|T191|ET|D008228|MSH|Non-Hodgkin Lymphoma|9590/3
C0024305|T191|ET|D008228|MSH|Non-Hodgkin's Lymphoma|9590/3
C0024305|T191|PM|D008228|MSH|Non-Hodgkins Lymphoma|9590/3
C0024305|T191|DSV|D008228|MSH|NONHODGKIN LYMPHOMA|9590/3
C0024305|T191|PM|D008228|MSH|Nonhodgkin's Lymphoma|9590/3
C0024305|T191|PM|D008228|MSH|Nonhodgkins Lymphoma|9590/3
C0024299|T191|ET|D008223|MSH|Reticulolymphosarcoma|9590/3
C0024299|T191|PM|D008223|MSH|Reticulolymphosarcomas|9590/3
C0024299|T191|ET|D008223|MSH|Sarcoma, Germinoblastic|9590/3
C0024299|T191|PM|D008223|MSH|Sarcomas, Germinoblastic|9590/3
C0024305|T191|PM|D008228|MSH|Small Cleaved Cell Lymphoma, Diffuse|9590/3
C0024305|T191|DEV|D008228|MSH|SMALL CLEAVED LYMPHOMA DIFFUSE|9590/3
C0024305|T191|ET|D008228|MSH|Small Cleaved-Cell Lymphoma, Diffuse|9590/3
C0024299|T191|PN|NOCODE|MTH|Lymphoma|9590/3
C0024305|T191|PN|NOCODE|MTH|Lymphoma, Non-Hodgkin|9590/3
C0024299|T191|ET|202.8|MTHICD9|Lymphoma NOS|9590/3
C0024299|T191|ET|202.8|MTHICD9|Malignant lymphoma NOS|9590/3
C0024299|T191|ET|200.8|MTHICD9|Reticulolymphosarcoma|9590/3
C0024299|T191|SY|TCGA|NCI|Lymphoma|9590/3
C0024299|T191|PT|C3208|NCI|Lymphoma|9590/3
C0024299|T191|AD|C3208|NCI|Lymphomatous|9590/3
C0024299|T191|SY|C3208|NCI|Malignant Lymphoma|9590/3
C0024305|T191|AB|C3211|NCI|NHL|9590/3
C0024305|T191|PT|C3211|NCI|Non-Hodgkin Lymphoma|9590/3
C0024305|T191|SY|C3211|NCI|Non-Hodgkin's Lymphoma|9590/3
C0024299|T191|PT|C3208|NCI_CDISC|LYMPHOMA, MALIGNANT|9590/3
C0024299|T191|SY|C3208|NCI_CDISC|Malignant Lymphoma|9590/3
C0024299|T191|PT|C3208|NCI_CPTAC|Lymphoma|9590/3
C0024305|T191|PT|C3211|NCI_CPTAC|Non-Hodgkin Lymphoma|9590/3
C0024299|T191|PT|10025316|NCI_CTEP-SDC|Lymphoma, NOS|9590/3
C0024305|T191|SY|10029593|NCI_CTEP-SDC|NHL, NOS|9590/3
C0024305|T191|PT|10029593|NCI_CTEP-SDC|Non-Hodgkin lymphoma, NOS|9590/3
C0024299|T191|DN|C3208|NCI_CTRP|Lymphoma|9590/3
C0024299|T191|PT|C3208|NCI_CTRP|Lymphoma|9590/3
C0024305|T191|PT|C3211|NCI_CTRP|Non-Hodgkin Lymphoma|9590/3
C0024305|T191|DN|C3211|NCI_CTRP|Non-Hodgkin Lymphoma|9590/3
C0024299|T191|PT|3263|NCI_FDA|Lymphoma|9590/3
C0024299|T191|PT|CDR0000045368|NCI_NCI-GLOSS|lymphoma|9590/3
C0024305|T191|PT|CDR0000430869|NCI_NCI-GLOSS|NHL|9590/3
C0024305|T191|PT|CDR0000045148|NCI_NCI-GLOSS|non-Hodgkin lymphoma|9590/3
C0024299|T191|PT|C3208|NCI_NICHD|Lymphoma|9590/3
C0024305|T191|PT|C3211|NCI_NICHD|Non-Hodgkin Lymphoma|9590/3
C0024305|T191|SY|C3211|NCI_NICHD|Non-Hodgkin's Lymphoma|9590/3
C0024299|T191|PT|CDR0000041429|PDQ|lymphoma|9590/3
C0024305|T191|SY|CDR0000038957|PDQ|lymphoma, non-Hodgkin's|9590/3
C0024299|T191|SY|CDR0000041429|PDQ|malignant lymphoma|9590/3
C0024305|T191|AB|CDR0000038957|PDQ|NHL|9590/3
C0024305|T191|PT|CDR0000038957|PDQ|non-Hodgkin lymphoma|9590/3
C0024305|T191|SY|CDR0000038957|PDQ|Non-Hodgkin's Lymphoma|9590/3
C0024305|T191|PT|R0121804|QMR|MALIGNANT LYMPHOMA NON HODGKINS TYPE|9590/3
C0024299|T191|PT|X77q5|RCD|Lymphoma morphology|9590/3
C0024305|T191|AB|B627.|RCD|Malig lymphoma, non-Hodgkin's|9590/3
C0024299|T191|OA|B62y0|RCD|Malig.lymphoma NOS-unspec site|9590/3
C0024299|T191|PT|Xa99k|RCD|Malignant lymphoma|9590/3
C0024299|T191|OP|B62y.|RCD|Malignant lymphoma NOS|9590/3
C0024299|T191|OP|B62y0|RCD|Malignant lymphoma NOS of unspecified site|9590/3
C0024305|T191|SY|B627.|RCD|Malignant lymphoma, non-Hodgkin's type|9590/3
C0024305|T191|SY|B627.|RCD|NHL - Non-Hodgkin's lymphoma|9590/3
C0024305|T191|PT|B627.|RCD|Non-Hodgkin's lymphoma|9590/3
C0024305|T191|IS|XE2t9|RCD|Non-Hodgkin's lymphoma NOS|9590/3
C0024299|T191|IS|BBg1.|RCDSY|Lymphoma NOS|9590/3
C0024305|T191|OA|BBg2.|RCDSY|Mal lymphoma, non-Hodg type|9590/3
C0024305|T191|OA|BBgM.|RCDSY|Malg lymph,smal cleav,difus|9590/3
C0024299|T191|OP|BBg1.|RCDSY|Malignant lymphoma NOS|9590/3
C0024305|T191|OP|BBg2.|RCDSY|Malignant lymphoma, non-Hodgkin's type|9590/3
C0024305|T191|OP|BBgM.|RCDSY|Malignant lymphoma, small cleaved cell, diffuse|9590/3
C0024305|T191|OA|XE2t9|RCDSY|Non-Hod lympha, unspec type|9590/3
C0024305|T191|IS|BBg2.|RCDSY|Non-Hodgkin's lymphoma|9590/3
C0024305|T191|OP|XE2t9|RCDSY|Non-Hodgkin's lymphoma, unspecified type|9590/3
C0024299|T191|SY|118600007|SNOMEDCT_US|Lymphoma|9590/3
C0024299|T191|SY|21964009|SNOMEDCT_US|Lymphoma|9590/3
C0024299|T191|OAS|269627002|SNOMEDCT_US|Lymphoma|9590/3
C0024299|T191|OAP|134218000|SNOMEDCT_US|Lymphoma morphology|9590/3
C0024299|T191|IS|21964009|SNOMEDCT_US|Lymphoma, NOS|9590/3
C0024299|T191|PT|118600007|SNOMEDCT_US|Malignant lymphoma|9590/3
C0024299|T191|PT|21964009|SNOMEDCT_US|Malignant lymphoma|9590/3
C0024299|T191|PT|115244002|SNOMEDCT_US|Malignant lymphoma - category|9590/3
C0024299|T191|OF|188704004|SNOMEDCT_US|Malignant lymphoma NOS|9590/3
C0024299|T191|OAP|188694002|SNOMEDCT_US|Malignant lymphoma NOS|9590/3
C0024299|T191|OAP|188704004|SNOMEDCT_US|Malignant lymphoma NOS|9590/3
C0024299|T191|OAP|188695001|SNOMEDCT_US|Malignant lymphoma NOS of unspecified site|9590/3
C0024299|T191|SY|21964009|SNOMEDCT_US|Malignant lymphoma, no ICD-O subtype|9590/3
C0024299|T191|SY|21964009|SNOMEDCT_US|Malignant lymphoma, no International Classification of Diseases for Oncology subtype|9590/3
C0024305|T191|PT|1929004|SNOMEDCT_US|Malignant lymphoma, non-Hodgkin|9590/3
C0024305|T191|SY|1929004|SNOMEDCT_US|Malignant lymphoma, non-Hodgkin's|9590/3
C0024305|T191|SY|118601006|SNOMEDCT_US|Malignant lymphoma, non-Hodgkin's type|9590/3
C0024305|T191|IS|1929004|SNOMEDCT_US|Malignant lymphoma, non-Hodgkin's, NOS|9590/3
C0024299|T191|IS|21964009|SNOMEDCT_US|Malignant lymphoma, NOS|9590/3
C0024305|T191|IS|63086004|SNOMEDCT_US|Malignant lymphoma, small cleaved cell, diffuse -RETIRED-|9590/3
C0024305|T191|OF|63086004|SNOMEDCT_US|Malignant lymphoma, small cleaved cell, diffuse -RETIRED-|9590/3
C0024305|T191|SY|118601006|SNOMEDCT_US|NHL - Non-Hodgkin's lymphoma|9590/3
C0024305|T191|SY|118601006|SNOMEDCT_US|Non-Hodgkin lymphoma|9590/3
C0024305|T191|SY|128929007|SNOMEDCT_US|Non-Hodgkin lymphoma - category|9590/3
C0024305|T191|SY|1929004|SNOMEDCT_US|Non-Hodgkin lymphoma, no ICD-O subtype|9590/3
C0024305|T191|SY|1929004|SNOMEDCT_US|Non-Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype|9590/3
C0024305|T191|OAS|154583006|SNOMEDCT_US|Non-Hodgkin's lymphoma|9590/3
C0024305|T191|OAS|269628007|SNOMEDCT_US|Non-Hodgkin's lymphoma|9590/3
C0024305|T191|SY|118601006|SNOMEDCT_US|Non-Hodgkin's lymphoma|9590/3
C0024305|T191|SY|1929004|SNOMEDCT_US|Non-Hodgkin's lymphoma|9590/3
C0024305|T191|SY|118601006|SNOMEDCT_US|Non-Hodgkin's lymphoma - disorder|9590/3
C0024305|T191|OAS|271385002|SNOMEDCT_US|Non-Hodgkin's lymphoma NOS|9590/3
C0024305|T191|IS|1929004|SNOMEDCT_US|Non-Hodgkin's lymphoma, NOS|9590/3
C0024299|T191|SY|188676008|SNOMEDCT_US|Reticulolymphosarcoma|9590/3
C0024299|T191|PT|1110|WHO|LYMPHOMA MALIGNANT|9590/3
C0024305|T191|PT|1544|WHO|NON-HODGKIN'S LYMPHOMA|9590/3
C1266190|T191|LLT|10071541|MDR|Metastatic lymphoma|9590/6
C1266190|T191|PT|10071541|MDR|Metastatic lymphoma|9590/6
C1266190|T191|SY|110459008|SNOMEDCT_US|Lymphoma, metastatic|9590/6
C1266190|T191|PT|110459008|SNOMEDCT_US|Malignant lymphoma, metastatic|9590/6
C0024302|T191|ET|0000004626|AOD|histiocytic lymphoma|9591/3
C0024305|T191|AB|BI00323|BI|nhl|9591/3
C0024305|T191|PT|BI00323|BI|non-hodgkin's lymphoma|9591/3
C0024302|T191|PT|0047637|CCPSS|LYMPHOMA LARGE CELL|9591/3
C0024305|T191|PT|0001640|CCPSS|LYMPHOMA NON HODGKIN|9591/3
C0024305|T191|SD|38|CCS|Non-Hodgkin`s lymphoma|9591/3
C0024305|T191|MD|2.10.2|CCS|Non-Hodgkins lymphoma|9591/3
C0024305|T191|SD|NEO058|CCSR_10|Non-Hodgkin lymphoma|9591/3
C0024302|T191|SY|0000007619|CHV|cell large lymphomas|9591/3
C0024302|T191|SY|0000007619|CHV|cell reticulum sarcomas|9591/3
C0431132|T191|SY|0000034150|CHV|cells lymphoma stem|9591/3
C0024302|T191|SY|0000007619|CHV|cells reticulum sarcoma|9591/3
C0349633|T191|SY|0000007335|CHV|hairy cell leukaemia variant|9591/3
C0349633|T191|SY|0000007335|CHV|hairy cell leukemia variant|9591/3
C0024302|T191|SY|0000007619|CHV|histiocytic lymphoma|9591/3
C0024302|T191|PT|0000007619|CHV|large cell lymphoma|9591/3
C0024302|T191|SY|0000007619|CHV|lymphoma large cell|9591/3
C0431132|T191|SY|0000034150|CHV|lymphoma stem cell|9591/3
C0024305|T191|SY|0000007621|CHV|nhl|9591/3
C0024305|T191|SY|0000007621|CHV|non hodgkin lymphoma|9591/3
C0024305|T191|SY|0000007621|CHV|non hodgkin's lymphoma|9591/3
C0024305|T191|SY|0000007621|CHV|non hodgkins lymphoma|9591/3
C0024305|T191|SY|0000007621|CHV|non-hodgkin lymphoma|9591/3
C0024305|T191|SY|0000007621|CHV|non-hodgkin's lymphoma|9591/3
C0024305|T191|SY|0000007621|CHV|non-hodgkins lymphoma|9591/3
C0024305|T191|SY|0000007621|CHV|nonhodgkin lymphoma|9591/3
C0024305|T191|SY|0000007621|CHV|nonhodgkin's lymphoma|9591/3
C0024305|T191|SY|0000007621|CHV|nonhodgkins lymphoma|9591/3
C0024302|T191|SY|0000007619|CHV|reticulosarcoma|9591/3
C0024302|T191|SY|0000007619|CHV|reticulum cell sarcoma|9591/3
C0431132|T191|PT|0000034150|CHV|stem cell lymphoma|9591/3
C0024305|T191|PT|U000045|COSTAR|NON HODGKINS LYMPHOMA|9591/3
C0024305|T191|PT|525|COSTAR|NONHODGKINS LYMPHOMA|9591/3
C0024302|T191|PT|NOCODE|COSTAR|Reticulum Cell Sarcoma|9591/3
C0024302|T191|PT|2004-7036|CSP|histiocytic lymphoma|9591/3
C0024305|T191|PT|4001-0094|CSP|nonHodgkin's lymphoma|9591/3
C0024305|T191|SY|NOCODE|DXP|LYMPHOMA, NON HODGKIN|9591/3
C0024305|T191|SY|NOCODE|DXP|NHL|9591/3
C0024305|T191|FI|U002830|DXP|NON-HODGKIN LYMPHOMA|9591/3
C0024305|T191|PT|HP:0012539|HPO|Non-Hodgkin lymphoma|9591/3
C0024305|T191|PT|C85.9|ICD10|Non-Hodgkin's lymphoma, unspecified type|9591/3
C0024305|T191|ET|C85.9|ICD10CM|Non-Hodgkin lymphoma NOS|9591/3
C0024302|T191|HT|200.7|ICD9CM|Large cell lymphoma|9591/3
C0024302|T191|HT|200.0|ICD9CM|Reticulosarcoma|9591/3
C0024305|T191|PT|MTHU023065|ICPC2ICD10ENG|diffuse; lymphoma, small cell, cleaved|9591/3
C0024302|T191|PT|MTHU023078|ICPC2ICD10ENG|diffuse; reticulosarcoma|9591/3
C0024302|T191|PT|MTHU035166|ICPC2ICD10ENG|histiocytic; lymphoma|9591/3
C0024305|T191|PT|MTHU046759|ICPC2ICD10ENG|lymphoma; diffuse, small cell, cleaved|9591/3
C0024302|T191|PT|MTHU046800|ICPC2ICD10ENG|lymphoma; histiocytic|9591/3
C0024305|T191|PT|MTHU046842|ICPC2ICD10ENG|lymphoma; non-Hodgkin's|9591/3
C0024305|T191|PT|MTHU053464|ICPC2ICD10ENG|non-Hodgkin's lymphoma|9591/3
C0024305|T191|PT|MTHU053462|ICPC2ICD10ENG|non-Hodgkin's; lymphoma|9591/3
C0431136|T191|PT|MTHU060032|ICPC2ICD10ENG|pleomorphic cell type; reticulosarcoma|9591/3
C0024302|T191|PT|MTHU064360|ICPC2ICD10ENG|reticulosarcoma|9591/3
C0024302|T191|PT|MTHU064361|ICPC2ICD10ENG|reticulosarcoma; diffuse|9591/3
C0431136|T191|PT|MTHU064362|ICPC2ICD10ENG|reticulosarcoma; pleomorphic cell type|9591/3
C0024302|T191|PT|MTHU064376|ICPC2ICD10ENG|reticulum cell sarcoma|9591/3
C0024302|T191|PT|MTHU064373|ICPC2ICD10ENG|reticulum cell; sarcoma|9591/3
C0431136|T191|PT|MTHU064375|ICPC2ICD10ENG|reticulum cell; sarcoma, pleomorphic cell type|9591/3
C0024302|T191|PT|MTHU065928|ICPC2ICD10ENG|sarcoma; reticulum cell|9591/3
C0431136|T191|PT|MTHU065930|ICPC2ICD10ENG|sarcoma; reticulum cell, pleomorphic cell type|9591/3
C0024305|T191|PT|B74002|ICPC2P|Lymphoma;non Hodgkins|9591/3
C0024305|T191|PTN|B74002|ICPC2P|non hodgkins lymphoma|9591/3
C0024302|T191|PT|B74009|ICPC2P|Reticulosarcoma|9591/3
C0024302|T191|PTN|B74009|ICPC2P|reticulosarcoma|9591/3
C0024302|T191|PT|sh85113321|LCH_NW|Reticulum cell sarcoma|9591/3
C0349633|T191|LLT|10019054|MDR|Hairy cell leukaemia variant|9591/3
C0349633|T191|LLT|10019056|MDR|Hairy cell leukemia variant|9591/3
C4524190|T191|LLT|10080217|MDR|High-grade B-cell lymphoma, with MYC and BCL2 and/or BCL6 rearrangements|9591/3
C0024305|T191|PT|10029547|MDR|Non-Hodgkin's lymphoma|9591/3
C0024305|T191|LLT|10029547|MDR|Non-Hodgkin's lymphoma|9591/3
C0024305|T191|LLT|10029593|MDR|Non-Hodgkin's lymphoma NOS|9591/3
C0024302|T191|LLT|10038804|MDR|Reticulosarcoma|9591/3
C0349633|T191|PT|350013|MEDCIN|hairy-cell leukemia variant|9591/3
C0024302|T191|PT|312620|MEDCIN|large cell lymphoma|9591/3
C0349633|T191|SY|350013|MEDCIN|leukemia hairy-cell - variant|9591/3
C0024305|T191|PT|35839|MEDCIN|non-Hodgkin's lymphoma|9591/3
C0024302|T191|PT|92518|MEDCIN|reticulosarcoma|9591/3
C0024305|T191|SY|117|MEDLINEPLUS|Non-Hodgkin lymphoma|9591/3
C0024305|T191|ET|117|MEDLINEPLUS|Non-Hodgkin Lymphoma|9591/3
C0024305|T191|PM|D008228|MSH|Diffuse Small Cleaved Cell Lymphoma|9591/3
C0024305|T191|DEV|D008228|MSH|DIFFUSE SMALL CLEAVED LYMPHOMA|9591/3
C0024305|T191|ET|D008228|MSH|Diffuse Small Cleaved-Cell Lymphoma|9591/3
C0024305|T191|DEV|D008228|MSH|LYMPHOMA SMALL CLEAVED DIFFUSE|9591/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Atypical Diffuse Small Lymphoid|9591/3
C0024305|T191|PM|D008228|MSH|Lymphoma, Non Hodgkin|9591/3
C0024305|T191|PM|D008228|MSH|Lymphoma, Non Hodgkin's|9591/3
C0024305|T191|PM|D008228|MSH|Lymphoma, Non Hodgkins|9591/3
C0024305|T191|MH|D008228|MSH|Lymphoma, Non-Hodgkin|9591/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Non-Hodgkin's|9591/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Non-Hodgkins|9591/3
C0024305|T191|PM|D008228|MSH|Lymphoma, Nonhodgkin|9591/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Nonhodgkin's|9591/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Nonhodgkins|9591/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Small Cleaved Cell, Diffuse|9591/3
C0024305|T191|ET|D008228|MSH|Lymphoma, Small Cleaved-Cell, Diffuse|9591/3
C0024305|T191|PM|D008228|MSH|Non Hodgkin Lymphoma|9591/3
C0024305|T191|PM|D008228|MSH|Non Hodgkin's Lymphoma|9591/3
C0024305|T191|ET|D008228|MSH|Non-Hodgkin Lymphoma|9591/3
C0024305|T191|ET|D008228|MSH|Non-Hodgkin's Lymphoma|9591/3
C0024305|T191|PM|D008228|MSH|Non-Hodgkins Lymphoma|9591/3
C0024305|T191|DSV|D008228|MSH|NONHODGKIN LYMPHOMA|9591/3
C0024305|T191|PM|D008228|MSH|Nonhodgkin's Lymphoma|9591/3
C0024305|T191|PM|D008228|MSH|Nonhodgkins Lymphoma|9591/3
C0024302|T191|ET|D008228|MSH|Reticulosarcoma|9591/3
C0024302|T191|PM|D008228|MSH|Reticulosarcomas|9591/3
C0024302|T191|ET|D008228|MSH|Reticulum Cell Sarcoma|9591/3
C0024302|T191|PM|D008228|MSH|Reticulum Cell Sarcomas|9591/3
C0024302|T191|PEP|D008228|MSH|Reticulum-Cell Sarcoma|9591/3
C0024302|T191|PM|D008228|MSH|Reticulum-Cell Sarcomas|9591/3
C0024302|T191|PM|D008228|MSH|Sarcoma, Reticulum Cell|9591/3
C0024302|T191|ET|D008228|MSH|Sarcoma, Reticulum-Cell|9591/3
C0024305|T191|PM|D008228|MSH|Small Cleaved Cell Lymphoma, Diffuse|9591/3
C0024305|T191|DEV|D008228|MSH|SMALL CLEAVED LYMPHOMA DIFFUSE|9591/3
C0024305|T191|ET|D008228|MSH|Small Cleaved-Cell Lymphoma, Diffuse|9591/3
C0024305|T191|PN|NOCODE|MTH|Lymphoma, Non-Hodgkin|9591/3
C0024302|T191|PN|NOCODE|MTH|Reticulosarcoma|9591/3
C0431136|T191|ET|200.0|MTHICD9|Malignant lymphoma histiocytic pleomorphic cell type|9591/3
C0024302|T191|ET|200.0|MTHICD9|Malignant lymphoma reticulum cell type|9591/3
C0431136|T191|ET|200.0|MTHICD9|Pleomorphic cell type reticulum cell sarcoma|9591/3
C0024302|T191|ET|200.0|MTHICD9|Reticulum cell sarcoma NOS|9591/3
C0349633|T191|PT|C7401|NCI|Hairy Cell Leukemia Variant|9591/3
C0349633|T191|AB|C7401|NCI|HCL-V|9591/3
C4524190|T191|SY|C138195|NCI|HGBL with MYC and BCL2 and/or BCL6 Rearrangements|9591/3
C4524190|T191|PT|C138195|NCI|High Grade B-Cell Lymphoma with MYC and BCL2 and/or BCL6 Rearrangements|9591/3
C4524676|T191|PT|C133494|NCI|Large B-Cell Lymphoma with IRF4 Rearrangement|9591/3
C4524676|T191|SY|C133494|NCI|LBCL with IRF4 Rearrangement|9591/3
C0024305|T191|AB|C3211|NCI|NHL|9591/3
C0024305|T191|PT|C3211|NCI|Non-Hodgkin Lymphoma|9591/3
C0024305|T191|SY|C3211|NCI|Non-Hodgkin's Lymphoma|9591/3
C0349633|T191|SY|C7401|NCI|Prolymphocytic Variant of Hairy Cell Leukemia|9591/3
C0024302|T191|PT|C27824|NCI|Reticulosarcoma|9591/3
C0024302|T191|OP|C27824|NCI|Reticulosarcoma|9591/3
C2699507|T191|PT|C80308|NCI|Splenic B-Cell Lymphoma/Leukemia, Unclassifiable|9591/3
C2699508|T191|PT|C80309|NCI|Splenic Diffuse Red Pulp Small B-Cell Lymphoma|9591/3
C0024305|T191|PT|C3211|NCI_CPTAC|Non-Hodgkin Lymphoma|9591/3
C0024305|T191|SY|10029593|NCI_CTEP-SDC|NHL, NOS|9591/3
C0024305|T191|PT|10029593|NCI_CTEP-SDC|Non-Hodgkin lymphoma, NOS|9591/3
C4524190|T191|DN|C138195|NCI_CTRP|High Grade B-Cell Lymphoma with MYC and BCL2 and/or BCL6 Rearrangements|9591/3
C4524676|T191|DN|C133494|NCI_CTRP|Large B-Cell Lymphoma with IRF4 Rearrangement|9591/3
C0024305|T191|DN|C3211|NCI_CTRP|Non-Hodgkin Lymphoma|9591/3
C0024305|T191|PT|C3211|NCI_CTRP|Non-Hodgkin Lymphoma|9591/3
C0024305|T191|PT|CDR0000430869|NCI_NCI-GLOSS|NHL|9591/3
C0024305|T191|PT|CDR0000045148|NCI_NCI-GLOSS|non-Hodgkin lymphoma|9591/3
C0024305|T191|PT|C3211|NCI_NICHD|Non-Hodgkin Lymphoma|9591/3
C0024305|T191|SY|C3211|NCI_NICHD|Non-Hodgkin's Lymphoma|9591/3
C0024305|T191|SY|CDR0000038957|PDQ|lymphoma, non-Hodgkin's|9591/3
C0024305|T191|AB|CDR0000038957|PDQ|NHL|9591/3
C0024305|T191|PT|CDR0000038957|PDQ|non-Hodgkin lymphoma|9591/3
C0024305|T191|SY|CDR0000038957|PDQ|Non-Hodgkin's Lymphoma|9591/3
C0024305|T191|PT|R0121804|QMR|MALIGNANT LYMPHOMA NON HODGKINS TYPE|9591/3
C0349633|T191|PT|Xa0SA|RCD|Hairy cell leukaemia variant|9591/3
C0024305|T191|AB|B627.|RCD|Malig lymphoma, non-Hodgkin's|9591/3
C0431132|T191|OA|BBg4.|RCD|Malig lymphoma,stem cell type|9591/3
C0024305|T191|SY|B627.|RCD|Malignant lymphoma, non-Hodgkin's type|9591/3
C0431132|T191|OP|BBg4.|RCD|Malignant lymphoma, stem cell type|9591/3
C0024305|T191|SY|B627.|RCD|NHL - Non-Hodgkin's lymphoma|9591/3
C0024305|T191|PT|B627.|RCD|Non-Hodgkin's lymphoma|9591/3
C0024305|T191|IS|XE2t9|RCD|Non-Hodgkin's lymphoma NOS|9591/3
C0431136|T191|AB|BBh1.|RCD|Reticulosarc, pleomorph cell|9591/3
C0024302|T191|PT|B600.|RCD|Reticulosarcoma|9591/3
C0024302|T191|OA|B6000|RCD|Reticulosarcoma - unspec site|9591/3
C0024302|T191|PT|BBh..|RCD|Reticulosarcoma morphology|9591/3
C0024302|T191|OP|B600z|RCD|Reticulosarcoma NOS|9591/3
C0024302|T191|OP|B6000|RCD|Reticulosarcoma of unspecified site|9591/3
C0547066|T191|PT|BBh2.|RCD|Reticulosarcoma, nodular|9591/3
C0431136|T191|PT|BBh1.|RCD|Reticulosarcoma, pleomorphic cell type|9591/3
C0024302|T191|SY|B600.|RCD|Reticulum cell sarcoma|9591/3
C0024302|T191|SY|BBh..|RCD|Reticulum cell sarcoma morphol|9591/3
C0349633|T191|PT|Xa0SA|RCDAE|Hairy cell leukemia variant|9591/3
C0024302|T191|OP|BBmH.|RCDSY|Large cell lymphoma|9591/3
C0024305|T191|OA|BBg2.|RCDSY|Mal lymphoma, non-Hodg type|9591/3
C0024305|T191|OA|BBgM.|RCDSY|Malg lymph,smal cleav,difus|9591/3
C0024305|T191|OP|BBg2.|RCDSY|Malignant lymphoma, non-Hodgkin's type|9591/3
C0024305|T191|OP|BBgM.|RCDSY|Malignant lymphoma, small cleaved cell, diffuse|9591/3
C0024305|T191|OA|XE2t9|RCDSY|Non-Hod lympha, unspec type|9591/3
C0024305|T191|IS|BBg2.|RCDSY|Non-Hodgkin's lymphoma|9591/3
C0024305|T191|OP|XE2t9|RCDSY|Non-Hodgkin's lymphoma, unspecified type|9591/3
C0024302|T191|SY|BBh..|RCDSY|Reticulosarcoma NOS|9591/3
C1282448|T191|PT|314922006|SNOMEDCT_US|B-cell lymphoma morphology|9591/3
C1282460|T191|PT|314934003|SNOMEDCT_US|Diffuse high grade B-cell lymphoma morphology|9591/3
C0349633|T191|SYGB|54087003|SNOMEDCT_US|Hairy cell leukaemia variant|9591/3
C0349633|T191|PTGB|277568007|SNOMEDCT_US|Hairy cell leukaemia variant|9591/3
C0349633|T191|PT|277568007|SNOMEDCT_US|Hairy cell leukemia variant|9591/3
C0349633|T191|SY|54087003|SNOMEDCT_US|Hairy cell leukemia variant|9591/3
C1282451|T191|PT|314925008|SNOMEDCT_US|High grade B-cell lymphoma morphology|9591/3
C4524190|T191|PT|786909001|SNOMEDCT_US|High grade B-cell lymphoma with MYC and BCL2 and/or BCL6 rearrangements|9591/3
C0024302|T191|SY|715664005|SNOMEDCT_US|Interdigitating cell sarcoma|9591/3
C0024302|T191|PT|715664005|SNOMEDCT_US|Interdigitating dendritic cell sarcoma|9591/3
C4524676|T191|SY|786960000|SNOMEDCT_US|Large B-cell lymphoma with interferon regulatory factor 4 rearrangement|9591/3
C4524676|T191|PT|786960000|SNOMEDCT_US|Large B-cell lymphoma with IRF4 rearrangement|9591/3
C1282449|T191|PT|314923001|SNOMEDCT_US|Low grade B-cell lymphoma morphology|9591/3
C0024305|T191|PT|1929004|SNOMEDCT_US|Malignant lymphoma, non-Hodgkin|9591/3
C0024305|T191|SY|1929004|SNOMEDCT_US|Malignant lymphoma, non-Hodgkin's|9591/3
C0024305|T191|SY|118601006|SNOMEDCT_US|Malignant lymphoma, non-Hodgkin's type|9591/3
C0024305|T191|IS|1929004|SNOMEDCT_US|Malignant lymphoma, non-Hodgkin's, NOS|9591/3
C0024305|T191|OF|63086004|SNOMEDCT_US|Malignant lymphoma, small cleaved cell, diffuse -RETIRED-|9591/3
C0024305|T191|IS|63086004|SNOMEDCT_US|Malignant lymphoma, small cleaved cell, diffuse -RETIRED-|9591/3
C0431132|T191|PT|189962004|SNOMEDCT_US|Malignant lymphoma, stem cell type|9591/3
C0024305|T191|SY|118601006|SNOMEDCT_US|NHL - Non-Hodgkin's lymphoma|9591/3
C1282457|T191|PT|314931006|SNOMEDCT_US|Nodular high grade B-cell lymphoma morphology|9591/3
C0024305|T191|SY|118601006|SNOMEDCT_US|Non-Hodgkin lymphoma|9591/3
C0024305|T191|SY|128929007|SNOMEDCT_US|Non-Hodgkin lymphoma - category|9591/3
C0024305|T191|SY|1929004|SNOMEDCT_US|Non-Hodgkin lymphoma, no ICD-O subtype|9591/3
C0024305|T191|SY|1929004|SNOMEDCT_US|Non-Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype|9591/3
C0024305|T191|OAS|154583006|SNOMEDCT_US|Non-Hodgkin's lymphoma|9591/3
C0024305|T191|OAS|269628007|SNOMEDCT_US|Non-Hodgkin's lymphoma|9591/3
C0024305|T191|SY|118601006|SNOMEDCT_US|Non-Hodgkin's lymphoma|9591/3
C0024305|T191|SY|1929004|SNOMEDCT_US|Non-Hodgkin's lymphoma|9591/3
C0024305|T191|SY|118601006|SNOMEDCT_US|Non-Hodgkin's lymphoma - disorder|9591/3
C0024305|T191|OAS|271385002|SNOMEDCT_US|Non-Hodgkin's lymphoma NOS|9591/3
C0024305|T191|IS|1929004|SNOMEDCT_US|Non-Hodgkin's lymphoma, NOS|9591/3
C1688594|T191|PT|418265009|SNOMEDCT_US|Primary cutaneous B-cell lymphoma - category|9591/3
C0024302|T191|OAP|154579006|SNOMEDCT_US|Reticulosarcoma|9591/3
C0024302|T191|PT|373168002|SNOMEDCT_US|Reticulosarcoma|9591/3
C0024302|T191|OAP|40152000|SNOMEDCT_US|Reticulosarcoma|9591/3
C0024302|T191|OAP|118604003|SNOMEDCT_US|Reticulosarcoma|9591/3
C0024302|T191|OF|154579006|SNOMEDCT_US|Reticulosarcoma|9591/3
C0024302|T191|IS|40152000|SNOMEDCT_US|Reticulosarcoma -RETIRED-|9591/3
C0024302|T191|OF|40152000|SNOMEDCT_US|Reticulosarcoma -RETIRED-|9591/3
C0024302|T191|OAP|189983005|SNOMEDCT_US|Reticulosarcoma morphology|9591/3
C0024302|T191|OAP|189986002|SNOMEDCT_US|Reticulosarcoma morphology|9591/3
C0024302|T191|OF|189983005|SNOMEDCT_US|Reticulosarcoma morphology|9591/3
C0024302|T191|OF|189986002|SNOMEDCT_US|Reticulosarcoma morphology|9591/3
C0024302|T191|PT|189982000|SNOMEDCT_US|Reticulosarcoma morphology|9591/3
C0024302|T191|OAP|188497004|SNOMEDCT_US|Reticulosarcoma NOS|9591/3
C0024302|T191|OAP|188488003|SNOMEDCT_US|Reticulosarcoma of unspecified site|9591/3
C0024302|T191|IS|40152000|SNOMEDCT_US|Reticulosarcoma, diffuse|9591/3
C0547066|T191|PT|189985003|SNOMEDCT_US|Reticulosarcoma, nodular|9591/3
C0024302|T191|IS|40152000|SNOMEDCT_US|Reticulosarcoma, NOS|9591/3
C0431136|T191|PT|189984004|SNOMEDCT_US|Reticulosarcoma, pleomorphic cell type|9591/3
C0024302|T191|SY|715664005|SNOMEDCT_US|Reticulum cell sarcoma|9591/3
C0024302|T191|SY|373168002|SNOMEDCT_US|Reticulum cell sarcoma|9591/3
C0024302|T191|OAS|118604003|SNOMEDCT_US|Reticulum cell sarcoma|9591/3
C0024302|T191|IS|189982000|SNOMEDCT_US|Reticulum cell sarcoma morphol|9591/3
C0024302|T191|SY|189982000|SNOMEDCT_US|Reticulum cell sarcoma morphology|9591/3
C0024302|T191|IS|40152000|SNOMEDCT_US|Reticulum cell sarcoma, diffuse|9591/3
C0024302|T191|IS|40152000|SNOMEDCT_US|Reticulum cell sarcoma, NOS|9591/3
C4518419|T191|PT|734141009|SNOMEDCT_US|Splenic B-cell lymphoma|9591/3
C2699508|T191|PT|763884007|SNOMEDCT_US|Splenic diffuse red pulp small B-cell lymphoma|9591/3
C2699508|T191|PT|734067001|SNOMEDCT_US|Splenic diffuse red pulp small B-cell lymphoma|9591/3
C0024305|T191|PT|1544|WHO|NON-HODGKIN'S LYMPHOMA|9591/3
C0545080|T191|PT|10073957|MDR|Composite lymphoma|9596/3
C0545080|T191|LLT|10073957|MDR|Composite lymphoma|9596/3
C1333878|T191|PT|366686|MEDCIN|B-cell lymphoma unclassifiable with features intermediate between classical Hodgkin lymphoma and diffuse large B-cell lymphoma|9596/3
C0545080|T191|MH|D058617|MSH|Composite Lymphoma|9596/3
C0545080|T191|PM|D058617|MSH|Composite Lymphomas|9596/3
C0545080|T191|PM|D058617|MSH|Lymphoma, Composite|9596/3
C0545080|T191|PM|D058617|MSH|Lymphomas, Composite|9596/3
C1333878|T191|PT|C37869|NCI|B-Cell Lymphoma, Unclassifiable, with Features Intermediate between Diffuse Large B-Cell Lymphoma and Classic Hodgkin Lymphoma|9596/3
C1333878|T191|SY|C37869|NCI|B-Cell Lymphoma, Unclassifiable, with Features Intermediate between Diffuse Large B-Cell Lymphoma and Classical Hodgkin Lymphoma|9596/3
C0545080|T191|PT|C38661|NCI|Composite Lymphoma|9596/3
C1333878|T191|SY|C37869|NCI|Gray Zone Lymphoma|9596/3
C1333878|T191|SY|C37869|NCI|Hodgkin-Like Anaplastic Large Cell Lymphoma|9596/3
C1333878|T191|SY|C37869|NCI|Large B-Cell Lymphoma with Hodgkin Features|9596/3
C1333878|T191|PT|C37869|NCI_CPTAC|B-Cell Lymphoma, Unclassifiable, with Features Intermediate between Diffuse Large B-Cell Lymphoma and Classic Hodgkin Lymphoma|9596/3
C0545080|T191|PT|C38661|NCI_CPTAC|Composite Lymphoma|9596/3
C1333878|T191|DN|C37869|NCI_CTRP|B-Cell Lymphoma, Unclassifiable, with Features Intermediate between Diffuse Large B-Cell Lymphoma and Classic Hodgkin Lymphoma|9596/3
C0545080|T191|PT|C38661|NCI_CTRP|Composite Lymphoma|9596/3
C0545080|T191|DN|C38661|NCI_CTRP|Composite Lymphoma|9596/3
C0545080|T191|PT|CDR0000633086|NCI_NCI-GLOSS|composite lymphoma|9596/3
C1333878|T191|PT|722954005|SNOMEDCT_US|B-cell lymphoma unclassifiable with features intermediate between classical Hodgkin lymphoma and diffuse large B-cell lymphoma|9596/3
C4301998|T191|PT|12351000132102|SNOMEDCT_US|B-cell lymphoma, unclassifiable, with features intermediate between diffuse large B-cell lymphoma and Hodgkin lymphoma|9596/3
C1266191|T191|PT|128798004|SNOMEDCT_US|Composite Hodgkin and non-Hodgkin lymphoma|9596/3
C1333171|T191|SY|357441|MEDCIN|malignant neoplasm lymphoma b-cell primary cutaneous follicular center|9597/3
C1333171|T191|PT|357441|MEDCIN|Primary cutaneous follicular center B-cell lymphoma|9597/3
C1333171|T191|PN|NOCODE|MTH|Primary Cutaneous Follicle Center Lymphoma|9597/3
C1333171|T191|SY|C7217|NCI|Crosti's Disease|9597/3
C1333171|T191|SY|C7217|NCI|Cutaneous Follicle Center Lymphoma|9597/3
C1333171|T191|SY|C7217|NCI|Cutaneous Follicle Centre Lymphoma|9597/3
C1333171|T191|AB|C7217|NCI|PCFCL|9597/3
C1333171|T191|PT|C7217|NCI|Primary Cutaneous Follicle Center Lymphoma|9597/3
C1333171|T191|SY|C7217|NCI|Reticulohistiocytoma of the Dorsum|9597/3
C1333171|T191|SY|404143002|SNOMEDCT_US|Crosti's lymphoma|9597/3
C1333171|T191|PT|419662008|SNOMEDCT_US|Primary cutaneous follicle center cell lymphoma|9597/3
C1333171|T191|SY|419662008|SNOMEDCT_US|Primary cutaneous follicle center lymphoma|9597/3
C1333171|T191|SY|404143002|SNOMEDCT_US|Primary cutaneous follicle center lymphoma|9597/3
C1333171|T191|PTGB|419662008|SNOMEDCT_US|Primary cutaneous follicle centre cell lymphoma|9597/3
C1333171|T191|SYGB|419662008|SNOMEDCT_US|Primary cutaneous follicle centre lymphoma|9597/3
C1333171|T191|SYGB|404143002|SNOMEDCT_US|Primary cutaneous follicle centre lymphoma|9597/3
C1333171|T191|SYGB|404143002|SNOMEDCT_US|Primary cutaneous follicle centre-cell B-cell lymphoma|9597/3
C1333171|T191|PT|404143002|SNOMEDCT_US|Primary cutaneous follicular center B-cell lymphoma|9597/3
C1333171|T191|PTGB|404143002|SNOMEDCT_US|Primary cutaneous follicular centre B-cell lymphoma|9597/3
C1333171|T191|IS|404143002|SNOMEDCT_US|Reticulohistiocytome du dos de l'adulte|9597/3
C0019829|T191|ET|0000004628|AOD|Hodgkin's disease|9650/3
C0019829|T191|AB|BI00314|BI|hd|9650/3
C0019829|T191|PT|BI00314|BI|hodgkin's disease|9650/3
C0019829|T191|RT|BI00314|BI|hodgkin's lymphoma|9650/3
C0019829|T191|PT|1006070|CCPSS|LYMPHOMA HODGKIN|9650/3
C0019829|T191|SD|37|CCS|Hodgkin`s disease|9650/3
C0019829|T191|MD|2.10.1|CCS|Hodgkins disease|9650/3
C0019829|T191|SD|NEO057|CCSR_10|Hodgkin lymphoma|9650/3
C0019829|T191|SY|0000006210|CHV|HD|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkin disease|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkin lymphoma|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkin lymphomas|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkin's disease|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphoma|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphoma disease|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphomas|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkins disease|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkins diseases|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkins lymphoma|9650/3
C0019829|T191|SY|0000006210|CHV|hodgkins lymphomas|9650/3
C0019829|T191|SY|0000006210|CHV|lymphogranulomatosis|9650/3
C0019829|T191|PT|U000356|COSTAR|HODGKIN'S DISEASE|9650/3
C0019829|T191|PT|376|COSTAR|HODGKINS DISEASE|9650/3
C0019829|T191|PT|2004-1208|CSP|Hodgkin's disease|9650/3
C0019829|T191|ET|2004-1208|CSP|lymphogranulomatosis|9650/3
C0019829|T191|GT|LYMPHOMA LIKE REACT|CST|HODGINS|9650/3
C0019829|T191|DI|U000853|DXP|HODGKINS DISEASE|9650/3
C0019829|T191|SY|HP:0012189|HPO|Hodgkin disease|9650/3
C0019829|T191|PT|HP:0012189|HPO|Hodgkin lymphoma|9650/3
C0019829|T191|SY|HP:0012189|HPO|Hodgkin's lymphoma|9650/3
C0019829|T191|HT|C81|ICD10|Hodgkin's disease|9650/3
C0019829|T191|PT|C81.9|ICD10|Hodgkin's disease, unspecified|9650/3
C1333064|T191|ET|C81.7|ICD10CM|Classical Hodgkin lymphoma NOS|9650/3
C0019829|T191|AB|C81|ICD10CM|Hodgkin lymphoma|9650/3
C0019829|T191|HT|C81|ICD10CM|Hodgkin lymphoma|9650/3
C0019829|T191|AB|C81.9|ICD10CM|Hodgkin lymphoma, unspecified|9650/3
C0019829|T191|HT|C81.9|ICD10CM|Hodgkin lymphoma, unspecified|9650/3
C0019829|T191|HT|201|ICD9CM|Hodgkin's disease|9650/3
C0019829|T191|HT|201.9|ICD9CM|Hodgkin's disease, unspecified type|9650/3
C0019829|T191|HT|201.1|ICD9CM|Hodgkin's granuloma|9650/3
C0019829|T191|HT|201.0|ICD9CM|Hodgkin's paragranuloma|9650/3
C0019829|T191|HT|201.2|ICD9CM|Hodgkin's sarcoma|9650/3
C0019829|T191|PT|B72|ICPC|Hodgkins disease|9650/3
C0019829|T191|AB|B72|ICPC2EENG|Hodgkin's disease/lymphoma|9650/3
C0019829|T191|PT|B72|ICPC2EENG|Hodgkin's disease/lymphoma|9650/3
C0019829|T191|PT|MTHU083121|ICPC2ICD10ENG|disease; Hodgkin|9650/3
C0019829|T191|PT|MTHU032756|ICPC2ICD10ENG|granuloma; Hodgkin|9650/3
C0019829|T191|PT|MTHU032780|ICPC2ICD10ENG|granuloma; malignant|9650/3
C0019829|T191|PT|MTHU035331|ICPC2ICD10ENG|Hodgkin|9650/3
C0019829|T191|PT|MTHU035334|ICPC2ICD10ENG|Hodgkin; granuloma|9650/3
C0019829|T191|PT|MTHU035344|ICPC2ICD10ENG|Hodgkin; lymphoma|9650/3
C0019829|T191|PT|MTHU035351|ICPC2ICD10ENG|Hodgkin; paragranuloma|9650/3
C0019829|T191|PT|MTHU035352|ICPC2ICD10ENG|Hodgkin; sarcoma|9650/3
C0019829|T191|PT|MTHU046802|ICPC2ICD10ENG|lymphoma; Hodgkin|9650/3
C0019829|T191|PT|MTHU047288|ICPC2ICD10ENG|malignant; granuloma|9650/3
C0019829|T191|PT|MTHU057409|ICPC2ICD10ENG|paragranuloma; Hodgkin|9650/3
C0019829|T191|PT|MTHU065903|ICPC2ICD10ENG|sarcoma; Hodgkin|9650/3
C0019829|T191|PT|B72001|ICPC2P|Disease;Hodgkins|9650/3
C0019829|T191|PTN|B72001|ICPC2P|Hodgkins disease|9650/3
C0019829|T191|PTN|B72003|ICPC2P|hodgkins lymphoma|9650/3
C0019829|T191|PTN|B72004|ICPC2P|Hodgkins sarcoma|9650/3
C0019829|T191|PT|B72003|ICPC2P|Lymphoma;Hodgkins|9650/3
C0019829|T191|PT|B72004|ICPC2P|Sarcoma;Hodgkins|9650/3
C0019829|T191|PT|U002210|LCH|Hodgkin's disease|9650/3
C0019829|T191|PT|sh85061347|LCH_NW|Hodgkin's disease|9650/3
C0019829|T191|LA|LA26792-4|LNC|Hodgkin lymphoma|9650/3
C1333064|T191|LLT|10080208|MDR|Classical Hodgkin lymphoma|9650/3
C0019829|T191|OL|10020205|MDR|Hodgins|9650/3
C0019829|T191|PT|10020206|MDR|Hodgkin's disease|9650/3
C0019829|T191|LLT|10020206|MDR|Hodgkin's disease|9650/3
C0019829|T191|LLT|10020255|MDR|Hodgkin's disease NOS|9650/3
C0019829|T191|LLT|10020309|MDR|Hodgkin's disease, unspecified type|9650/3
C0019829|T191|LLT|10020318|MDR|Hodgkin's granuloma|9650/3
C0019829|T191|LLT|10020328|MDR|Hodgkin's lymphoma|9650/3
C0019829|T191|LLT|10020329|MDR|Hodgkin's paragranuloma|9650/3
C0019829|T191|LLT|10020339|MDR|Hodgkin's sarcoma|9650/3
C0019829|T191|LLT|10063666|MDR|Lymphogranulomatosis|9650/3
C0019829|T191|HG|10025319|MDR|Lymphomas Hodgkin's disease|9650/3
C0019829|T191|PT|31691|MEDCIN|Hodgkin disease|9650/3
C0019829|T191|PT|92514|MEDCIN|Hodgkin disease granuloma|9650/3
C0019829|T191|PT|92513|MEDCIN|Hodgkin disease paragranuloma|9650/3
C0019829|T191|PT|92515|MEDCIN|Hodgkin disease sarcoma|9650/3
C0019829|T191|PT|1262|MEDLINEPLUS|Hodgkin Disease|9650/3
C0019829|T191|SY|1262|MEDLINEPLUS|Hodgkin lymphoma|9650/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkin|9650/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkin's|9650/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkins|9650/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkin|9650/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkin's|9650/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkins|9650/3
C0019829|T191|ET|D006689|MSH|Granuloma, Malignant|9650/3
C0019829|T191|DEV|D006689|MSH|HODGKIN DIS|9650/3
C0019829|T191|MH|D006689|MSH|Hodgkin Disease|9650/3
C0019829|T191|PM|D006689|MSH|Hodgkin Granuloma|9650/3
C0019829|T191|ET|D006689|MSH|Hodgkin Lymphoma|9650/3
C0019829|T191|ET|D006689|MSH|Hodgkin's Disease|9650/3
C0019829|T191|PM|D006689|MSH|Hodgkin's Granuloma|9650/3
C0019829|T191|ET|D006689|MSH|Hodgkin's Lymphoma|9650/3
C0019829|T191|DEV|D006689|MSH|HODGKINS DIS|9650/3
C0019829|T191|ET|D006689|MSH|Hodgkins Disease|9650/3
C0019829|T191|PM|D006689|MSH|Hodgkins Granuloma|9650/3
C0019829|T191|PM|D006689|MSH|Hodgkins Lymphoma|9650/3
C0019829|T191|ET|D006689|MSH|Lymphogranuloma, Malignant|9650/3
C0019829|T191|PM|D006689|MSH|Lymphogranulomas, Malignant|9650/3
C0019829|T191|PM|D006689|MSH|Lymphoma, Hodgkin|9650/3
C0019829|T191|PM|D006689|MSH|Lymphoma, Hodgkin's|9650/3
C0019829|T191|PM|D006689|MSH|Malignant Granuloma|9650/3
C0019829|T191|PM|D006689|MSH|Malignant Granulomas|9650/3
C0019829|T191|PM|D006689|MSH|Malignant Lymphogranuloma|9650/3
C0019829|T191|PM|D006689|MSH|Malignant Lymphogranulomas|9650/3
C1333064|T191|PN|NOCODE|MTH|Classical Hodgkin's Lymphoma|9650/3
C0019829|T191|PN|NOCODE|MTH|Hodgkin Disease|9650/3
C0019829|T191|PT|376|MTH|Hodgkin's Disease|9650/3
C0019829|T191|ET|201.9|MTHICD9|Hodgkin's disease NOS|9650/3
C0019829|T191|ET|201.9|MTHICD9|Hodgkin's lymphoma NOS|9650/3
C0019829|T191|ET|201.9|MTHICD9|Malignant lymphogranuloma|9650/3
C0019829|T191|ET|201.9|MTHICD9|Malignant lymphogranulomatosis|9650/3
C1333064|T191|AB|C7164|NCI|cHL|9650/3
C1333064|T191|PT|C7164|NCI|Classic Hodgkin Lymphoma|9650/3
C1333064|T191|SY|C7164|NCI|Classical Hodgkin Lymphoma|9650/3
C1333064|T191|SY|C7164|NCI|Classical Hodgkin's Lymphoma|9650/3
C0019829|T191|AB|C9357|NCI|HL|9650/3
C0019829|T191|PT|C9357|NCI|Hodgkin Lymphoma|9650/3
C0019829|T191|SY|C9357|NCI|Hodgkin's Disease|9650/3
C0019829|T191|PT|C6914|NCI|Hodgkin's Granuloma|9650/3
C0019829|T191|OP|C6914|NCI|Hodgkin's Granuloma|9650/3
C0019829|T191|SY|C9357|NCI|Hodgkin's Lymphoma|9650/3
C0019829|T191|PT|C26956|NCI|Hodgkin's Paragranuloma|9650/3
C0019829|T191|OP|C26956|NCI|Hodgkin's Paragranuloma|9650/3
C1333064|T191|PT|C7164|NCI_CPTAC|Classic Hodgkin Lymphoma|9650/3
C0019829|T191|PT|C9357|NCI_CPTAC|Hodgkin Lymphoma|9650/3
C0019829|T191|SY|C9357|NCI_CPTAC|Hodgkin's Disease|9650/3
C0019829|T191|PT|C26956|NCI_CPTAC|Hodgkins Paragranuloma|9650/3
C0019829|T191|PT|10020255|NCI_CTEP-SDC|Hodgkin lymphoma, NOS|9650/3
C1333064|T191|DN|C7164|NCI_CTRP|Classical Hodgkin Lymphoma|9650/3
C0019829|T191|DN|C9357|NCI_CTRP|Hodgkin Lymphoma|9650/3
C0019829|T191|PT|C9357|NCI_CTRP|Hodgkin Lymphoma|9650/3
C1333064|T191|PT|CDR0000574284|NCI_NCI-GLOSS|classical Hodgkin lymphoma|9650/3
C0019829|T191|PT|CDR0000045012|NCI_NCI-GLOSS|Hodgkin disease|9650/3
C0019829|T191|PT|CDR0000270800|NCI_NCI-GLOSS|Hodgkin lymphoma|9650/3
C0019829|T191|PT|C9357|NCI_NICHD|Hodgkin Lymphoma|9650/3
C0019829|T191|SY|C9357|NCI_NICHD|Hodgkin's Disease|9650/3
C0019829|T191|SY|C9357|NCI_NICHD|Hodgkin's Lymphoma|9650/3
C0019829|T191|AB|CDR0000041646|PDQ|HL|9650/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkin disease|9650/3
C0019829|T191|PT|CDR0000041646|PDQ|Hodgkin lymphoma|9650/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkin's disease|9650/3
C0019829|T191|LV|CDR0000041646|PDQ|Hodgkin's lymphoma|9650/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkins disease|9650/3
C0019829|T191|LV|CDR0000041646|PDQ|Hodgkins lymphoma|9650/3
C0019829|T191|PT|R0121435|QMR|HODGKINS DISEASE SYSTEMIC|9650/3
C0019829|T191|SY|B61..|RCD|HD - Hodgkin's disease|9650/3
C0019829|T191|OA|B61z0|RCD|Hodgkin's dis.NOS-unspec. site|9650/3
C0019829|T191|PT|B61..|RCD|Hodgkin's disease|9650/3
C0019829|T191|OP|B61z.|RCD|Hodgkin's disease NOS|9650/3
C0019829|T191|OP|B61z0|RCD|Hodgkin's disease NOS, unspecified site|9650/3
C0019829|T191|PT|B611.|RCD|Hodgkin's granuloma|9650/3
C0019829|T191|OP|B611z|RCD|Hodgkin's granuloma NOS|9650/3
C0019829|T191|OP|B6110|RCD|Hodgkin's granuloma of unspecified site|9650/3
C0019829|T191|OA|B6110|RCD|Hodgkin's granuloma-unsp. site|9650/3
C0019829|T191|OA|B6100|RCD|Hodgkin's paragran-unspec site|9650/3
C0019829|T191|PT|B610.|RCD|Hodgkin's paragranuloma|9650/3
C0019829|T191|OP|B610z|RCD|Hodgkin's paragranuloma NOS|9650/3
C0019829|T191|OP|B6100|RCD|Hodgkin's paragranuloma of unspecified site|9650/3
C0019829|T191|PT|B612.|RCD|Hodgkin's sarcoma|9650/3
C0019829|T191|OP|B612z|RCD|Hodgkin's sarcoma NOS|9650/3
C0019829|T191|OP|B6120|RCD|Hodgkin's sarcoma of unspecified site|9650/3
C0019829|T191|OA|B6120|RCD|Hodgkin's sarcoma-unspec. site|9650/3
C0019829|T191|SY|B61..|RCD|Malignant Hodgkin's lymphoma|9650/3
C0019829|T191|PT|BBj..|RCDSY|Hodgkin's disease|9650/3
C0019829|T191|OP|XaC2n|RCDSY|Hodgkin's disease NOS|9650/3
C0019829|T191|OP|BBj9.|RCDSY|Hodgkin's granuloma|9650/3
C0019829|T191|OP|BBj8.|RCDSY|Hodgkin's paragranuloma|9650/3
C0019829|T191|OP|BBjA.|RCDSY|Hodgkin's sarcoma|9650/3
C0019829|T191|OP|XE1we|RCDSY|Lymphogranuloma, malignant|9650/3
C1333064|T191|PT|762690000|SNOMEDCT_US|Classical Hodgkin lymphoma|9650/3
C1333064|T191|PT|762691001|SNOMEDCT_US|Classical Hodgkin lymphoma|9650/3
C0019829|T191|SY|118599009|SNOMEDCT_US|HD - Hodgkin's disease|9650/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Hodgkin disease|9650/3
C0019829|T191|SY|118602004|SNOMEDCT_US|Hodgkin granuloma|9650/3
C0019829|T191|PT|14537002|SNOMEDCT_US|Hodgkin lymphoma|9650/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin lymphoma, no ICD-O subtype|9650/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype|9650/3
C0019829|T191|SY|118606001|SNOMEDCT_US|Hodgkin sarcoma|9650/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Hodgkin's disease|9650/3
C0019829|T191|OAP|154582001|SNOMEDCT_US|Hodgkin's disease|9650/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin's disease|9650/3
C0019829|T191|OF|154582001|SNOMEDCT_US|Hodgkin's disease|9650/3
C0019829|T191|OAP|188595005|SNOMEDCT_US|Hodgkin's disease NOS|9650/3
C0019829|T191|OAP|188605006|SNOMEDCT_US|Hodgkin's disease NOS|9650/3
C0019829|T191|OF|188605006|SNOMEDCT_US|Hodgkin's disease NOS|9650/3
C0019829|T191|OAP|188596006|SNOMEDCT_US|Hodgkin's disease NOS, unspecified site|9650/3
C0019829|T191|IS|14537002|SNOMEDCT_US|Hodgkin's disease, NOS|9650/3
C0019829|T191|SY|118602004|SNOMEDCT_US|Hodgkin's granuloma|9650/3
C0019829|T191|SY|74189002|SNOMEDCT_US|Hodgkin's granuloma|9650/3
C0019829|T191|OAP|188542007|SNOMEDCT_US|Hodgkin's granuloma NOS|9650/3
C0019829|T191|OAP|188533000|SNOMEDCT_US|Hodgkin's granuloma of unspecified site|9650/3
C0019829|T191|OAP|52337003|SNOMEDCT_US|Hodgkin's paragranuloma|9650/3
C0019829|T191|OAP|188521005|SNOMEDCT_US|Hodgkin's paragranuloma|9650/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma -RETIRED-|9650/3
C0019829|T191|OF|52337003|SNOMEDCT_US|Hodgkin's paragranuloma -RETIRED-|9650/3
C0019829|T191|OAP|188532005|SNOMEDCT_US|Hodgkin's paragranuloma NOS|9650/3
C0019829|T191|OAP|188522003|SNOMEDCT_US|Hodgkin's paragranuloma of unspecified site|9650/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma, nodular|9650/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma, NOS|9650/3
C0019829|T191|SY|118606001|SNOMEDCT_US|Hodgkin's sarcoma|9650/3
C0019829|T191|SY|46923007|SNOMEDCT_US|Hodgkin's sarcoma|9650/3
C0019829|T191|OAP|188552006|SNOMEDCT_US|Hodgkin's sarcoma NOS|9650/3
C0019829|T191|OAP|188543002|SNOMEDCT_US|Hodgkin's sarcoma of unspecified site|9650/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Lymphoma, Hodgkins|9650/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Malignant Hodgkin's lymphoma|9650/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Malignant lymphoma, Hodgkin's|9650/3
C1266194|T191|PX|C81.0|ICD10|Hodgkin's disease with lymphocytic predominance|9651/3
C1266194|T191|PS|C81.0|ICD10|Lymphocytic predominance|9651/3
C1266194|T191|ET|C81.4|ICD10CM|Lymphocyte-rich classical Hodgkin lymphoma|9651/3
C1266194|T191|AB|C81.4|ICD10CM|Lymphocyte-rich Hodgkin lymphoma|9651/3
C1266194|T191|HT|C81.4|ICD10CM|Lymphocyte-rich Hodgkin lymphoma|9651/3
C1266194|T191|HT|201.4|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance|9651/3
C1266194|T191|PT|MTHU083128|ICPC2ICD10ENG|disease; Hodgkin's, lymphocytic predominance|9651/3
C1266194|T191|PT|MTHU083124|ICPC2ICD10ENG|disease; Hodgkin's, lymphocytic-histiocytic predominance|9651/3
C1266194|T191|PT|MTHU035340|ICPC2ICD10ENG|Hodgkin; lymphocytic predominance|9651/3
C1266194|T191|PT|MTHU035335|ICPC2ICD10ENG|Hodgkin; lymphocytic-histiocytic predominance|9651/3
C1266194|T191|LLT|10020231|MDR|Hodgkin's disease lymphocyte predominance type stage unspecified|9651/3
C1266194|T191|PT|10020231|MDR|Hodgkin's disease lymphocyte predominance type stage unspecified|9651/3
C1266194|T191|LLT|10020281|MDR|Hodgkin's disease, lymphocytic-histiocytic predominance|9651/3
C1266194|T191|SY|31693|MEDCIN|Hodgkin's disease lymphocyte predominant|9651/3
C1266194|T191|SY|273312|MEDCIN|Hodgkin's disease with lymphocytic-histiocytic predominance|9651/3
C1266194|T191|PT|273312|MEDCIN|Hodgkin's disease, lymphocytic-histiocytic predominance|9651/3
C1266194|T191|PT|31693|MEDCIN|lymphocyte-rich Hodgkin lymphoma|9651/3
C1266194|T191|PM|D006689|MSH|Lymphocyte Rich Classical Hodgkin's Lymphoma|9651/3
C1266194|T191|PEP|D006689|MSH|Lymphocyte-Rich Classical Hodgkin's Lymphoma|9651/3
C1266194|T191|PN|NOCODE|MTH|Lymphocyte Rich Classical Hodgkin Lymphoma|9651/3
C1266194|T191|AB|C6913|NCI|LRCHL|9651/3
C1266194|T191|SY|C6913|NCI|Lymphocyte Rich Classical Hodgkin Lymphoma|9651/3
C1266194|T191|SY|C6913|NCI|Lymphocyte Rich Classical Hodgkin's Disease|9651/3
C1266194|T191|SY|C6913|NCI|Lymphocyte Rich Classical Hodgkin's Lymphoma|9651/3
C1266194|T191|SY|C6913|NCI|Lymphocyte Rich Hodgkin Lymphoma|9651/3
C1266194|T191|SY|C6913|NCI|Lymphocyte Rich Hodgkin's Disease|9651/3
C1266194|T191|SY|C6913|NCI|Lymphocyte Rich Hodgkin's Lymphoma|9651/3
C1266194|T191|PT|C6913|NCI|Lymphocyte-Rich Classic Hodgkin Lymphoma|9651/3
C1266194|T191|SY|C6913|NCI|Lymphocyte-Rich Classical Hodgkin Lymphoma|9651/3
C1266194|T191|SY|C6913|NCI|Lymphocyte-Rich Classical Hodgkin's Lymphoma|9651/3
C1266194|T191|PT|C6913|NCI_CPTAC|Lymphocyte-Rich Classic Hodgkin Lymphoma|9651/3
C1266194|T191|DN|C6913|NCI_CTRP|Lymphocyte-Rich Classical Hodgkin Lymphoma|9651/3
C1266194|T191|AB|B613.|RCD|Hodgkin dis, lymphocyt predom|9651/3
C1266194|T191|PT|B613.|RCD|Hodgkin's disease, lymphocytic predominance|9651/3
C1266194|T191|SY|B613.|RCD|Hodgkin's disease, lymphocytic-histiocytic predominance|9651/3
C1266194|T191|OP|B6130|RCD|Hodgkin's disease, lymphocytic-histiocytic predominance of unspecified site|9651/3
C1266194|T191|AB|B613.|RCD|Hodgkin's lympho-histio predom|9651/3
C1266194|T191|OP|B613z|RCD|Hodgkin's, lymphocytic-histiocytic predominance NOS|9651/3
C1266194|T191|OA|B6130|RCD|Hodgkin's, lymphocytic-histiocytic predominance unspec site|9651/3
C1266194|T191|OA|B6130|RCD|Lymph-histio-Hodgkin,unsp.site|9651/3
C1266194|T191|OA|B613z|RCD|Lympho-histiocytic Hodgkin NOS|9651/3
C1266194|T191|OP|BBj1.|RCDSY|Hodgkin's disease, lymphocytic predominance|9651/3
C1266194|T191|OA|BBj1.|RCDSY|Hodgkin's,lymphocytic pred.|9651/3
C1266194|T191|SY|128799007|SNOMEDCT_US|Classical Hodgkin lymphoma, lymphocyte-rich|9651/3
C1266194|T191|PT|128799007|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte-rich|9651/3
C1266194|T191|SY|118607005|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte-rich|9651/3
C1266194|T191|IS|118607005|SNOMEDCT_US|Hodgkin's disease, lymphocytic predominance|9651/3
C1266194|T191|OAP|59668005|SNOMEDCT_US|Hodgkin's disease, lymphocytic predominance|9651/3
C1266194|T191|IS|59668005|SNOMEDCT_US|Hodgkin's disease, lymphocytic predominance -RETIRED-|9651/3
C1266194|T191|OF|59668005|SNOMEDCT_US|Hodgkin's disease, lymphocytic predominance -RETIRED-|9651/3
C1266194|T191|IS|59668005|SNOMEDCT_US|Hodgkin's disease, lymphocytic predominance, NOS|9651/3
C1266194|T191|IS|59668005|SNOMEDCT_US|Hodgkin's disease, lymphocytic-histiocytic predominance|9651/3
C1266194|T191|OAP|188553001|SNOMEDCT_US|Hodgkin's disease, lymphocytic-histiocytic predominance of unspecified site|9651/3
C1266194|T191|OAP|188563009|SNOMEDCT_US|Hodgkin's, lymphocytic-histiocytic predominance NOS|9651/3
C1266194|T191|PT|118607005|SNOMEDCT_US|Lymphocyte-rich classical Hodgkin lymphoma|9651/3
C0152266|T191|PX|C81.2|ICD10|Hodgkin's disease with mixed cellularity|9652/3
C0152266|T191|PS|C81.2|ICD10|Mixed cellularity|9652/3
C0152266|T191|ET|C81.2|ICD10CM|Mixed cellularity classical Hodgkin lymphoma|9652/3
C0152266|T191|AB|C81.2|ICD10CM|Mixed cellularity Hodgkin lymphoma|9652/3
C0152266|T191|HT|C81.2|ICD10CM|Mixed cellularity Hodgkin lymphoma|9652/3
C0152266|T191|HT|201.6|ICD9CM|Hodgkin's disease, mixed cellularity|9652/3
C0152266|T191|PT|MTHU083122|ICPC2ICD10ENG|disease; Hodgkin's, mixed cellularity|9652/3
C0152266|T191|PT|MTHU035332|ICPC2ICD10ENG|Hodgkin; mixed cellularity|9652/3
C0152266|T191|LLT|10020232|MDR|Hodgkin's disease mixed cellularity|9652/3
C0152266|T191|PT|10020242|MDR|Hodgkin's disease mixed cellularity stage unspecified|9652/3
C0152266|T191|LLT|10020242|MDR|Hodgkin's disease mixed cellularity stage unspecified|9652/3
C0152266|T191|LLT|10020290|MDR|Hodgkin's disease, mixed cellularity|9652/3
C0152266|T191|PT|31694|MEDCIN|mixed cellularity Hodgkin's disease|9652/3
C0152266|T191|PEP|D006689|MSH|Mixed Cellularity Hodgkin's Lymphoma|9652/3
C0152266|T191|PN|NOCODE|MTH|Mixed Cellularity Hodgkin Lymphoma|9652/3
C0152266|T191|SY|C3517|NCI|Hodgkin's Disease Mixed Cellularity|9652/3
C0152266|T191|SY|C3517|NCI|Hodgkin's Lymphoma Mixed Cellularity|9652/3
C0152266|T191|AB|C3517|NCI|MCCHL|9652/3
C0152266|T191|AB|C3517|NCI|MCHL|9652/3
C0152266|T191|PT|C3517|NCI|Mixed Cellularity Classic Hodgkin Lymphoma|9652/3
C0152266|T191|SY|C3517|NCI|Mixed Cellularity Classical Hodgkin Lymphoma|9652/3
C0152266|T191|SY|CIBMTR|NCI|Mixed Cellularity Classical Hodgkin Lymphoma|9652/3
C0152266|T191|SY|C3517|NCI|Mixed Cellularity Hodgkin Lymphoma|9652/3
C0152266|T191|SY|C3517|NCI|Mixed Cellularity Hodgkin's Disease|9652/3
C0152266|T191|SY|C3517|NCI|Mixed Cellularity Hodgkin's Lymphoma|9652/3
C0152266|T191|PT|C3517|NCI_CPTAC|Mixed Cellularity Classic Hodgkin Lymphoma|9652/3
C0152266|T191|DN|C3517|NCI_CTRP|Mixed Cellularity Classical Hodgkin Lymphoma|9652/3
C0152266|T191|AB|B615.|RCD|Hodgkin's - mixed cellularity|9652/3
C0152266|T191|PT|B615.|RCD|Hodgkin's disease, mixed cellularity|9652/3
C0152266|T191|OP|B615z|RCD|Hodgkin's disease, mixed cellularity NOS|9652/3
C0152266|T191|OP|B6150|RCD|Hodgkin's disease, mixed cellularity of unspecified site|9652/3
C0152266|T191|OA|B6150|RCD|Hodgkin's mix cell-unspec site|9652/3
C0152266|T191|OA|B615z|RCD|Hodgkin's mixed cellular. NOS|9652/3
C0152266|T191|PT|BBj2.|RCDSY|Hodgkin's disease, mixed cellularity|9652/3
C0152266|T191|AB|BBj2.|RCDSY|Hodgkin's,mixed cellularity|9652/3
C0152266|T191|SY|41529000|SNOMEDCT_US|Classical Hodgkin lymphoma, mixed cellularity|9652/3
C0152266|T191|SY|118609008|SNOMEDCT_US|Hodgkin disease, mixed cellularity|9652/3
C0152266|T191|PT|41529000|SNOMEDCT_US|Hodgkin lymphoma, mixed cellularity|9652/3
C0152266|T191|SY|118609008|SNOMEDCT_US|Hodgkin mixed cellularity lymphoma|9652/3
C0152266|T191|SY|118609008|SNOMEDCT_US|Hodgkin's disease, mixed cellularity|9652/3
C0152266|T191|SY|41529000|SNOMEDCT_US|Hodgkin's disease, mixed cellularity|9652/3
C0152266|T191|OAP|188583005|SNOMEDCT_US|Hodgkin's disease, mixed cellularity NOS|9652/3
C0152266|T191|OAP|188574000|SNOMEDCT_US|Hodgkin's disease, mixed cellularity of unspecified site|9652/3
C0152266|T191|IS|41529000|SNOMEDCT_US|Hodgkin's disease, mixed cellularity, NOS|9652/3
C0152267|T191|PX|C81.3|ICD10|Hodgkin's disease with lymphocytic depletion|9653/3
C0152267|T191|PS|C81.3|ICD10|Lymphocytic depletion|9653/3
C0152267|T191|ET|C81.3|ICD10CM|Lymphocyte depleted classical Hodgkin lymphoma|9653/3
C0152267|T191|AB|C81.3|ICD10CM|Lymphocyte depleted Hodgkin lymphoma|9653/3
C0152267|T191|HT|C81.3|ICD10CM|Lymphocyte depleted Hodgkin lymphoma|9653/3
C0152267|T191|HT|201.7|ICD9CM|Hodgkin's disease, lymphocytic depletion|9653/3
C0152267|T191|PT|MTHU083125|ICPC2ICD10ENG|disease; Hodgkin's, lymphocytic depletion|9653/3
C0152267|T191|PT|MTHU035336|ICPC2ICD10ENG|Hodgkin; lymphocytic depletion|9653/3
C0152267|T191|LLT|10020219|MDR|Hodgkin's disease lymphocyte depletion type stage unspecified|9653/3
C0152267|T191|PT|10020219|MDR|Hodgkin's disease lymphocyte depletion type stage unspecified|9653/3
C0152267|T191|LLT|10020272|MDR|Hodgkin's disease, lymphocytic depletion|9653/3
C0152267|T191|PT|31692|MEDCIN|Hodgkin's disease lymphocytic depletion|9653/3
C0152267|T191|PEP|D006689|MSH|Lymphocyte Depletion Hodgkin's Lymphoma|9653/3
C0152267|T191|PN|NOCODE|MTH|Hodgkin lymphoma, lymphocyte depletion|9653/3
C0152267|T191|ET|201.7|MTHICD9|Hodgkin's disease, lymphocytic depletion NOS|9653/3
C0152267|T191|SY|C9283|NCI|Hodgkin Lymphoma Lymphocyte Depleted|9653/3
C0152267|T191|SY|C9283|NCI|Hodgkin's Disease Lymphocyte Depletion|9653/3
C0152267|T191|SY|C9283|NCI|Hodgkin's Lymphoma Lymphocyte Depleted|9653/3
C0152267|T191|AB|C9283|NCI|LDCHL|9653/3
C0152267|T191|AB|C9283|NCI|LDHL|9653/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Classical Hodgkin Lymphoma|9653/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Classical Hodgkin's Lymphoma|9653/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Hodgkin Lymphoma|9653/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Hodgkin's Disease|9653/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Hodgkin's Lymphoma|9653/3
C0152267|T191|PT|C9283|NCI|Lymphocyte-Depleted Classic Hodgkin Lymphoma|9653/3
C0152267|T191|SY|C9283|NCI|Lymphocyte-Depleted Classical Hodgkin Lymphoma|9653/3
C0152267|T191|SY|C9283|NCI|Lymphocyte-Depleted Hodgkin's Disease|9653/3
C0152267|T191|SY|C9283|NCI|Lymphocyte-Depleted Hodgkin's Lymphoma|9653/3
C0152267|T191|PT|C9283|NCI_CPTAC|Lymphocyte-Depleted Classic Hodgkin Lymphoma|9653/3
C0152267|T191|DN|C9283|NCI_CTRP|Lymphocyte-Depleted Classical Hodgkin Lymphoma|9653/3
C0152267|T191|PT|B616.|RCD|Hodgkin's disease, lymphocytic depletion|9653/3
C0152267|T191|OP|B616z|RCD|Hodgkin's disease, lymphocytic depletion NOS|9653/3
C0152267|T191|OA|B6160|RCD|Hodgkin's lymp.dep.-unsp. site|9653/3
C0152267|T191|OA|B616z|RCD|Hodgkin's lymphocyt. depl. NOS|9653/3
C0152267|T191|AB|B616.|RCD|Hodgkin's lymphocyt. depletion|9653/3
C0152267|T191|OP|B6160|RCD|Hodgkin's lymphocytic depletion of unspecified site|9653/3
C0152267|T191|OP|BBj3.|RCDSY|Hodgkin's disease, lymphocytic depletion NOS|9653/3
C0152267|T191|OA|BBj3.|RCDSY|Hodgkin's,lymphocyt.dep.NOS|9653/3
C0152267|T191|SY|112687003|SNOMEDCT_US|Classical Hodgkin lymphoma, lymphocyte depletion|9653/3
C0152267|T191|SY|118610003|SNOMEDCT_US|Hodgkin disease, lymphocytic depletion|9653/3
C0152267|T191|PT|112687003|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte depletion|9653/3
C0152267|T191|SY|118610003|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion|9653/3
C0152267|T191|SY|112687003|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion|9653/3
C0152267|T191|OAP|188594009|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion NOS|9653/3
C0152267|T191|IS|112687003|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion, NOS|9653/3
C0152267|T191|OAP|188584004|SNOMEDCT_US|Hodgkin's lymphocytic depletion of unspecified site|9653/3
C0334622|T191|PT|MTHU083126|ICPC2ICD10ENG|disease; Hodgkin's, lymphocytic depletion, diffuse fibrosis|9654/3
C0334622|T191|PT|MTHU035337|ICPC2ICD10ENG|Hodgkin; lymphocytic depletion, diffuse fibrosis|9654/3
C0334622|T191|PT|92516|MEDCIN|Hodgkin's disease lymphocyte depleted diffuse fibrosis|9654/3
C0334622|T191|ET|201.7|MTHICD9|Hodgkin's disease, lymphocytic depletion diffuse fibrosis|9654/3
C1881058|T191|OP|C66846|NCI|Hodgkin's Disease, Lymphocyte Depletion, Diffuse Fibrosis|9654/3
C1881058|T191|PT|C66846|NCI|Hodgkin's Disease, Lymphocyte Depletion, Diffuse Fibrosis|9654/3
C0334622|T191|AB|XaBBZ|RCD|Hodg,lymphocyt depl,dif fib|9654/3
C0334622|T191|PT|XaBBZ|RCD|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis|9654/3
C0334622|T191|PT|BBj4.|RCDSY|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis|9654/3
C0334622|T191|AB|BBj4.|RCDSY|Hodgkin's disease,lymphocytic depletion,diffuse fibrosis|9654/3
C0334622|T191|AB|BBj4.|RCDSY|Hodgkin's,lymp.dep.,dif.fib|9654/3
C0334622|T191|IS|16893006|SNOMEDCT_US|Classical Hodgkin lymphoma, lymphocyte depletion, diffuse fibrosis|9654/3
C0334622|T191|SY|16893006|SNOMEDCT_US|Classical Hodgkin lymphoma, lymphocyte depletion, diffuse fibrosis|9654/3
C0334622|T191|SY|307633009|SNOMEDCT_US|Hodgkin disease, lymphocytic depletion, diffuse fibrosis|9654/3
C0334622|T191|IS|16893006|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte depletion, diffuse fibrosis|9654/3
C0334622|T191|PT|16893006|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte depletion, diffuse fibrosis|9654/3
C0334622|T191|SY|16893006|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis|9654/3
C0334622|T191|PT|307633009|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis|9654/3
C0431137|T191|PT|MTHU083127|ICPC2ICD10ENG|disease; Hodgkin's, lymphocytic depletion, reticular|9655/3
C0431137|T191|PT|MTHU035339|ICPC2ICD10ENG|Hodgkin; lymphocytic depletion, reticular|9655/3
C0431137|T191|PT|92517|MEDCIN|Hodgkin's disease lymphocyte depleted reticular type|9655/3
C0431137|T191|PT|236529|MEDCIN|Hodgkin's lymphoma of lymph node with reticular lymphocytic depletion|9655/3
C0431137|T191|ET|201.7|MTHICD9|Hodgkin's disease, lymphocytic depletion reticular type|9655/3
C1881059|T191|OP|C66847|NCI|Hodgkin's Disease, Lymphocyte Depletion, Reticular|9655/3
C1881059|T191|PT|C66847|NCI|Hodgkin's Disease, Lymphocyte Depletion, Reticular|9655/3
C0431137|T191|AB|XaBBb|RCD|Hodg dis,lymphocyt depl,retic|9655/3
C0431137|T191|PT|XaBBb|RCD|Hodgkin's disease, lymphocytic depletion, reticular type|9655/3
C0431137|T191|PT|BBj5.|RCDSY|Hodgkin's disease, lymphocytic depletion, reticular type|9655/3
C0431137|T191|AB|BBj5.|RCDSY|Hodgkin's,lymp.dep.ret.type|9655/3
C0431137|T191|IS|71109004|SNOMEDCT_US|Classical Hodgkin lymphoma, lymphocyte depletion, reticular|9655/3
C0431137|T191|SY|71109004|SNOMEDCT_US|Classical Hodgkin lymphoma, lymphocyte depletion, reticular|9655/3
C0431137|T191|SY|307634003|SNOMEDCT_US|Hodgkin disease, lymphocytic depletion, reticular type|9655/3
C0431137|T191|IS|71109004|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte depletion, reticular|9655/3
C0431137|T191|PT|71109004|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte depletion, reticular|9655/3
C0431137|T191|SY|71109004|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion, reticular|9655/3
C0431137|T191|PT|307634003|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion, reticular type|9655/3
C1334968|T191|HT|C81.0|ICD10CM|Nodular lymphocyte predominant Hodgkin lymphoma|9659/3
C1334968|T191|AB|C81.0|ICD10CM|Nodular lymphocyte predominant Hodgkin lymphoma|9659/3
C2239290|T191|PT|MTHU083130|ICPC2ICD10ENG|disease; Hodgkin's, lymphocytic predominance, nodular|9659/3
C2239290|T191|PT|MTHU035342|ICPC2ICD10ENG|Hodgkin; lymphocytic predominance, nodular|9659/3
C1334968|T191|LLT|10080201|MDR|Nodular lymphocyte predominant Hodgkin lymphoma|9659/3
C1334968|T191|PT|10080201|MDR|Nodular lymphocyte predominant Hodgkin lymphoma|9659/3
C2239290|T191|SY|91367|MEDCIN|Hodgkin's disease lymphocyte predominant nodular|9659/3
C2239290|T191|PT|91367|MEDCIN|Hodgkin's disease lymphocyte predominant, nodular|9659/3
C2239290|T191|PT|273314|MEDCIN|nodular Hodgkin's disease with lymphocytic-histiocytic predominance|9659/3
C1334968|T191|PM|D006689|MSH|Nodular Lymphocyte Predominant Hodgkin's Lymphoma|9659/3
C1334968|T191|PEP|D006689|MSH|Nodular Lymphocyte-Predominant Hodgkin's Lymphoma|9659/3
C1334968|T191|ET|D006689|MSH|Nodular Sclerosing Hodgkin's Lymphoma|9659/3
C2239290|T191|PN|NOCODE|MTH|Hodgkin lymphoma, nodular lymphocyte predominance|9659/3
C1334968|T191|PN|NOCODE|MTH|Nodular Lymphocyte Predominant Hodgkin Lymphoma|9659/3
C1334968|T191|AB|C7258|NCI|NLPHL|9659/3
C1334968|T191|PT|C7258|NCI|Nodular Lymphocyte Predominant Hodgkin Lymphoma|9659/3
C1334968|T191|SY|TCGA|NCI|Nodular Lymphocyte Predominant Hodgkin Lymphoma|9659/3
C1334968|T191|SY|C7258|NCI|Nodular Lymphocyte Predominant Hodgkin's Lymphoma|9659/3
C1334968|T191|PT|C7258|NCI_CPTAC|Nodular Lymphocyte Predominant Hodgkin Lymphoma|9659/3
C1334968|T191|SY|10020231|NCI_CTEP-SDC|Hodgkin lymphoma nodular LP, NOS|9659/3
C1334968|T191|PT|10020231|NCI_CTEP-SDC|Hodgkin lymphoma nodular lymphocyte predominant type, NOS|9659/3
C1334968|T191|DN|C7258|NCI_CTRP|Nodular Lymphocyte Predominant Hodgkin Lymphoma|9659/3
C1334968|T191|PT|CDR0000574285|NCI_NCI-GLOSS|NLPHL|9659/3
C1334968|T191|PT|CDR0000574286|NCI_NCI-GLOSS|nodular lymphocyte-predominant Hodgkin lymphoma|9659/3
C2239290|T191|AB|Xa0St|RCD|Hodgk dis, lymph predomin-nod|9659/3
C2239290|T191|PT|Xa0St|RCD|Hodgkin's disease, lymphocytic predominance - nodular|9659/3
C2239290|T191|OA|BBj11|RCDSY|Hodgk,lymphocy predom,nodul|9659/3
C2239290|T191|OP|BBj11|RCDSY|Hodgkin,s disease, lymphocytic predominance, nodular|9659/3
C2239290|T191|OAS|277608004|SNOMEDCT_US|Hodgkin disease, lymphocytic predominance - nodular|9659/3
C2239290|T191|SY|70600005|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte predominance, nodular|9659/3
C2239290|T191|SY|118605002|SNOMEDCT_US|Hodgkin lymphoma, nodular lymphocyte predominance|9659/3
C2239290|T191|PT|70600005|SNOMEDCT_US|Hodgkin lymphoma, nodular lymphocyte predominance|9659/3
C2239290|T191|OAP|277608004|SNOMEDCT_US|Hodgkin's disease, lymphocytic predominance - nodular|9659/3
C2239290|T191|SY|70600005|SNOMEDCT_US|Hodgkin's disease, lymphocytic predominance, nodular|9659/3
C0019829|T191|ET|0000004628|AOD|Hodgkin's disease|9661/3
C0019829|T191|AB|BI00314|BI|hd|9661/3
C0019829|T191|PT|BI00314|BI|hodgkin's disease|9661/3
C0019829|T191|RT|BI00314|BI|hodgkin's lymphoma|9661/3
C0019829|T191|PT|1006070|CCPSS|LYMPHOMA HODGKIN|9661/3
C0019829|T191|SD|37|CCS|Hodgkin`s disease|9661/3
C0019829|T191|MD|2.10.1|CCS|Hodgkins disease|9661/3
C0019829|T191|SD|NEO057|CCSR_10|Hodgkin lymphoma|9661/3
C0019829|T191|SY|0000006210|CHV|HD|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkin disease|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkin lymphoma|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkin lymphomas|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkin's disease|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphoma|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphoma disease|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphomas|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkins disease|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkins diseases|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkins lymphoma|9661/3
C0019829|T191|SY|0000006210|CHV|hodgkins lymphomas|9661/3
C0019829|T191|SY|0000006210|CHV|lymphogranulomatosis|9661/3
C0019829|T191|PT|U000356|COSTAR|HODGKIN'S DISEASE|9661/3
C0019829|T191|PT|376|COSTAR|HODGKINS DISEASE|9661/3
C0019829|T191|PT|2004-1208|CSP|Hodgkin's disease|9661/3
C0019829|T191|ET|2004-1208|CSP|lymphogranulomatosis|9661/3
C0019829|T191|GT|LYMPHOMA LIKE REACT|CST|HODGINS|9661/3
C0019829|T191|DI|U000853|DXP|HODGKINS DISEASE|9661/3
C0019829|T191|SY|HP:0012189|HPO|Hodgkin disease|9661/3
C0019829|T191|PT|HP:0012189|HPO|Hodgkin lymphoma|9661/3
C0019829|T191|SY|HP:0012189|HPO|Hodgkin's lymphoma|9661/3
C0019829|T191|HT|C81|ICD10|Hodgkin's disease|9661/3
C0019829|T191|PT|C81.9|ICD10|Hodgkin's disease, unspecified|9661/3
C0019829|T191|AB|C81|ICD10CM|Hodgkin lymphoma|9661/3
C0019829|T191|HT|C81|ICD10CM|Hodgkin lymphoma|9661/3
C0019829|T191|AB|C81.9|ICD10CM|Hodgkin lymphoma, unspecified|9661/3
C0019829|T191|HT|C81.9|ICD10CM|Hodgkin lymphoma, unspecified|9661/3
C0019829|T191|HT|201|ICD9CM|Hodgkin's disease|9661/3
C0019829|T191|HT|201.9|ICD9CM|Hodgkin's disease, unspecified type|9661/3
C0019829|T191|HT|201.1|ICD9CM|Hodgkin's granuloma|9661/3
C0019829|T191|HT|201.0|ICD9CM|Hodgkin's paragranuloma|9661/3
C0019829|T191|HT|201.2|ICD9CM|Hodgkin's sarcoma|9661/3
C0019829|T191|PT|B72|ICPC|Hodgkins disease|9661/3
C0019829|T191|AB|B72|ICPC2EENG|Hodgkin's disease/lymphoma|9661/3
C0019829|T191|PT|B72|ICPC2EENG|Hodgkin's disease/lymphoma|9661/3
C0019829|T191|PT|MTHU083121|ICPC2ICD10ENG|disease; Hodgkin|9661/3
C0019829|T191|PT|MTHU032756|ICPC2ICD10ENG|granuloma; Hodgkin|9661/3
C0019829|T191|PT|MTHU032780|ICPC2ICD10ENG|granuloma; malignant|9661/3
C0019829|T191|PT|MTHU035331|ICPC2ICD10ENG|Hodgkin|9661/3
C0019829|T191|PT|MTHU035334|ICPC2ICD10ENG|Hodgkin; granuloma|9661/3
C0019829|T191|PT|MTHU035344|ICPC2ICD10ENG|Hodgkin; lymphoma|9661/3
C0019829|T191|PT|MTHU035351|ICPC2ICD10ENG|Hodgkin; paragranuloma|9661/3
C0019829|T191|PT|MTHU035352|ICPC2ICD10ENG|Hodgkin; sarcoma|9661/3
C0019829|T191|PT|MTHU046802|ICPC2ICD10ENG|lymphoma; Hodgkin|9661/3
C0019829|T191|PT|MTHU047288|ICPC2ICD10ENG|malignant; granuloma|9661/3
C0019829|T191|PT|MTHU057409|ICPC2ICD10ENG|paragranuloma; Hodgkin|9661/3
C0019829|T191|PT|MTHU065903|ICPC2ICD10ENG|sarcoma; Hodgkin|9661/3
C0019829|T191|PT|B72001|ICPC2P|Disease;Hodgkins|9661/3
C0019829|T191|PTN|B72001|ICPC2P|Hodgkins disease|9661/3
C0019829|T191|PTN|B72003|ICPC2P|hodgkins lymphoma|9661/3
C0019829|T191|PTN|B72004|ICPC2P|Hodgkins sarcoma|9661/3
C0019829|T191|PT|B72003|ICPC2P|Lymphoma;Hodgkins|9661/3
C0019829|T191|PT|B72004|ICPC2P|Sarcoma;Hodgkins|9661/3
C0019829|T191|PT|U002210|LCH|Hodgkin's disease|9661/3
C0019829|T191|PT|sh85061347|LCH_NW|Hodgkin's disease|9661/3
C0019829|T191|LA|LA26792-4|LNC|Hodgkin lymphoma|9661/3
C0019829|T191|OL|10020205|MDR|Hodgins|9661/3
C0019829|T191|LLT|10020206|MDR|Hodgkin's disease|9661/3
C0019829|T191|PT|10020206|MDR|Hodgkin's disease|9661/3
C0019829|T191|LLT|10020255|MDR|Hodgkin's disease NOS|9661/3
C0019829|T191|LLT|10020309|MDR|Hodgkin's disease, unspecified type|9661/3
C0019829|T191|LLT|10020318|MDR|Hodgkin's granuloma|9661/3
C0019829|T191|LLT|10020328|MDR|Hodgkin's lymphoma|9661/3
C0019829|T191|LLT|10020329|MDR|Hodgkin's paragranuloma|9661/3
C0019829|T191|LLT|10020339|MDR|Hodgkin's sarcoma|9661/3
C0019829|T191|LLT|10063666|MDR|Lymphogranulomatosis|9661/3
C0019829|T191|HG|10025319|MDR|Lymphomas Hodgkin's disease|9661/3
C0019829|T191|PT|31691|MEDCIN|Hodgkin disease|9661/3
C0019829|T191|PT|92514|MEDCIN|Hodgkin disease granuloma|9661/3
C0019829|T191|PT|92513|MEDCIN|Hodgkin disease paragranuloma|9661/3
C0019829|T191|PT|92515|MEDCIN|Hodgkin disease sarcoma|9661/3
C0019829|T191|PT|1262|MEDLINEPLUS|Hodgkin Disease|9661/3
C0019829|T191|SY|1262|MEDLINEPLUS|Hodgkin lymphoma|9661/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkin|9661/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkin's|9661/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkins|9661/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkin|9661/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkin's|9661/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkins|9661/3
C0019829|T191|ET|D006689|MSH|Granuloma, Malignant|9661/3
C0019829|T191|DEV|D006689|MSH|HODGKIN DIS|9661/3
C0019829|T191|MH|D006689|MSH|Hodgkin Disease|9661/3
C0019829|T191|PM|D006689|MSH|Hodgkin Granuloma|9661/3
C0019829|T191|ET|D006689|MSH|Hodgkin Lymphoma|9661/3
C0019829|T191|ET|D006689|MSH|Hodgkin's Disease|9661/3
C0019829|T191|PM|D006689|MSH|Hodgkin's Granuloma|9661/3
C0019829|T191|ET|D006689|MSH|Hodgkin's Lymphoma|9661/3
C0019829|T191|DEV|D006689|MSH|HODGKINS DIS|9661/3
C0019829|T191|ET|D006689|MSH|Hodgkins Disease|9661/3
C0019829|T191|PM|D006689|MSH|Hodgkins Granuloma|9661/3
C0019829|T191|PM|D006689|MSH|Hodgkins Lymphoma|9661/3
C0019829|T191|ET|D006689|MSH|Lymphogranuloma, Malignant|9661/3
C0019829|T191|PM|D006689|MSH|Lymphogranulomas, Malignant|9661/3
C0019829|T191|PM|D006689|MSH|Lymphoma, Hodgkin|9661/3
C0019829|T191|PM|D006689|MSH|Lymphoma, Hodgkin's|9661/3
C0019829|T191|PM|D006689|MSH|Malignant Granuloma|9661/3
C0019829|T191|PM|D006689|MSH|Malignant Granulomas|9661/3
C0019829|T191|PM|D006689|MSH|Malignant Lymphogranuloma|9661/3
C0019829|T191|PM|D006689|MSH|Malignant Lymphogranulomas|9661/3
C0019829|T191|PN|NOCODE|MTH|Hodgkin Disease|9661/3
C0019829|T191|PT|376|MTH|Hodgkin's Disease|9661/3
C0019829|T191|ET|201.9|MTHICD9|Hodgkin's disease NOS|9661/3
C0019829|T191|ET|201.9|MTHICD9|Hodgkin's lymphoma NOS|9661/3
C0019829|T191|ET|201.9|MTHICD9|Malignant lymphogranuloma|9661/3
C0019829|T191|ET|201.9|MTHICD9|Malignant lymphogranulomatosis|9661/3
C0019829|T191|AB|C9357|NCI|HL|9661/3
C0019829|T191|PT|C9357|NCI|Hodgkin Lymphoma|9661/3
C0019829|T191|SY|C9357|NCI|Hodgkin's Disease|9661/3
C0019829|T191|OP|C6914|NCI|Hodgkin's Granuloma|9661/3
C0019829|T191|PT|C6914|NCI|Hodgkin's Granuloma|9661/3
C0019829|T191|SY|C9357|NCI|Hodgkin's Lymphoma|9661/3
C0019829|T191|OP|C26956|NCI|Hodgkin's Paragranuloma|9661/3
C0019829|T191|PT|C26956|NCI|Hodgkin's Paragranuloma|9661/3
C0019829|T191|PT|C9357|NCI_CPTAC|Hodgkin Lymphoma|9661/3
C0019829|T191|SY|C9357|NCI_CPTAC|Hodgkin's Disease|9661/3
C0019829|T191|PT|C26956|NCI_CPTAC|Hodgkins Paragranuloma|9661/3
C0019829|T191|PT|10020255|NCI_CTEP-SDC|Hodgkin lymphoma, NOS|9661/3
C0019829|T191|DN|C9357|NCI_CTRP|Hodgkin Lymphoma|9661/3
C0019829|T191|PT|C9357|NCI_CTRP|Hodgkin Lymphoma|9661/3
C0019829|T191|PT|CDR0000045012|NCI_NCI-GLOSS|Hodgkin disease|9661/3
C0019829|T191|PT|CDR0000270800|NCI_NCI-GLOSS|Hodgkin lymphoma|9661/3
C0019829|T191|PT|C9357|NCI_NICHD|Hodgkin Lymphoma|9661/3
C0019829|T191|SY|C9357|NCI_NICHD|Hodgkin's Disease|9661/3
C0019829|T191|SY|C9357|NCI_NICHD|Hodgkin's Lymphoma|9661/3
C0019829|T191|AB|CDR0000041646|PDQ|HL|9661/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkin disease|9661/3
C0019829|T191|PT|CDR0000041646|PDQ|Hodgkin lymphoma|9661/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkin's disease|9661/3
C0019829|T191|LV|CDR0000041646|PDQ|Hodgkin's lymphoma|9661/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkins disease|9661/3
C0019829|T191|LV|CDR0000041646|PDQ|Hodgkins lymphoma|9661/3
C0019829|T191|PT|R0121435|QMR|HODGKINS DISEASE SYSTEMIC|9661/3
C0019829|T191|SY|B61..|RCD|HD - Hodgkin's disease|9661/3
C0019829|T191|OA|B61z0|RCD|Hodgkin's dis.NOS-unspec. site|9661/3
C0019829|T191|PT|B61..|RCD|Hodgkin's disease|9661/3
C0019829|T191|OP|B61z.|RCD|Hodgkin's disease NOS|9661/3
C0019829|T191|OP|B61z0|RCD|Hodgkin's disease NOS, unspecified site|9661/3
C0019829|T191|PT|B611.|RCD|Hodgkin's granuloma|9661/3
C0019829|T191|OP|B611z|RCD|Hodgkin's granuloma NOS|9661/3
C0019829|T191|OP|B6110|RCD|Hodgkin's granuloma of unspecified site|9661/3
C0019829|T191|OA|B6110|RCD|Hodgkin's granuloma-unsp. site|9661/3
C0019829|T191|OA|B6100|RCD|Hodgkin's paragran-unspec site|9661/3
C0019829|T191|PT|B610.|RCD|Hodgkin's paragranuloma|9661/3
C0019829|T191|OP|B610z|RCD|Hodgkin's paragranuloma NOS|9661/3
C0019829|T191|OP|B6100|RCD|Hodgkin's paragranuloma of unspecified site|9661/3
C0019829|T191|PT|B612.|RCD|Hodgkin's sarcoma|9661/3
C0019829|T191|OP|B612z|RCD|Hodgkin's sarcoma NOS|9661/3
C0019829|T191|OP|B6120|RCD|Hodgkin's sarcoma of unspecified site|9661/3
C0019829|T191|OA|B6120|RCD|Hodgkin's sarcoma-unspec. site|9661/3
C0019829|T191|SY|B61..|RCD|Malignant Hodgkin's lymphoma|9661/3
C0019829|T191|PT|BBj..|RCDSY|Hodgkin's disease|9661/3
C0019829|T191|OP|XaC2n|RCDSY|Hodgkin's disease NOS|9661/3
C0019829|T191|OP|BBj9.|RCDSY|Hodgkin's granuloma|9661/3
C0019829|T191|OP|BBj8.|RCDSY|Hodgkin's paragranuloma|9661/3
C0019829|T191|OP|BBjA.|RCDSY|Hodgkin's sarcoma|9661/3
C0019829|T191|OP|XE1we|RCDSY|Lymphogranuloma, malignant|9661/3
C0019829|T191|SY|118599009|SNOMEDCT_US|HD - Hodgkin's disease|9661/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Hodgkin disease|9661/3
C0019829|T191|SY|118602004|SNOMEDCT_US|Hodgkin granuloma|9661/3
C0019829|T191|PT|14537002|SNOMEDCT_US|Hodgkin lymphoma|9661/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin lymphoma, no ICD-O subtype|9661/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype|9661/3
C0019829|T191|SY|118606001|SNOMEDCT_US|Hodgkin sarcoma|9661/3
C0019829|T191|OAP|154582001|SNOMEDCT_US|Hodgkin's disease|9661/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin's disease|9661/3
C0019829|T191|OF|154582001|SNOMEDCT_US|Hodgkin's disease|9661/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Hodgkin's disease|9661/3
C0019829|T191|OAP|188595005|SNOMEDCT_US|Hodgkin's disease NOS|9661/3
C0019829|T191|OAP|188605006|SNOMEDCT_US|Hodgkin's disease NOS|9661/3
C0019829|T191|OF|188605006|SNOMEDCT_US|Hodgkin's disease NOS|9661/3
C0019829|T191|OAP|188596006|SNOMEDCT_US|Hodgkin's disease NOS, unspecified site|9661/3
C0019829|T191|IS|14537002|SNOMEDCT_US|Hodgkin's disease, NOS|9661/3
C0019829|T191|SY|74189002|SNOMEDCT_US|Hodgkin's granuloma|9661/3
C0019829|T191|SY|118602004|SNOMEDCT_US|Hodgkin's granuloma|9661/3
C0019829|T191|OAP|188542007|SNOMEDCT_US|Hodgkin's granuloma NOS|9661/3
C0019829|T191|OAP|188533000|SNOMEDCT_US|Hodgkin's granuloma of unspecified site|9661/3
C0019829|T191|OAP|52337003|SNOMEDCT_US|Hodgkin's paragranuloma|9661/3
C0019829|T191|OAP|188521005|SNOMEDCT_US|Hodgkin's paragranuloma|9661/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma -RETIRED-|9661/3
C0019829|T191|OF|52337003|SNOMEDCT_US|Hodgkin's paragranuloma -RETIRED-|9661/3
C0019829|T191|OAP|188532005|SNOMEDCT_US|Hodgkin's paragranuloma NOS|9661/3
C0019829|T191|OAP|188522003|SNOMEDCT_US|Hodgkin's paragranuloma of unspecified site|9661/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma, nodular|9661/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma, NOS|9661/3
C0019829|T191|SY|46923007|SNOMEDCT_US|Hodgkin's sarcoma|9661/3
C0019829|T191|SY|118606001|SNOMEDCT_US|Hodgkin's sarcoma|9661/3
C0019829|T191|OAP|188552006|SNOMEDCT_US|Hodgkin's sarcoma NOS|9661/3
C0019829|T191|OAP|188543002|SNOMEDCT_US|Hodgkin's sarcoma of unspecified site|9661/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Lymphoma, Hodgkins|9661/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Malignant Hodgkin's lymphoma|9661/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Malignant lymphoma, Hodgkin's|9661/3
C0019829|T191|ET|0000004628|AOD|Hodgkin's disease|9662/3
C0019829|T191|AB|BI00314|BI|hd|9662/3
C0019829|T191|PT|BI00314|BI|hodgkin's disease|9662/3
C0019829|T191|RT|BI00314|BI|hodgkin's lymphoma|9662/3
C0019829|T191|PT|1006070|CCPSS|LYMPHOMA HODGKIN|9662/3
C0019829|T191|SD|37|CCS|Hodgkin`s disease|9662/3
C0019829|T191|MD|2.10.1|CCS|Hodgkins disease|9662/3
C0019829|T191|SD|NEO057|CCSR_10|Hodgkin lymphoma|9662/3
C0019829|T191|SY|0000006210|CHV|HD|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkin disease|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkin lymphoma|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkin lymphomas|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkin's disease|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphoma|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphoma disease|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkin's lymphomas|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkins disease|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkins diseases|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkins lymphoma|9662/3
C0019829|T191|SY|0000006210|CHV|hodgkins lymphomas|9662/3
C0019829|T191|SY|0000006210|CHV|lymphogranulomatosis|9662/3
C0019829|T191|PT|U000356|COSTAR|HODGKIN'S DISEASE|9662/3
C0019829|T191|PT|376|COSTAR|HODGKINS DISEASE|9662/3
C0019829|T191|PT|2004-1208|CSP|Hodgkin's disease|9662/3
C0019829|T191|ET|2004-1208|CSP|lymphogranulomatosis|9662/3
C0019829|T191|GT|LYMPHOMA LIKE REACT|CST|HODGINS|9662/3
C0019829|T191|DI|U000853|DXP|HODGKINS DISEASE|9662/3
C0019829|T191|SY|HP:0012189|HPO|Hodgkin disease|9662/3
C0019829|T191|PT|HP:0012189|HPO|Hodgkin lymphoma|9662/3
C0019829|T191|SY|HP:0012189|HPO|Hodgkin's lymphoma|9662/3
C0019829|T191|HT|C81|ICD10|Hodgkin's disease|9662/3
C0152267|T191|PX|C81.3|ICD10|Hodgkin's disease with lymphocytic depletion|9662/3
C0019829|T191|PT|C81.9|ICD10|Hodgkin's disease, unspecified|9662/3
C0152267|T191|PS|C81.3|ICD10|Lymphocytic depletion|9662/3
C0019829|T191|HT|C81|ICD10CM|Hodgkin lymphoma|9662/3
C0019829|T191|AB|C81|ICD10CM|Hodgkin lymphoma|9662/3
C0019829|T191|AB|C81.9|ICD10CM|Hodgkin lymphoma, unspecified|9662/3
C0019829|T191|HT|C81.9|ICD10CM|Hodgkin lymphoma, unspecified|9662/3
C0152267|T191|ET|C81.3|ICD10CM|Lymphocyte depleted classical Hodgkin lymphoma|9662/3
C0152267|T191|AB|C81.3|ICD10CM|Lymphocyte depleted Hodgkin lymphoma|9662/3
C0152267|T191|HT|C81.3|ICD10CM|Lymphocyte depleted Hodgkin lymphoma|9662/3
C0019829|T191|HT|201|ICD9CM|Hodgkin's disease|9662/3
C0152267|T191|HT|201.7|ICD9CM|Hodgkin's disease, lymphocytic depletion|9662/3
C0019829|T191|HT|201.9|ICD9CM|Hodgkin's disease, unspecified type|9662/3
C0019829|T191|HT|201.1|ICD9CM|Hodgkin's granuloma|9662/3
C0019829|T191|HT|201.0|ICD9CM|Hodgkin's paragranuloma|9662/3
C0019829|T191|HT|201.2|ICD9CM|Hodgkin's sarcoma|9662/3
C0019829|T191|PT|B72|ICPC|Hodgkins disease|9662/3
C0019829|T191|AB|B72|ICPC2EENG|Hodgkin's disease/lymphoma|9662/3
C0019829|T191|PT|B72|ICPC2EENG|Hodgkin's disease/lymphoma|9662/3
C0019829|T191|PT|MTHU083121|ICPC2ICD10ENG|disease; Hodgkin|9662/3
C0152267|T191|PT|MTHU083125|ICPC2ICD10ENG|disease; Hodgkin's, lymphocytic depletion|9662/3
C0019829|T191|PT|MTHU032756|ICPC2ICD10ENG|granuloma; Hodgkin|9662/3
C0019829|T191|PT|MTHU032780|ICPC2ICD10ENG|granuloma; malignant|9662/3
C0019829|T191|PT|MTHU035331|ICPC2ICD10ENG|Hodgkin|9662/3
C0019829|T191|PT|MTHU035334|ICPC2ICD10ENG|Hodgkin; granuloma|9662/3
C0152267|T191|PT|MTHU035336|ICPC2ICD10ENG|Hodgkin; lymphocytic depletion|9662/3
C0019829|T191|PT|MTHU035344|ICPC2ICD10ENG|Hodgkin; lymphoma|9662/3
C0019829|T191|PT|MTHU035351|ICPC2ICD10ENG|Hodgkin; paragranuloma|9662/3
C0019829|T191|PT|MTHU035352|ICPC2ICD10ENG|Hodgkin; sarcoma|9662/3
C0019829|T191|PT|MTHU046802|ICPC2ICD10ENG|lymphoma; Hodgkin|9662/3
C0019829|T191|PT|MTHU047288|ICPC2ICD10ENG|malignant; granuloma|9662/3
C0019829|T191|PT|MTHU057409|ICPC2ICD10ENG|paragranuloma; Hodgkin|9662/3
C0019829|T191|PT|MTHU065903|ICPC2ICD10ENG|sarcoma; Hodgkin|9662/3
C0019829|T191|PT|B72001|ICPC2P|Disease;Hodgkins|9662/3
C0019829|T191|PTN|B72001|ICPC2P|Hodgkins disease|9662/3
C0019829|T191|PTN|B72003|ICPC2P|hodgkins lymphoma|9662/3
C0019829|T191|PTN|B72004|ICPC2P|Hodgkins sarcoma|9662/3
C0019829|T191|PT|B72003|ICPC2P|Lymphoma;Hodgkins|9662/3
C0019829|T191|PT|B72004|ICPC2P|Sarcoma;Hodgkins|9662/3
C0019829|T191|PT|U002210|LCH|Hodgkin's disease|9662/3
C0019829|T191|PT|sh85061347|LCH_NW|Hodgkin's disease|9662/3
C0019829|T191|LA|LA26792-4|LNC|Hodgkin lymphoma|9662/3
C0019829|T191|OL|10020205|MDR|Hodgins|9662/3
C0019829|T191|PT|10020206|MDR|Hodgkin's disease|9662/3
C0019829|T191|LLT|10020206|MDR|Hodgkin's disease|9662/3
C0152267|T191|LLT|10020219|MDR|Hodgkin's disease lymphocyte depletion type stage unspecified|9662/3
C0152267|T191|PT|10020219|MDR|Hodgkin's disease lymphocyte depletion type stage unspecified|9662/3
C0019829|T191|LLT|10020255|MDR|Hodgkin's disease NOS|9662/3
C0152267|T191|LLT|10020272|MDR|Hodgkin's disease, lymphocytic depletion|9662/3
C0019829|T191|LLT|10020309|MDR|Hodgkin's disease, unspecified type|9662/3
C0019829|T191|LLT|10020318|MDR|Hodgkin's granuloma|9662/3
C0019829|T191|LLT|10020328|MDR|Hodgkin's lymphoma|9662/3
C0019829|T191|LLT|10020329|MDR|Hodgkin's paragranuloma|9662/3
C0019829|T191|LLT|10020339|MDR|Hodgkin's sarcoma|9662/3
C0019829|T191|LLT|10063666|MDR|Lymphogranulomatosis|9662/3
C0019829|T191|HG|10025319|MDR|Lymphomas Hodgkin's disease|9662/3
C0019829|T191|PT|31691|MEDCIN|Hodgkin disease|9662/3
C0019829|T191|PT|92514|MEDCIN|Hodgkin disease granuloma|9662/3
C0019829|T191|PT|92513|MEDCIN|Hodgkin disease paragranuloma|9662/3
C0019829|T191|PT|92515|MEDCIN|Hodgkin disease sarcoma|9662/3
C0152267|T191|PT|31692|MEDCIN|Hodgkin's disease lymphocytic depletion|9662/3
C0019829|T191|PT|1262|MEDLINEPLUS|Hodgkin Disease|9662/3
C0019829|T191|SY|1262|MEDLINEPLUS|Hodgkin lymphoma|9662/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkin|9662/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkin's|9662/3
C0019829|T191|PM|D006689|MSH|Disease, Hodgkins|9662/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkin|9662/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkin's|9662/3
C0019829|T191|ET|D006689|MSH|Granuloma, Hodgkins|9662/3
C0019829|T191|ET|D006689|MSH|Granuloma, Malignant|9662/3
C0019829|T191|DEV|D006689|MSH|HODGKIN DIS|9662/3
C0019829|T191|MH|D006689|MSH|Hodgkin Disease|9662/3
C0019829|T191|PM|D006689|MSH|Hodgkin Granuloma|9662/3
C0019829|T191|ET|D006689|MSH|Hodgkin Lymphoma|9662/3
C0019829|T191|ET|D006689|MSH|Hodgkin's Disease|9662/3
C0019829|T191|PM|D006689|MSH|Hodgkin's Granuloma|9662/3
C0019829|T191|ET|D006689|MSH|Hodgkin's Lymphoma|9662/3
C0019829|T191|DEV|D006689|MSH|HODGKINS DIS|9662/3
C0019829|T191|ET|D006689|MSH|Hodgkins Disease|9662/3
C0019829|T191|PM|D006689|MSH|Hodgkins Granuloma|9662/3
C0019829|T191|PM|D006689|MSH|Hodgkins Lymphoma|9662/3
C0152267|T191|PEP|D006689|MSH|Lymphocyte Depletion Hodgkin's Lymphoma|9662/3
C0019829|T191|ET|D006689|MSH|Lymphogranuloma, Malignant|9662/3
C0019829|T191|PM|D006689|MSH|Lymphogranulomas, Malignant|9662/3
C0019829|T191|PM|D006689|MSH|Lymphoma, Hodgkin|9662/3
C0019829|T191|PM|D006689|MSH|Lymphoma, Hodgkin's|9662/3
C0019829|T191|PM|D006689|MSH|Malignant Granuloma|9662/3
C0019829|T191|PM|D006689|MSH|Malignant Granulomas|9662/3
C0019829|T191|PM|D006689|MSH|Malignant Lymphogranuloma|9662/3
C0019829|T191|PM|D006689|MSH|Malignant Lymphogranulomas|9662/3
C0019829|T191|PN|NOCODE|MTH|Hodgkin Disease|9662/3
C0152267|T191|PN|NOCODE|MTH|Hodgkin lymphoma, lymphocyte depletion|9662/3
C0019829|T191|PT|376|MTH|Hodgkin's Disease|9662/3
C0019829|T191|ET|201.9|MTHICD9|Hodgkin's disease NOS|9662/3
C0152267|T191|ET|201.7|MTHICD9|Hodgkin's disease, lymphocytic depletion NOS|9662/3
C0019829|T191|ET|201.9|MTHICD9|Hodgkin's lymphoma NOS|9662/3
C0019829|T191|ET|201.9|MTHICD9|Malignant lymphogranuloma|9662/3
C0019829|T191|ET|201.9|MTHICD9|Malignant lymphogranulomatosis|9662/3
C0019829|T191|AB|C9357|NCI|HL|9662/3
C0019829|T191|PT|C9357|NCI|Hodgkin Lymphoma|9662/3
C0152267|T191|SY|C9283|NCI|Hodgkin Lymphoma Lymphocyte Depleted|9662/3
C0019829|T191|SY|C9357|NCI|Hodgkin's Disease|9662/3
C0152267|T191|SY|C9283|NCI|Hodgkin's Disease Lymphocyte Depletion|9662/3
C0019829|T191|PT|C6914|NCI|Hodgkin's Granuloma|9662/3
C0019829|T191|OP|C6914|NCI|Hodgkin's Granuloma|9662/3
C0019829|T191|SY|C9357|NCI|Hodgkin's Lymphoma|9662/3
C0152267|T191|SY|C9283|NCI|Hodgkin's Lymphoma Lymphocyte Depleted|9662/3
C0019829|T191|PT|C26956|NCI|Hodgkin's Paragranuloma|9662/3
C0019829|T191|OP|C26956|NCI|Hodgkin's Paragranuloma|9662/3
C0152267|T191|AB|C9283|NCI|LDCHL|9662/3
C0152267|T191|AB|C9283|NCI|LDHL|9662/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Classical Hodgkin Lymphoma|9662/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Classical Hodgkin's Lymphoma|9662/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Hodgkin Lymphoma|9662/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Hodgkin's Disease|9662/3
C0152267|T191|SY|C9283|NCI|Lymphocyte Depleted Hodgkin's Lymphoma|9662/3
C0152267|T191|PT|C9283|NCI|Lymphocyte-Depleted Classic Hodgkin Lymphoma|9662/3
C0152267|T191|SY|C9283|NCI|Lymphocyte-Depleted Classical Hodgkin Lymphoma|9662/3
C0152267|T191|SY|C9283|NCI|Lymphocyte-Depleted Hodgkin's Disease|9662/3
C0152267|T191|SY|C9283|NCI|Lymphocyte-Depleted Hodgkin's Lymphoma|9662/3
C0019829|T191|PT|C9357|NCI_CPTAC|Hodgkin Lymphoma|9662/3
C0019829|T191|SY|C9357|NCI_CPTAC|Hodgkin's Disease|9662/3
C0019829|T191|PT|C26956|NCI_CPTAC|Hodgkins Paragranuloma|9662/3
C0152267|T191|PT|C9283|NCI_CPTAC|Lymphocyte-Depleted Classic Hodgkin Lymphoma|9662/3
C0019829|T191|PT|10020255|NCI_CTEP-SDC|Hodgkin lymphoma, NOS|9662/3
C0019829|T191|PT|C9357|NCI_CTRP|Hodgkin Lymphoma|9662/3
C0019829|T191|DN|C9357|NCI_CTRP|Hodgkin Lymphoma|9662/3
C0152267|T191|DN|C9283|NCI_CTRP|Lymphocyte-Depleted Classical Hodgkin Lymphoma|9662/3
C0019829|T191|PT|CDR0000045012|NCI_NCI-GLOSS|Hodgkin disease|9662/3
C0019829|T191|PT|CDR0000270800|NCI_NCI-GLOSS|Hodgkin lymphoma|9662/3
C0019829|T191|PT|C9357|NCI_NICHD|Hodgkin Lymphoma|9662/3
C0019829|T191|SY|C9357|NCI_NICHD|Hodgkin's Disease|9662/3
C0019829|T191|SY|C9357|NCI_NICHD|Hodgkin's Lymphoma|9662/3
C0019829|T191|AB|CDR0000041646|PDQ|HL|9662/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkin disease|9662/3
C0019829|T191|PT|CDR0000041646|PDQ|Hodgkin lymphoma|9662/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkin's disease|9662/3
C0019829|T191|LV|CDR0000041646|PDQ|Hodgkin's lymphoma|9662/3
C0019829|T191|SY|CDR0000041646|PDQ|Hodgkins disease|9662/3
C0019829|T191|LV|CDR0000041646|PDQ|Hodgkins lymphoma|9662/3
C0019829|T191|PT|R0121435|QMR|HODGKINS DISEASE SYSTEMIC|9662/3
C0019829|T191|SY|B61..|RCD|HD - Hodgkin's disease|9662/3
C0019829|T191|OA|B61z0|RCD|Hodgkin's dis.NOS-unspec. site|9662/3
C0019829|T191|PT|B61..|RCD|Hodgkin's disease|9662/3
C0019829|T191|OP|B61z.|RCD|Hodgkin's disease NOS|9662/3
C0019829|T191|OP|B61z0|RCD|Hodgkin's disease NOS, unspecified site|9662/3
C0152267|T191|PT|B616.|RCD|Hodgkin's disease, lymphocytic depletion|9662/3
C0152267|T191|OP|B616z|RCD|Hodgkin's disease, lymphocytic depletion NOS|9662/3
C0019829|T191|PT|B611.|RCD|Hodgkin's granuloma|9662/3
C0019829|T191|OP|B611z|RCD|Hodgkin's granuloma NOS|9662/3
C0019829|T191|OP|B6110|RCD|Hodgkin's granuloma of unspecified site|9662/3
C0019829|T191|OA|B6110|RCD|Hodgkin's granuloma-unsp. site|9662/3
C0152267|T191|OA|B6160|RCD|Hodgkin's lymp.dep.-unsp. site|9662/3
C0152267|T191|OA|B616z|RCD|Hodgkin's lymphocyt. depl. NOS|9662/3
C0152267|T191|AB|B616.|RCD|Hodgkin's lymphocyt. depletion|9662/3
C0152267|T191|OP|B6160|RCD|Hodgkin's lymphocytic depletion of unspecified site|9662/3
C0019829|T191|OA|B6100|RCD|Hodgkin's paragran-unspec site|9662/3
C0019829|T191|PT|B610.|RCD|Hodgkin's paragranuloma|9662/3
C0019829|T191|OP|B610z|RCD|Hodgkin's paragranuloma NOS|9662/3
C0019829|T191|OP|B6100|RCD|Hodgkin's paragranuloma of unspecified site|9662/3
C0019829|T191|PT|B612.|RCD|Hodgkin's sarcoma|9662/3
C0019829|T191|OP|B612z|RCD|Hodgkin's sarcoma NOS|9662/3
C0019829|T191|OP|B6120|RCD|Hodgkin's sarcoma of unspecified site|9662/3
C0019829|T191|OA|B6120|RCD|Hodgkin's sarcoma-unspec. site|9662/3
C0019829|T191|SY|B61..|RCD|Malignant Hodgkin's lymphoma|9662/3
C0019829|T191|PT|BBj..|RCDSY|Hodgkin's disease|9662/3
C0019829|T191|OP|XaC2n|RCDSY|Hodgkin's disease NOS|9662/3
C0152267|T191|OP|BBj3.|RCDSY|Hodgkin's disease, lymphocytic depletion NOS|9662/3
C0019829|T191|OP|BBj9.|RCDSY|Hodgkin's granuloma|9662/3
C0019829|T191|OP|BBj8.|RCDSY|Hodgkin's paragranuloma|9662/3
C0019829|T191|OP|BBjA.|RCDSY|Hodgkin's sarcoma|9662/3
C0152267|T191|OA|BBj3.|RCDSY|Hodgkin's,lymphocyt.dep.NOS|9662/3
C0019829|T191|OP|XE1we|RCDSY|Lymphogranuloma, malignant|9662/3
C0152267|T191|SY|112687003|SNOMEDCT_US|Classical Hodgkin lymphoma, lymphocyte depletion|9662/3
C0019829|T191|SY|118599009|SNOMEDCT_US|HD - Hodgkin's disease|9662/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Hodgkin disease|9662/3
C0152267|T191|SY|118610003|SNOMEDCT_US|Hodgkin disease, lymphocytic depletion|9662/3
C0019829|T191|SY|118602004|SNOMEDCT_US|Hodgkin granuloma|9662/3
C0019829|T191|PT|14537002|SNOMEDCT_US|Hodgkin lymphoma|9662/3
C0152267|T191|PT|112687003|SNOMEDCT_US|Hodgkin lymphoma, lymphocyte depletion|9662/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin lymphoma, no ICD-O subtype|9662/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype|9662/3
C0019829|T191|SY|118606001|SNOMEDCT_US|Hodgkin sarcoma|9662/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Hodgkin's disease|9662/3
C0019829|T191|OAP|154582001|SNOMEDCT_US|Hodgkin's disease|9662/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Hodgkin's disease|9662/3
C0019829|T191|OF|154582001|SNOMEDCT_US|Hodgkin's disease|9662/3
C0019829|T191|OAP|188595005|SNOMEDCT_US|Hodgkin's disease NOS|9662/3
C0019829|T191|OAP|188605006|SNOMEDCT_US|Hodgkin's disease NOS|9662/3
C0019829|T191|OF|188605006|SNOMEDCT_US|Hodgkin's disease NOS|9662/3
C0019829|T191|OAP|188596006|SNOMEDCT_US|Hodgkin's disease NOS, unspecified site|9662/3
C0152267|T191|SY|118610003|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion|9662/3
C0152267|T191|SY|112687003|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion|9662/3
C0152267|T191|OAP|188594009|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion NOS|9662/3
C0152267|T191|IS|112687003|SNOMEDCT_US|Hodgkin's disease, lymphocytic depletion, NOS|9662/3
C0019829|T191|IS|14537002|SNOMEDCT_US|Hodgkin's disease, NOS|9662/3
C0019829|T191|SY|118602004|SNOMEDCT_US|Hodgkin's granuloma|9662/3
C0019829|T191|SY|74189002|SNOMEDCT_US|Hodgkin's granuloma|9662/3
C0019829|T191|OAP|188542007|SNOMEDCT_US|Hodgkin's granuloma NOS|9662/3
C0019829|T191|OAP|188533000|SNOMEDCT_US|Hodgkin's granuloma of unspecified site|9662/3
C0152267|T191|OAP|188584004|SNOMEDCT_US|Hodgkin's lymphocytic depletion of unspecified site|9662/3
C0019829|T191|OAP|52337003|SNOMEDCT_US|Hodgkin's paragranuloma|9662/3
C0019829|T191|OAP|188521005|SNOMEDCT_US|Hodgkin's paragranuloma|9662/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma -RETIRED-|9662/3
C0019829|T191|OF|52337003|SNOMEDCT_US|Hodgkin's paragranuloma -RETIRED-|9662/3
C0019829|T191|OAP|188532005|SNOMEDCT_US|Hodgkin's paragranuloma NOS|9662/3
C0019829|T191|OAP|188522003|SNOMEDCT_US|Hodgkin's paragranuloma of unspecified site|9662/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma, nodular|9662/3
C0019829|T191|IS|52337003|SNOMEDCT_US|Hodgkin's paragranuloma, NOS|9662/3
C0019829|T191|SY|118606001|SNOMEDCT_US|Hodgkin's sarcoma|9662/3
C0019829|T191|SY|46923007|SNOMEDCT_US|Hodgkin's sarcoma|9662/3
C0019829|T191|OAP|188552006|SNOMEDCT_US|Hodgkin's sarcoma NOS|9662/3
C0019829|T191|OAP|188543002|SNOMEDCT_US|Hodgkin's sarcoma of unspecified site|9662/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Lymphoma, Hodgkins|9662/3
C0019829|T191|SY|118599009|SNOMEDCT_US|Malignant Hodgkin's lymphoma|9662/3
C0019829|T191|SY|14537002|SNOMEDCT_US|Malignant lymphoma, Hodgkin's|9662/3
C0152268|T191|PT|0052318|CCPSS|LYMPHOMA HODGKIN NODULAR SCLEROSIS|9663/3
C0152268|T191|PT|0000017244|CHV|nodular sclerosis|9663/3
C0152268|T191|PX|C81.1|ICD10|Hodgkin's disease with nodular sclerosis|9663/3
C0152268|T191|PS|C81.1|ICD10|Nodular sclerosis|9663/3
C0152268|T191|ET|C81.1|ICD10CM|Nodular sclerosis classical Hodgkin lymphoma|9663/3
C0152268|T191|HT|C81.1|ICD10CM|Nodular sclerosis Hodgkin lymphoma|9663/3
C0152268|T191|AB|C81.1|ICD10CM|Nodular sclerosis Hodgkin lymphoma|9663/3
C0152268|T191|HT|201.5|ICD9CM|Hodgkin's disease, nodular sclerosis|9663/3
C0152268|T191|PT|MTHU083131|ICPC2ICD10ENG|disease; Hodgkin's, nodular sclerosis|9663/3
C0152268|T191|PT|MTHU035345|ICPC2ICD10ENG|Hodgkin; nodular sclerosis|9663/3
C0152268|T191|LLT|10020244|MDR|Hodgkin's disease nodular sclerosis|9663/3
C0152268|T191|PT|10020244|MDR|Hodgkin's disease nodular sclerosis|9663/3
C0152268|T191|LLT|10020254|MDR|Hodgkin's disease nodular sclerosis stage unspecified|9663/3
C0152268|T191|LLT|10020299|MDR|Hodgkin's disease, nodular sclerosis|9663/3
C0152268|T191|OL|10029489|MDR|Nodular sclerosis|9663/3
C0152268|T191|PT|31695|MEDCIN|nodular sclerosing Hodgkin's disease|9663/3
C0152268|T191|PN|NOCODE|MTH|Nodular Sclerosis Classical Hodgkin Lymphoma|9663/3
C0152268|T191|ET|201.5|MTHICD9|Hodgkin's disease nodular sclerosis NOS|9663/3
C0152268|T191|SY|C3518|NCI|Hodgkin's Nodular Sclerosis|9663/3
C0152268|T191|PT|C3518|NCI|Nodular Sclerosis Classic Hodgkin Lymphoma|9663/3
C0152268|T191|SY|C3518|NCI|Nodular Sclerosis Classical Hodgkin Lymphoma|9663/3
C0152268|T191|SY|C3518|NCI|Nodular Sclerosis Hodgkin Lymphoma|9663/3
C0152268|T191|SY|C3518|NCI|Nodular Sclerosis Hodgkin's Disease|9663/3
C0152268|T191|SY|C3518|NCI|Nodular Sclerosis Hodgkin's Lymphoma|9663/3
C0152268|T191|AB|C3518|NCI|NSCHL|9663/3
C0152268|T191|AB|C3518|NCI|NSHD|9663/3
C0152268|T191|AB|C3518|NCI|NSHL|9663/3
C0152268|T191|PT|C3518|NCI_CPTAC|Nodular Sclerosis Classic Hodgkin Lymphoma|9663/3
C0152268|T191|DN|C3518|NCI_CTRP|Nodular Sclerosis Classical Hodgkin Lymphoma|9663/3
C0152268|T191|PT|B614.|RCD|Hodgkin's disease, nodular sclerosis|9663/3
C0152268|T191|OP|B614z|RCD|Hodgkin's disease, nodular sclerosis NOS|9663/3
C0152268|T191|OP|B6140|RCD|Hodgkin's disease, nodular sclerosis of unspecified site|9663/3
C0152268|T191|OA|B6140|RCD|Hodgkin's nod.scl. unspec site|9663/3
C0152268|T191|OA|B614z|RCD|Hodgkin's nodular scler. NOS|9663/3
C0152268|T191|AB|B614.|RCD|Hodgkin's nodular sclerosis|9663/3
C0152268|T191|OP|BBj6.|RCDSY|Hodgkin's disease, nodular sclerosis NOS|9663/3
C0152268|T191|OA|BBj6.|RCDSY|Hodgkin's,nodular scler.NOS|9663/3
C0152268|T191|SY|52248008|SNOMEDCT_US|Classical Hodgkin lymphoma, nodular sclerosis|9663/3
C0152268|T191|SY|118608000|SNOMEDCT_US|Hodgkin disease, nodular sclerosis|9663/3
C0152268|T191|PT|52248008|SNOMEDCT_US|Hodgkin lymphoma, nodular sclerosis|9663/3
C0152268|T191|SY|118608000|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis|9663/3
C0152268|T191|OAP|188573006|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis NOS|9663/3
C0152268|T191|OAP|188564003|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis of unspecified site|9663/3
C0152268|T191|IS|52248008|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis, NOS|9663/3
C0334627|T191|PT|MTHU083132|ICPC2ICD10ENG|disease; Hodgkin's, nodular sclerosis, cellular phase|9664/3
C0334627|T191|PT|MTHU035346|ICPC2ICD10ENG|Hodgkin; nodular sclerosis, cellular phase|9664/3
C0334627|T191|PT|91368|MEDCIN|nodular sclerosing Hodgkin's lymphoma in cellular phase|9664/3
C0334627|T191|ET|201.5|MTHICD9|Hodgkin's disease nodular sclerosis cellular phase|9664/3
C0334627|T191|OP|C67171|NCI|Hodgkin's Disease Nodular Sclerosis, Cellular Phase|9664/3
C0334627|T191|PT|C67171|NCI|Nodular Sclerosis Classic Hodgkin Lymphoma, Cellular Phase|9664/3
C0334627|T191|SY|C67171|NCI|Nodular Sclerosis Classical Hodgkin Lymphoma, Cellular Phase|9664/3
C0334627|T191|SY|C67171|NCI|Nodular Sclerosis Hodgkin Lymphoma, Cellular Phase|9664/3
C0334627|T191|AB|XaBBc|RCD|Hodg dis,nod scler,cell phase|9664/3
C0334627|T191|PT|XaBBc|RCD|Hodgkin's disease, nodular sclerosis - cellular phase|9664/3
C0334627|T191|PT|BBj7.|RCDSY|Hodgkin's disease, nodular sclerosis, cellular phase|9664/3
C0334627|T191|AB|BBj7.|RCDSY|Hodgkin's,nod.scler,cellul.|9664/3
C0334627|T191|SY|39086001|SNOMEDCT_US|Classical Hodgkin lymphoma, nodular sclerosis, cellular phase|9664/3
C0334627|T191|SY|307635002|SNOMEDCT_US|Hodgkin disease, nodular sclerosis - cellular phase|9664/3
C0334627|T191|PT|39086001|SNOMEDCT_US|Hodgkin lymphoma, nodular sclerosis, cellular phase|9664/3
C0334627|T191|PT|307635002|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis - cellular phase|9664/3
C0334627|T191|SY|39086001|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis, cellular phase|9664/3
C1521899|T191|PN|NOCODE|MTH|Grade I Nodular Sclerosis Hodgkin's Lymphoma|9665/3
C1521899|T191|PT|C7165|NCI|Grade 1 Nodular Sclerosis Classic Hodgkin Lymphoma|9665/3
C1521899|T191|SY|C7165|NCI|Grade 1 Nodular Sclerosis Classical Hodgkin Lymphoma|9665/3
C1521899|T191|SY|C7165|NCI|Grade 1 Nodular Sclerosis Hodgkin Lymphoma|9665/3
C1521899|T191|SY|C7165|NCI|Grade 1 Nodular Sclerosis Hodgkin's Lymphoma|9665/3
C1521899|T191|SY|C7165|NCI|Grade I Nodular Sclerosis Hodgkin's Lymphoma|9665/3
C1521899|T191|SY|45572000|SNOMEDCT_US|Classical Hodgkin lymphoma, nodular sclerosis, grade 1|9665/3
C1521899|T191|PT|45572000|SNOMEDCT_US|Hodgkin lymphoma, nodular sclerosis, grade 1|9665/3
C0334630|T191|PN|NOCODE|MTH|Grade 2 Nodular Sclerosis Classic Hodgkin Lymphoma|9667/3
C0334630|T191|PT|C7166|NCI|Grade 2 Nodular Sclerosis Classic Hodgkin Lymphoma|9667/3
C0334630|T191|SY|C7166|NCI|Grade 2 Nodular Sclerosis Classical Hodgkin Lymphoma|9667/3
C0334630|T191|SY|C7166|NCI|Grade 2 Nodular Sclerosis Hodgkin Lymphoma|9667/3
C0334630|T191|SY|C7166|NCI|Grade 2 Nodular Sclerosis Hodgkin's Lymphoma|9667/3
C0334630|T191|SY|C7166|NCI|Grade II Nodular Sclerosis Hodgkin's Lymphoma|9667/3
C0334630|T191|SY|43985008|SNOMEDCT_US|Classical Hodgkin lymphoma, nodular sclerosis, grade 2|9667/3
C0334630|T191|PT|43985008|SNOMEDCT_US|Hodgkin lymphoma, nodular sclerosis, grade 2|9667/3
C0334630|T191|SY|43985008|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis, lymphocyte depletion|9667/3
C0334630|T191|SY|43985008|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis, lymphocytic depletion|9667/3
C0334630|T191|SY|43985008|SNOMEDCT_US|Hodgkin's disease, nodular sclerosis, syncytial variant|9667/3
C0855095|T191|SY|0000015228|CHV|diffuse lymphocytic lymphoma|9670/3
C0855095|T191|PT|0000015228|CHV|lymphocytic lymphoma|9670/3
C0855095|T191|SY|0000015228|CHV|lymphoma small lymphocytic|9670/3
C0855095|T191|SY|0000015228|CHV|small lymphocytic lymphoma|9670/3
C0855095|T191|PT|MTHU023064|ICPC2ICD10ENG|diffuse; lymphoma, small cell|9670/3
C0855095|T191|PT|MTHU046693|ICPC2ICD10ENG|lymphocytic; lymphoma, small cell|9670/3
C0855095|T191|PT|MTHU046758|ICPC2ICD10ENG|lymphoma; diffuse, small cell|9670/3
C0855095|T191|PT|MTHU046816|ICPC2ICD10ENG|lymphoma; lymphocytic, small cell|9670/3
C0855095|T191|LLT|10003908|MDR|B-cell small lymphocytic lymphoma|9670/3
C0855095|T191|PT|10003908|MDR|B-cell small lymphocytic lymphoma|9670/3
C0855095|T191|LLT|10003910|MDR|B-cell small lymphocytic lymphoma NOS|9670/3
C0855095|T191|HT|10003909|MDR|B-cell small lymphocytic lymphomas|9670/3
C0855095|T191|LLT|10051812|MDR|Small cell lymphocytic lymphoma|9670/3
C0855095|T191|SY|335985|MEDCIN|malignant neoplasm lymphoma small b-cell lymphocytic|9670/3
C0855095|T191|PT|335985|MEDCIN|small B-cell lymphocytic lymphoma|9670/3
C0855095|T191|PN|NOCODE|MTH|Small Lymphocytic Lymphoma|9670/3
C0855095|T191|ET|200.1|MTHICD9|Diffuse lymphocytic lymphoma|9670/3
C0855095|T191|ET|200.1|MTHICD9|Diffuse lymphocytic lymphosarcoma|9670/3
C0855095|T191|ET|200.1|MTHICD9|Diffuse lymphocytic malignant lymphoma|9670/3
C0855095|T191|ET|200.1|MTHICD9|Lymphocytic lymphosarcoma|9670/3
C0855095|T191|SY|C7540|NCI|B-Cell Small Lymphocytic Lymphoma|9670/3
C0855095|T191|OP|C7540|NCI|Diffuse Well Differentiated Lymphocytic Lymphoma|9670/3
C0855095|T191|AB|C7540|NCI|SLL|9670/3
C0855095|T191|SY|C7540|NCI|Small B-Cell Lymphocytic Lymphoma|9670/3
C0855095|T191|PT|C7540|NCI|Small Lymphocytic Lymphoma|9670/3
C0855095|T191|SY|C7540|NCI_CDISC|B-Cell Small Lymphocytic Lymphoma|9670/3
C0855095|T191|SY|C7540|NCI_CDISC|Lymphoma, Lymphocytic, Malignant|9670/3
C0855095|T191|PT|C7540|NCI_CDISC|LYMPHOMA, SMALL LYMPHOCYTIC, MALIGNANT|9670/3
C0855095|T191|SY|C7540|NCI_CDISC|SLL|9670/3
C0855095|T191|SY|C7540|NCI_CDISC|Small B-Cell Lymphocytic Lymphoma|9670/3
C0855095|T191|PT|C7540|NCI_CPTAC|Small Lymphocytic Lymphoma|9670/3
C0855095|T191|PT|10003910|NCI_CTEP-SDC|Small lymphocytic lymphoma, NOS|9670/3
C0855095|T191|DN|C7540|NCI_CTRP|Small Lymphocytic Lymphoma|9670/3
C0855095|T191|PT|CDR0000641299|NCI_NCI-GLOSS|SLL|9670/3
C0855095|T191|PT|CDR0000407751|NCI_NCI-GLOSS|small lymphocytic lymphoma|9670/3
C0855095|T191|PT|CDR0000415910|NCI_NCI-GLOSS|well-differentiated lymphocytic lymphoma|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|B-Cell Small Lymphocytic Lymphoma|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|diffuse lymphocytic, well-differentiated lymphoma|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|diffuse WDL lymphoma|9670/3
C0855095|T191|IS|CDR0000038170|PDQ|Diffuse Well Differentiated Lymphocytic Lymphoma|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|diffuse well-differentiated lymphocytic lymphoma|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|DLWD lymphoma|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|DWDL lymphoma|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|lymphocytic lymphoma, small|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|lymphoma, diffuse lymphocytic, well-differentiated|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|lymphoma, small lymphocytic|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|SL lymphoma|9670/3
C0855095|T191|AB|CDR0000038170|PDQ|SLL|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|Small B-Cell Lymphocytic Lymphoma|9670/3
C0855095|T191|PT|CDR0000038170|PDQ|small lymphocytic lymphoma|9670/3
C0855095|T191|ET|CDR0000038170|PDQ|Small lymphocytic lymphoma|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|WDL, diffuse lymphocytic|9670/3
C0855095|T191|SY|CDR0000038170|PDQ|well-differentiated lymphoma, diffuse lymphocytic|9670/3
C0855095|T191|SY|Xa99l|RCD|Lymphocytic lymphoma|9670/3
C0855095|T191|SY|Xa99l|RCD|Lymphocytic lymphosarcoma|9670/3
C0855095|T191|AB|Xa99l|RCD|M lymphoma,lymphocyt,well dif|9670/3
C0855095|T191|AB|Xa99l|RCD|Malign lymph-small lymphocytic|9670/3
C0855095|T191|SY|Xa99l|RCD|Malignant lymphoma - small cell|9670/3
C0855095|T191|PT|Xa99l|RCD|Malignant lymphoma - small lymphocytic|9670/3
C0855095|T191|AB|Xa99l|RCD|Malignant lymphoma-small cell|9670/3
C0855095|T191|SY|Xa99l|RCD|Malignant lymphoma, lymphocytic, well differentiated|9670/3
C0855095|T191|IS|BBgC.|RCDSY|Lymphocytic lymphoma NOS|9670/3
C0855095|T191|OA|BBgC.|RCDSY|Lymphocytic lymphosarc NOS|9670/3
C0855095|T191|IS|BBgC.|RCDSY|Lymphocytic lymphosarcoma NOS|9670/3
C0855095|T191|OA|BBgC.|RCDSY|Malig.lymph,ly-cyt,well NOS|9670/3
C0855095|T191|OA|BBgL.|RCDSY|Malign lymph,small lymphocy|9670/3
C0855095|T191|OP|BBgC.|RCDSY|Malignant lymphoma, lymphocytic, well differentiated NOS|9670/3
C0855095|T191|OP|BBgL.|RCDSY|Malignant lymphoma, small lymphocytic NOS|9670/3
C0855095|T191|SY|302841002|SNOMEDCT_US|Lymphocytic lymphoma|9670/3
C0855095|T191|SY|302841002|SNOMEDCT_US|Lymphocytic lymphosarcoma|9670/3
C0855095|T191|SY|302841002|SNOMEDCT_US|Malignant lymphoma - small cell|9670/3
C0855095|T191|PT|302841002|SNOMEDCT_US|Malignant lymphoma - small lymphocytic|9670/3
C0855095|T191|SY|64575004|SNOMEDCT_US|Malignant lymphoma, lymphocytic|9670/3
C0855095|T191|SY|64575004|SNOMEDCT_US|Malignant lymphoma, lymphocytic, diffuse|9670/3
C0855095|T191|IS|64575004|SNOMEDCT_US|Malignant lymphoma, lymphocytic, diffuse, NOS|9670/3
C0855095|T191|IS|64575004|SNOMEDCT_US|Malignant lymphoma, lymphocytic, NOS|9670/3
C0855095|T191|SY|302841002|SNOMEDCT_US|Malignant lymphoma, lymphocytic, well differentiated|9670/3
C0855095|T191|SY|64575004|SNOMEDCT_US|Malignant lymphoma, lymphocytic, well differentiated, diffuse|9670/3
C0855095|T191|SY|64575004|SNOMEDCT_US|Malignant lymphoma, small B lymphocytic|9670/3
C0855095|T191|SY|64575004|SNOMEDCT_US|Malignant lymphoma, small cell|9670/3
C0855095|T191|SY|64575004|SNOMEDCT_US|Malignant lymphoma, small cell diffuse|9670/3
C0855095|T191|IS|64575004|SNOMEDCT_US|Malignant lymphoma, small cell, diffuse, NOS|9670/3
C0855095|T191|IS|64575004|SNOMEDCT_US|Malignant lymphoma, small cell, NOS|9670/3
C0855095|T191|PT|64575004|SNOMEDCT_US|Malignant lymphoma, small lymphocytic|9670/3
C0855095|T191|SY|64575004|SNOMEDCT_US|Malignant lymphoma, small lymphocytic, diffuse|9670/3
C0855095|T191|IS|64575004|SNOMEDCT_US|Malignant lymphoma, small lymphocytic, NOS|9670/3
C0855095|T191|SY|302841002|SNOMEDCT_US|Small lymphocytic lymphoma|9670/3
C0334633|T191|PT|0000030014|CHV|immunocytoma|9671/3
C0334633|T191|ET|C83.0|ICD10CM|Lymphoplasmacytic lymphoma|9671/3
C0334633|T191|PT|MTHU037619|ICPC2ICD10ENG|immunocytoma|9671/3
C0334633|T191|PT|MTHU046823|ICPC2ICD10ENG|lymphoma; lymphoplasmacytoid|9671/3
C0334633|T191|PT|MTHU046851|ICPC2ICD10ENG|lymphoma; plasmacytic|9671/3
C0334633|T191|PT|MTHU046868|ICPC2ICD10ENG|lymphoplasmacytoid; lymphoma|9671/3
C0334633|T191|PT|MTHU059930|ICPC2ICD10ENG|plasmacytic; lymphoma|9671/3
C0334633|T191|PT|355928|MEDCIN|malignant lymphoplasmacytic lymphoma|9671/3
C0334633|T191|SY|355928|MEDCIN|malignant neoplasm lymphoma lymphoplasmacytic|9671/3
C0334633|T191|PN|NOCODE|MTH|Malignant lymphoma - lymphoplasmacytic|9671/3
C0334633|T191|ET|200.8|MTHICD9|Malignant lymphoplasmacytoid type lymphoma|9671/3
C0334633|T191|OP|C3212|NCI|Immunocytoma, Lymphoplasmacytic Type|9671/3
C0334633|T191|PT|C3212|NCI|Lymphoplasmacytic Lymphoma|9671/3
C0334633|T191|SY|TCGA|NCI|Lymphoplasmacytic Lymphoma|9671/3
C0334633|T191|SY|C3212|NCI|Lymphoplasmacytoid Lymphoma|9671/3
C0334633|T191|SY|C3212|NCI_CDISC|Immunocytoma, Lymphoplasmacytic Type|9671/3
C0334633|T191|PT|C3212|NCI_CDISC|LYMPHOMA, LYMPHOPLASMACYTIC, MALIGNANT|9671/3
C0334633|T191|SY|C3212|NCI_CDISC|Lymphoma, Plasmacytic|9671/3
C0334633|T191|SY|C3212|NCI_CDISC|Lymphoplasmacytoid Lymphoma|9671/3
C0334633|T191|SY|10047803|NCI_CTEP-SDC|Lymphoplasmacytic lymphoma|9671/3
C0334633|T191|DN|C3212|NCI_CTRP|Lymphoplasmacytic Lymphoma|9671/3
C0334633|T191|PT|CDR0000409750|NCI_NCI-GLOSS|lymphoplasmacytic lymphoma|9671/3
C0334633|T191|SY|XaBBN|RCD|Immunocytoma|9671/3
C0334633|T191|AB|XaBBN|RCD|Mal lymphoma, lymphoplasmacyt|9671/3
C0334633|T191|AB|XaBBN|RCD|Malignant lymph-lymphoplasmac|9671/3
C0334633|T191|PT|XaBBN|RCD|Malignant lymphoma - lymphoplasmacytic|9671/3
C0334633|T191|SY|XaBBN|RCD|Malignant lymphoma, lymphoplasmacytoid type|9671/3
C0334633|T191|SY|XaBBN|RCD|Plasmacytic lymphoma|9671/3
C0334633|T191|AB|BBg7.|RCDSY|Malig.lymph,lymphoplasmacyt|9671/3
C0334633|T191|PT|BBg7.|RCDSY|Malignant lymphoma, lymphoplasmacytoid type|9671/3
C0334633|T191|SY|19340000|SNOMEDCT_US|Immunocytoma|9671/3
C0334633|T191|SY|307623001|SNOMEDCT_US|Immunocytoma|9671/3
C0334633|T191|PT|307623001|SNOMEDCT_US|Malignant lymphoma - lymphoplasmacytic|9671/3
C0334633|T191|PT|19340000|SNOMEDCT_US|Malignant lymphoma, lymphoplasmacytic|9671/3
C0334633|T191|SY|19340000|SNOMEDCT_US|Malignant lymphoma, lymphoplasmacytoid|9671/3
C0334633|T191|SY|307623001|SNOMEDCT_US|Malignant lymphoma, lymphoplasmacytoid type|9671/3
C0334633|T191|SY|19340000|SNOMEDCT_US|Malignant lymphoma, plasmacytoid|9671/3
C0334633|T191|SY|307623001|SNOMEDCT_US|Plasmacytic lymphoma|9671/3
C0334633|T191|SY|19340000|SNOMEDCT_US|Plasmacytic lymphoma|9671/3
C4721414|T191|SY|0000030015|CHV|cell lymphoma mantle|9673/3
C4721414|T191|PT|0000030015|CHV|mantle cell lymphoma|9673/3
C4721414|T191|SY|0000030015|CHV|mantle cell lymphomas|9673/3
C4721414|T191|SY|0000030015|CHV|mantle-cell lymphoma|9673/3
C4721414|T191|HT|C83.1|ICD10CM|Mantle cell lymphoma|9673/3
C4721414|T191|AB|C83.1|ICD10CM|Mantle cell lymphoma|9673/3
C4721414|T191|HT|200.4|ICD9CM|Mantle cell lymphoma|9673/3
C0334634|T191|PT|MTHU023070|ICPC2ICD10ENG|diffuse; lymphoma, lymphocytic, poorly differentiated|9673/3
C0334634|T191|PT|MTHU046764|ICPC2ICD10ENG|lymphoma; diffuse, lymphocytic, poorly differentiated|9673/3
C4721414|T191|PT|MTHU046825|ICPC2ICD10ENG|lymphoma; mantle zone|9673/3
C4721414|T191|PT|MTHU047542|ICPC2ICD10ENG|mantle zone; lymphoma|9673/3
C4721414|T191|LA|LA26524-1|LNC|Mantle cell lymphoma|9673/3
C4721414|T191|PT|10061275|MDR|Mantle cell lymphoma|9673/3
C4721414|T191|LLT|10061275|MDR|Mantle cell lymphoma|9673/3
C4721414|T191|LLT|10026799|MDR|Mantle cell lymphoma NOS|9673/3
C4721414|T191|HT|10026798|MDR|Mantle cell lymphomas|9673/3
C4721414|T191|LLT|10026806|MDR|Mantle zone lymphoma|9673/3
C4721414|T191|PT|312883|MEDCIN|mantle cell lymphoma|9673/3
C0334634|T191|PM|D020522|MSH|Centrocytic Small-Cell Lymphoma|9673/3
C0334634|T191|PM|D020522|MSH|Centrocytic Small-Cell Lymphomas|9673/3
C0334634|T191|DEV|D020522|MSH|DIFFUSE LYMPHOCYTIC LYMPHOMA POORLY DIFFER|9673/3
C0334634|T191|PM|D020522|MSH|Diffuse Lymphocytic Lymphoma, Poorly Differentiated|9673/3
C0334634|T191|ET|D020522|MSH|Diffuse Lymphocytic Lymphoma, Poorly-Differentiated|9673/3
C0334634|T191|DEV|D020522|MSH|LYMPHOCYTIC LYMPHOMA DIFFUSE POORLY DIFFER|9673/3
C0334634|T191|ET|D020522|MSH|Lymphocytic Lymphoma, Diffuse, Poorly Differentiated|9673/3
C0334634|T191|ET|D020522|MSH|Lymphocytic Lymphoma, Diffuse, Poorly-Differentiated|9673/3
C0334634|T191|DEV|D020522|MSH|LYMPHOMA LYMPHOCYTIC DIFFUSE INTERMEDIATE DIFFER|9673/3
C0334634|T191|DEV|D020522|MSH|LYMPHOMA LYMPHOCYTIC DIFFUSE POORLY DIFFER|9673/3
C0334634|T191|PM|D020522|MSH|Lymphoma, Centrocytic Small Cell|9673/3
C0334634|T191|ET|D020522|MSH|Lymphoma, Centrocytic Small-Cell|9673/3
C0334634|T191|ET|D020522|MSH|Lymphoma, Lymphocytic, Diffuse, Intermediate Differentiated|9673/3
C0334634|T191|ET|D020522|MSH|Lymphoma, Lymphocytic, Diffuse, Poorly-Differentiated|9673/3
C0334634|T191|PM|D020522|MSH|Lymphoma, Mantle Cell|9673/3
C0334634|T191|MH|D020522|MSH|Lymphoma, Mantle-Cell|9673/3
C0334634|T191|PM|D020522|MSH|Lymphoma, Mantle-Zone|9673/3
C0334634|T191|ET|D020522|MSH|Lymphoma, Small-Cell, Centrocytic|9673/3
C0334634|T191|PM|D020522|MSH|Lymphomas, Centrocytic Small-Cell|9673/3
C0334634|T191|PM|D020522|MSH|Lymphomas, Mantle-Cell|9673/3
C0334634|T191|PM|D020522|MSH|Lymphomas, Mantle-Zone|9673/3
C0334634|T191|PM|D020522|MSH|Mantle Cell Lymphoma|9673/3
C0334634|T191|PM|D020522|MSH|Mantle Zone Lymphoma|9673/3
C0334634|T191|ET|D020522|MSH|Mantle-Cell Lymphoma|9673/3
C0334634|T191|PM|D020522|MSH|Mantle-Cell Lymphomas|9673/3
C0334634|T191|ET|D020522|MSH|Mantle-Zone Lymphoma|9673/3
C0334634|T191|PM|D020522|MSH|Mantle-Zone Lymphomas|9673/3
C0334634|T191|PM|D020522|MSH|Small-Cell Lymphoma, Centrocytic|9673/3
C0334634|T191|PM|D020522|MSH|Small-Cell Lymphomas, Centrocytic|9673/3
C0334634|T191|PN|NOCODE|MTH|Malignant lymphoma, lymphocytic, intermediate differentiation, diffuse|9673/3
C4721414|T191|PN|NOCODE|MTH|Mantle cell lymphoma|9673/3
C4721414|T191|SY|C4337|NCI|Classical Mantle Cell Lymphoma|9673/3
C4721414|T191|PT|C4337|NCI|Mantle Cell Lymphoma|9673/3
C4721414|T191|SY|TCGA|NCI|Mantle Cell Lymphoma|9673/3
C4721414|T191|SY|C4337|NCI|Mantle Zone Lymphoma|9673/3
C4721414|T191|AB|C4337|NCI|MCL|9673/3
C4721414|T191|PT|C4337|NCI_CPTAC|Mantle Cell Lymphoma|9673/3
C4721414|T191|PT|10026799|NCI_CTEP-SDC|Mantle cell lymphoma|9673/3
C4721414|T191|DN|C4337|NCI_CTRP|Mantle Cell Lymphoma|9673/3
C4721414|T191|PT|CDR0000445048|NCI_NCI-GLOSS|mantle cell lymphoma|9673/3
C0334634|T191|SY|CDR0000038370|PDQ|diffuse PDL lymphoma|9673/3
C0334634|T191|SY|CDR0000038370|PDQ|diffuse poorly-differentiated lymphocytic lymphoma|9673/3
C0334634|T191|SY|CDR0000038370|PDQ|DPDL lymphoma|9673/3
C4721414|T191|SY|CDR0000042534|PDQ|lymphoma, mantle cell|9673/3
C4721414|T191|PT|CDR0000042534|PDQ|mantle cell lymphoma|9673/3
C4721414|T191|SY|CDR0000042534|PDQ|Mantle Zone Lymphoma|9673/3
C4721414|T191|AB|CDR0000042534|PDQ|MCL|9673/3
C0334634|T191|OA|BBgN.|RCDSY|Malg lymph,lym,int difn,dif|9673/3
C0334634|T191|OA|BBgN.|RCDSY|Malign lymphoma,lymphocytic,intermediate differn, diffuse|9673/3
C0334634|T191|OP|BBgN.|RCDSY|Malignant lymphoma, lymphocytic, intermediate differentiation, diffuse|9673/3
C0334634|T191|IS|74654000|SNOMEDCT_US|Malignant lymphoma, lymphocytic, intermediate differentiation, diffuse|9673/3
C0334634|T191|IS|63086004|SNOMEDCT_US|Malignant lymphoma, lymphocytic, poorly differentiated, diffuse|9673/3
C0334634|T191|PT|74654000|SNOMEDCT_US|Mantle cell lymphoma|9673/3
C4721414|T191|PT|443487006|SNOMEDCT_US|Mantle cell lymphoma|9673/3
C0334634|T191|IS|74654000|SNOMEDCT_US|Mantle zone lymphoma|9673/3
C0079757|T191|PT|MTHU023058|ICPC2ICD10ENG|diffuse; lymphoma, mixed cell type|9675/3
C0079757|T191|PT|MTHU023059|ICPC2ICD10ENG|diffuse; lymphoma, mixed cell type, small and large cell|9675/3
C0079757|T191|PT|MTHU046752|ICPC2ICD10ENG|lymphoma; diffuse, mixed cell type|9675/3
C0079757|T191|PT|MTHU046753|ICPC2ICD10ENG|lymphoma; diffuse, mixed cell type, small and large cell|9675/3
C0079757|T191|PT|MTHU046789|ICPC2ICD10ENG|lymphoma; mixed cell type, diffuse|9675/3
C0079757|T191|PM|D008228|MSH|Diffuse Mixed Cell Lymphoma|9675/3
C0079757|T191|DEV|D008228|MSH|DIFFUSE MIXED LYMPHOMA|9675/3
C0079757|T191|ET|D008228|MSH|Diffuse Mixed Small and Large Cell Lymphoma|9675/3
C0079757|T191|DEV|D008228|MSH|DIFFUSE MIXED SMALL LARGE LYMPHOMA|9675/3
C0079757|T191|ET|D008228|MSH|Diffuse Mixed-Cell Lymphoma|9675/3
C0079757|T191|PM|D008228|MSH|Diffuse Mixed-Cell Lymphomas|9675/3
C0079757|T191|DEV|D008228|MSH|LYMPHOMA DIFFUSE MIXED LYMPHOCYTIC HISTIOCYTIC|9675/3
C0079757|T191|DEV|D008228|MSH|LYMPHOMA MIXED DIFFUSE|9675/3
C0079757|T191|DEV|D008228|MSH|LYMPHOMA MIXED SMALL LARGE DIFFUSE|9675/3
C0079757|T191|DEV|D008228|MSH|LYMPHOMA SMALL LARGE CLEAVED DIFFUSE|9675/3
C0079757|T191|PM|D008228|MSH|Lymphoma, Diffuse Mixed-Cell|9675/3
C0079757|T191|ET|D008228|MSH|Lymphoma, Diffuse, Mixed Lymphocytic-Histiocytic|9675/3
C0079757|T191|ET|D008228|MSH|Lymphoma, Mixed Cell, Diffuse|9675/3
C0079757|T191|ET|D008228|MSH|Lymphoma, Mixed Small and Large Cell, Diffuse|9675/3
C0079757|T191|PEP|D008228|MSH|Lymphoma, Mixed-Cell, Diffuse|9675/3
C0079757|T191|ET|D008228|MSH|Lymphoma, Small and Large Cleaved-Cell, Diffuse|9675/3
C0079757|T191|PM|D008228|MSH|Mixed Cell Lymphoma, Diffuse|9675/3
C0079757|T191|DEV|D008228|MSH|MIXED LYMPHOMA DIFFUSE|9675/3
C0079757|T191|ET|D008228|MSH|Mixed Small and Large Cell Lymphoma, Diffuse|9675/3
C0079757|T191|DEV|D008228|MSH|MIXED SMALL LARGE LYMPHOMA DIFFUSE|9675/3
C0079757|T191|ET|D008228|MSH|Mixed-Cell Lymphoma, Diffuse|9675/3
C0079757|T191|PN|NOCODE|MTH|Diffuse Mixed-Cell Lymphoma|9675/3
C0334636|T191|ET|200.8|MTHICD9|Diffuse mixed cell type lymphosarcoma|9675/3
C0079757|T191|ET|200.8|MTHICD9|Diffuse mixed lymphocytic-histiocytic lymphoma|9675/3
C0334636|T191|ET|200.8|MTHICD9|Diffuse mixed lymphocytic-histiocytic malignant lymphoma|9675/3
C0079757|T191|PT|C3463|NCI|Diffuse Mixed Cell Lymphoma|9675/3
C0079757|T191|OP|C3463|NCI|Diffuse Mixed Cell Lymphoma|9675/3
C0079757|T191|OP|C3463|NCI|Diffuse Mixed Large and Small Cell Lymphoma|9675/3
C0334636|T191|OA|BBgP.|RCDSY|Malig lymph,small+larg,diff|9675/3
C0334636|T191|OP|BBgP.|RCDSY|Malignant lymphoma, mixed small and large cell, diffuse|9675/3
C0334636|T191|SY|50102004|SNOMEDCT_US|Malignant lymphoma, mixed cell type, diffuse|9675/3
C0334636|T191|SY|50102004|SNOMEDCT_US|Malignant lymphoma, mixed lymphocytic-histiocytic, diffuse|9675/3
C0334636|T191|PT|50102004|SNOMEDCT_US|Malignant lymphoma, mixed small and large cell, diffuse|9675/3
C1292753|T191|ET|C83.8|ICD10CM|Primary effusion B-cell lymphoma|9678/3
C1292753|T191|PT|10065857|MDR|Primary effusion lymphoma|9678/3
C1292753|T191|LLT|10065857|MDR|Primary effusion lymphoma|9678/3
C1292753|T191|SY|366463|MEDCIN|b-cell primary effusion lymphoma|9678/3
C1292753|T191|PT|366463|MEDCIN|Primary effusion lymphoma|9678/3
C1292753|T191|PM|D054685|MSH|Effusion Lymphoma, Primary|9678/3
C1292753|T191|PM|D054685|MSH|Effusion Lymphomas, Primary|9678/3
C1292753|T191|MH|D054685|MSH|Lymphoma, Primary Effusion|9678/3
C1292753|T191|PM|D054685|MSH|Lymphomas, Primary Effusion|9678/3
C1292753|T191|ET|D054685|MSH|Primary Effusion Lymphoma|9678/3
C1292753|T191|PM|D054685|MSH|Primary Effusion Lymphomas|9678/3
C1292753|T191|PN|NOCODE|MTH|Primary Effusion Lymphoma|9678/3
C1292753|T191|AB|C6915|NCI|PEL|9678/3
C1292753|T191|SY|TCGA|NCI|Primary Effusion Lymphoma|9678/3
C1292753|T191|PT|C6915|NCI|Primary Effusion Lymphoma|9678/3
C1292753|T191|PT|10065857|NCI_CTEP-SDC|Primary effusion lymphoma|9678/3
C1292753|T191|DN|C6915|NCI_CTRP|Primary Effusion Lymphoma|9678/3
C1292753|T191|PT|CDR0000455144|NCI_NCI-GLOSS|primary effusion lymphoma|9678/3
C1292753|T191|PT|713516007|SNOMEDCT_US|Primary effusion lymphoma|9678/3
C1292753|T191|IS|128800006|SNOMEDCT_US|Primary effusion lymphoma|9678/3
C1292753|T191|PT|128800006|SNOMEDCT_US|Primary effusion lymphoma|9678/3
C1292754|T191|CN|MTHU063569|LNC|Primary mediastinal large B-cell lymphoma|9679/3
C1292754|T191|LPN|LP411612-7|LNC|Primary mediastinal large B-cell lymphoma|9679/3
C1292754|T191|LLT|10036710|MDR|Primary mediastinal large B-cell lymphoma|9679/3
C1292754|T191|PT|10036710|MDR|Primary mediastinal large B-cell lymphoma|9679/3
C1292754|T191|LLT|10036712|MDR|Primary mediastinal large B-cell lymphoma NOS|9679/3
C1292754|T191|HT|10036711|MDR|Primary mediastinal large B-cell lymphomas|9679/3
C1292754|T191|PT|339510|MEDCIN|primary malignant mediastinal large b-cell lymphoma of thymus|9679/3
C1292754|T191|SY|339510|MEDCIN|thymus malignant lymphoma mediastinal large b-cell primary|9679/3
C1292754|T191|SY|C9280|NCI|B-Cell Diffuse Large Cell Lymphoma of Mediastinum|9679/3
C1292754|T191|SY|C9280|NCI|B-Cell Diffuse Large Cell Lymphoma of the Mediastinum|9679/3
C1292754|T191|SY|C9280|NCI|Mediastinal B-Cell Diffuse Large Cell Lymphoma|9679/3
C1292754|T191|OP|C9280|NCI|Mediastinal Diffuse Large Cell Lymphoma with Sclerosis|9679/3
C1292754|T191|AB|C9280|NCI|PMBL|9679/3
C1292754|T191|AB|C9280|NCI|PMLCL|9679/3
C1292754|T191|OP|C9280|NCI|Primary Mediastinal Clear Cell Lymphoma of B-Cell Type|9679/3
C1292754|T191|SY|C9280|NCI|Primary Mediastinal Large B-Cell Lymphoma|9679/3
C1292754|T191|SY|10036712|NCI_CTEP-SDC|Mediastinal large B-cell lymphoma|9679/3
C1292754|T191|SY|CDR0000771634|PDQ|B-cell diffuse large cell lymphoma of mediastinum|9679/3
C1292754|T191|SY|CDR0000771634|PDQ|B-cell diffuse large cell lymphoma of the mediastinum|9679/3
C1292754|T191|SY|CDR0000771634|PDQ|mediastinal B-cell diffuse large cell lymphoma|9679/3
C1292754|T191|AB|CDR0000771634|PDQ|PMBL|9679/3
C1292754|T191|AB|CDR0000771634|PDQ|PMLCL|9679/3
C1292754|T191|SY|CDR0000771634|PDQ|primary mediastinal large B-cell lymphoma|9679/3
C1292754|T191|PT|128801005|SNOMEDCT_US|Mediastinal large B-cell lymphoma|9679/3
C1292754|T191|SY|128801005|SNOMEDCT_US|Thymic large B-cell lymphoma|9679/3
C0079744|T191|SY|0000015222|CHV|diffuse histiocytic lymphoma|9680/3
C0079744|T191|SY|0000030016|CHV|diffuse large b cell lymphoma|9680/3
C0079744|T191|PT|0000030016|CHV|diffuse large b-cell lymphoma|9680/3
C0079744|T191|PT|0000015222|CHV|diffuse large cell lymphoma|9680/3
C0079744|T191|SY|0000015222|CHV|large cell diffuse lymphoma|9680/3
C0079744|T191|HT|C83.3|ICD10CM|Diffuse large B-cell lymphoma|9680/3
C0079744|T191|AB|C83.3|ICD10CM|Diffuse large B-cell lymphoma|9680/3
C0079744|T191|PT|MTHU023063|ICPC2ICD10ENG|diffuse; lymphoma, histiocytic|9680/3
C0079744|T191|PT|MTHU023061|ICPC2ICD10ENG|diffuse; lymphoma, large cell|9680/3
C0079744|T191|PT|MTHU046757|ICPC2ICD10ENG|lymphoma; diffuse, histiocytic|9680/3
C0079744|T191|PT|MTHU046755|ICPC2ICD10ENG|lymphoma; diffuse, large cell|9680/3
C2698294|T191|LA|LA26527-4|LNC|B-cell lymphoma, unclassifiable, with features intermediate between diffuse large B-cell lymphoma and Burkitt lymphoma|9680/3
C0079744|T191|LPN|LP411613-5|LNC|Diffuse large B-cell lymphoma|9680/3
C5192818|T191|CN|MTHU063570|LNC|Diffuse large B-cell lymphoma.activated B-cell subtype|9680/3
C5192818|T191|LPN|LP411618-4|LNC|Diffuse large B-cell lymphoma.activated B-cell subtype|9680/3
C0079744|T191|LLT|10012818|MDR|Diffuse large B-cell lymphoma|9680/3
C0079744|T191|PT|10012818|MDR|Diffuse large B-cell lymphoma|9680/3
C0079744|T191|LLT|10012820|MDR|Diffuse large B-cell lymphoma NOS|9680/3
C0079744|T191|HT|10012819|MDR|Diffuse large B-cell lymphomas|9680/3
C1321547|T191|LLT|10080211|MDR|T-cell/histiocyte-rich large B-cell lymphoma|9680/3
C2698294|T191|PT|366685|MEDCIN|B-cell lymphoma unclassifiable with features intermediate between Burkitt lymphoma and diffuse large B-cell lymphoma|9680/3
C0079744|T191|SY|31689|MEDCIN|DHL|9680/3
C2700007|T191|PT|366462|MEDCIN|Epstein-Barr virus positive diffuse large B-cell lymphoma of elderly|9680/3
C2026186|T191|PT|236170|MEDCIN|large B-cell diffuse lymphoma of central nervous system|9680/3
C0079744|T191|PM|D016403|MSH|Diffuse Histiocytic Lymphoma|9680/3
C0079744|T191|PM|D016403|MSH|Diffuse Histiocytic Lymphomas|9680/3
C0079744|T191|PM|D016403|MSH|Diffuse Large Cell Lymphoma|9680/3
C0079744|T191|DEV|D016403|MSH|DIFFUSE LARGE LYMPHOMA|9680/3
C0079744|T191|ET|D016403|MSH|Diffuse Large-Cell Lymphoma|9680/3
C0079744|T191|PM|D016403|MSH|Diffuse Large-Cell Lymphomas|9680/3
C0079744|T191|ET|D016403|MSH|Diffuse, Large B-Cell, Lymphoma|9680/3
C0079744|T191|ET|D016403|MSH|Histiocytic Lymphoma|9680/3
C0079744|T191|ET|D016403|MSH|Histiocytic Lymphoma, Diffuse|9680/3
C0079744|T191|PM|D016403|MSH|Histiocytic Lymphomas|9680/3
C0079744|T191|PM|D016403|MSH|Histiocytic Lymphomas, Diffuse|9680/3
C0079744|T191|PM|D016403|MSH|Large Cell Lymphoma, Diffuse|9680/3
C0079744|T191|ET|D016403|MSH|Large Lymphoid Lymphoma, Diffuse|9680/3
C0079744|T191|DEV|D016403|MSH|LARGE LYMPHOMA DIFFUSE|9680/3
C0079744|T191|ET|D016403|MSH|Large-Cell Lymphoma, Diffuse|9680/3
C0079744|T191|PM|D016403|MSH|Large-Cell Lymphomas, Diffuse|9680/3
C0079744|T191|DEV|D016403|MSH|LYMPHOMA DIFFUSE LARGE|9680/3
C0079744|T191|DEV|D016403|MSH|LYMPHOMA LARGE DIFFUSE|9680/3
C0079744|T191|PM|D016403|MSH|Lymphoma, Diffuse Histiocytic|9680/3
C0079744|T191|PM|D016403|MSH|Lymphoma, Diffuse Large Cell|9680/3
C0079744|T191|ET|D016403|MSH|Lymphoma, Diffuse Large-Cell|9680/3
C0079744|T191|ET|D016403|MSH|Lymphoma, Histiocytic|9680/3
C0079744|T191|ET|D016403|MSH|Lymphoma, Histiocytic, Diffuse|9680/3
C0079744|T191|MH|D016403|MSH|Lymphoma, Large B-Cell, Diffuse|9680/3
C0079744|T191|ET|D016403|MSH|Lymphoma, Large Cell, Diffuse|9680/3
C0079744|T191|ET|D016403|MSH|Lymphoma, Large Lymphoid, Diffuse|9680/3
C0079744|T191|ET|D016403|MSH|Lymphoma, Large-Cell, Diffuse|9680/3
C0079744|T191|PM|D016403|MSH|Lymphomas, Diffuse Histiocytic|9680/3
C0079744|T191|PM|D016403|MSH|Lymphomas, Diffuse Large-Cell|9680/3
C0079744|T191|PM|D016403|MSH|Lymphomas, Histiocytic|9680/3
C0079744|T191|PN|NOCODE|MTH|Diffuse Large B-Cell Lymphoma|9680/3
C2698294|T191|PN|NOCODE|MTH|High Grade B-Cell Lymphoma, Not Otherwise Specified|9680/3
C2700007|T191|OP|C80281|NCI|Age-Related EBV Positive B-Cell Lymphoproliferative Disorder|9680/3
C2698294|T191|OP|C80291|NCI|B-Cell Lymphoma, Unclassifiable, with Features Intermediate between Diffuse Large B-Cell Lymphoma and Burkitt Lymphoma|9680/3
C2698294|T191|AB|C80291|NCI|BCLU|9680/3
C2026186|T191|SY|C71720|NCI|Central Nervous System Diffuse Large B-Cell Lymphoma|9680/3
C2026186|T191|AB|C71720|NCI|CNS DLBCL|9680/3
C0079744|T191|SY|TCGA|NCI|Diffuse Large B-Cell Lymphoma|9680/3
C0079744|T191|PT|C8851|NCI|Diffuse Large B-Cell Lymphoma|9680/3
C2699776|T191|PT|C80289|NCI|Diffuse Large B-Cell Lymphoma Associated with Chronic Inflammation|9680/3
C0079744|T191|AB|C8851|NCI|DLBCL|9680/3
C2699776|T191|AB|C80289|NCI|DLBCL-CI|9680/3
C2700007|T191|OP|C80281|NCI|EBV Positive Diffuse Large B-Cell Lymphoma of the Elderly|9680/3
C2700007|T191|PT|C80281|NCI|EBV-Positive Diffuse Large B-Cell Lymphoma, Not Otherwise Specified|9680/3
C2700007|T191|SY|C80281|NCI|EBV-Positive DLBCL, NOS|9680/3
C2700007|T191|OP|C80281|NCI|Epstein-Barr Virus Positive Diffuse Large B-Cell Lymphoma of the Elderly|9680/3
C2700007|T191|SY|C80281|NCI|Epstein-Barr Virus Positive DLBCL, NOS|9680/3
C2700007|T191|SY|C80281|NCI|Epstein-Barr Virus-Positive Diffuse Large B-Cell Lymphoma, Not Otherwise Specified|9680/3
C2698294|T191|AB|C80291|NCI|HGBL, NOS|9680/3
C2698294|T191|SY|C80291|NCI|High Grade B-Cell Lymphoma, NOS|9680/3
C2698294|T191|PT|C80291|NCI|High Grade B-Cell Lymphoma, Not Otherwise Specified|9680/3
C2698294|T191|SY|C80291|NCI|High-Grade B-Cell Lymphoma, NOS|9680/3
C2698294|T191|SY|C80291|NCI|High-Grade B-Cell Lymphoma, Not Otherwise Specified|9680/3
C1709656|T191|PT|C45194|NCI|Primary Cutaneous Diffuse Large B-Cell Lymphoma, Leg Type|9680/3
C2026186|T191|PT|C71720|NCI|Primary Diffuse Large B-Cell Lymphoma of the Central Nervous System|9680/3
C2026186|T191|SY|C71720|NCI|Primary DLBCL of the CNS|9680/3
C2700007|T191|OP|C80281|NCI|Senile EBV-Associated B-Cell Lymphoproliferative Disorder|9680/3
C1321547|T191|SY|C9496|NCI|T-Cell Rich/Histiocyte-Rich Large B-Cell Lymphoma|9680/3
C1321547|T191|SY|C9496|NCI|T-Cell/Histiocyte Rich Lymphoma|9680/3
C1321547|T191|PT|C9496|NCI|T-Cell/Histiocyte-Rich Large B-Cell Lymphoma|9680/3
C1321547|T191|SY|C9496|NCI|THRLBCL|9680/3
C0079744|T191|PT|C8851|NCI_CPTAC|Diffuse Large B-Cell Lymphoma|9680/3
C0079744|T191|PT|10012820|NCI_CTEP-SDC|Diffuse large B-cell lymphoma|9680/3
C0079744|T191|DN|C8851|NCI_CTRP|Diffuse Large B-Cell Lymphoma|9680/3
C2700007|T191|DN|C80281|NCI_CTRP|EBV-Positive Diffuse Large B-Cell Lymphoma, NOS|9680/3
C1321547|T191|DN|C9496|NCI_CTRP|T-Cell/Histiocyte-Rich Large B-Cell Lymphoma|9680/3
C0079744|T191|PT|CDR0000428286|NCI_NCI-GLOSS|diffuse large B-cell lymphoma|9680/3
C0079744|T191|AB|Xa0TG|RCD|Diff malig lymphoma-histiocyt|9680/3
C0079744|T191|AB|Xa0TG|RCD|Diff malig lymphoma-large cell|9680/3
C0079744|T191|SY|Xa0TG|RCD|Diffuse malignant lymphoma - histiocytic|9680/3
C0079744|T191|PT|Xa0TG|RCD|Diffuse malignant lymphoma - large cell|9680/3
C0079744|T191|AB|Xa0TG|RCD|Mal lymphom-large cleav+non cl|9680/3
C0079744|T191|SY|Xa0TG|RCD|Malignant lymphoma - large cell cleaved and non-cleaved|9680/3
C0079744|T191|OA|BBgR.|RCDSY|Malig lymph,large cell,diff|9680/3
C0079744|T191|OP|BBgR.|RCDSY|Malignant lymphoma, large cell, diffuse NOS|9680/3
C2698294|T191|PT|722953004|SNOMEDCT_US|B-cell lymphoma unclassifiable with features intermediate between Burkitt lymphoma and diffuse large B-cell lymphoma|9680/3
C4518409|T191|PT|734142002|SNOMEDCT_US|B-cell lymphoma with features intermediate between diffuse large B-cell lymphoma and Burkitt lymphoma|9680/3
C2698294|T191|PT|12341000132100|SNOMEDCT_US|B-cell lymphoma, unclassifiable, with features intermediate between diffuse large B-cell lymphoma and Burkitt lymphoma|9680/3
C0079744|T191|SY|46732000|SNOMEDCT_US|Diffuse large B-cell lymphoma|9680/3
C1531683|T191|PT|413990004|SNOMEDCT_US|Diffuse large B-cell lymphoma - category|9680/3
C5192818|T191|PT|787565006|SNOMEDCT_US|Diffuse large B-cell lymphoma activated B-cell subtype|9680/3
C2699776|T191|PT|734076008|SNOMEDCT_US|Diffuse large B-cell lymphoma associated with chronic inflammation|9680/3
C5192843|T191|PT|787594004|SNOMEDCT_US|Diffuse large B-cell lymphoma germinal center B-cell subtype|9680/3
C5192843|T191|PTGB|787594004|SNOMEDCT_US|Diffuse large B-cell lymphoma germinal centre B-cell subtype|9680/3
C2026186|T191|PT|734066005|SNOMEDCT_US|Diffuse large B-cell lymphoma of central nervous system|9680/3
C0079744|T191|SY|109969005|SNOMEDCT_US|Diffuse malignant lymphoma - histiocytic|9680/3
C0079744|T191|SY|109969005|SNOMEDCT_US|Diffuse malignant lymphoma - large cell|9680/3
C0079744|T191|SY|109969005|SNOMEDCT_US|Diffuse non-Hodgkin lymphoma, large cell|9680/3
C0079744|T191|SY|109969005|SNOMEDCT_US|Diffuse non-Hodgkin's lymphoma, large cell|9680/3
C2700007|T191|PT|716789004|SNOMEDCT_US|Epstein-Barr virus positive diffuse large B-cell lymphoma of elderly|9680/3
C2700007|T191|PT|716788007|SNOMEDCT_US|Epstein-Barr virus positive diffuse large B-cell lymphoma of elderly|9680/3
C1321547|T191|IS|46732000|SNOMEDCT_US|Histiocyte-rich large B-cell lymphoma|9680/3
C1321547|T191|SY|450959001|SNOMEDCT_US|Histiocyte-rich large B-cell lymphoma|9680/3
C0079744|T191|SY|109969005|SNOMEDCT_US|Lymphoma, diffuse large B cell, non Hodgkins|9680/3
C0079744|T191|SY|109969005|SNOMEDCT_US|Malignant lymphoma - large cell cleaved and non-cleaved|9680/3
C0079744|T191|SY|46732000|SNOMEDCT_US|Malignant lymphoma, histiocytic|9680/3
C0079744|T191|SY|46732000|SNOMEDCT_US|Malignant lymphoma, histiocytic, diffuse|9680/3
C0079744|T191|IS|46732000|SNOMEDCT_US|Malignant lymphoma, histiocytic, NOS|9680/3
C0079744|T191|SY|46732000|SNOMEDCT_US|Malignant lymphoma, large B-cell|9680/3
C0079744|T191|PT|46732000|SNOMEDCT_US|Malignant lymphoma, large B-cell, diffuse|9680/3
C0079744|T191|SY|46732000|SNOMEDCT_US|Malignant lymphoma, large B-cell, diffuse, no ICD-O subtype|9680/3
C0079744|T191|SY|46732000|SNOMEDCT_US|Malignant lymphoma, large B-cell, diffuse, no International Classification of Diseases for Oncology subtype|9680/3
C0079744|T191|SY|46732000|SNOMEDCT_US|Malignant lymphoma, large cell|9680/3
C0079744|T191|SY|46732000|SNOMEDCT_US|Malignant lymphoma, large cell, cleaved and noncleaved|9680/3
C0079744|T191|IS|46732000|SNOMEDCT_US|Malignant lymphoma, large cell, diffuse, NOS|9680/3
C0079744|T191|IS|46732000|SNOMEDCT_US|Malignant lymphoma, large cell, NOS|9680/3
C1636152|T191|OAP|419427007|SNOMEDCT_US|Primary cutaneous large B-cell lymphoma of the leg|9680/3
C1321547|T191|PT|724645006|SNOMEDCT_US|T-cell histiocyte rich large B-cell lymphoma|9680/3
C1321547|T191|SY|724645006|SNOMEDCT_US|T-cell hystiocyte rich large B-cell lymphoma|9680/3
C1321547|T191|IS|46732000|SNOMEDCT_US|T-cell rich large B-cell lymphoma|9680/3
C1321547|T191|SY|450959001|SNOMEDCT_US|T-cell rich large B-cell lymphoma|9680/3
C1321547|T191|IS|46732000|SNOMEDCT_US|T-cell rich/histiocyte-rich large B-cell lymphoma|9680/3
C1321547|T191|SY|450959001|SNOMEDCT_US|T-cell rich/histiocyte-rich large B-cell lymphoma|9680/3
C1321547|T191|PT|450959001|SNOMEDCT_US|T-cell/histiocyte rich large B-cell lymphoma|9680/3
C0079746|T191|PT|0000015224|CHV|immunoblastic lymphoma|9684/3
C0079746|T191|SY|0000015224|CHV|immunoblastic sarcoma|9684/3
C0079746|T191|SY|0000015224|CHV|plasmablastic lymphoma|9684/3
C3472614|T191|ET|C83.3|ICD10CM|Plasmablastic diffuse large B-cell lymphoma|9684/3
C0079746|T191|PT|MTHU037617|ICPC2ICD10ENG|immunoblastic; lymphoma|9684/3
C0079746|T191|PT|MTHU037618|ICPC2ICD10ENG|immunoblastic; sarcoma|9684/3
C0079746|T191|PT|MTHU046803|ICPC2ICD10ENG|lymphoma; immunoblastic|9684/3
C0079746|T191|PT|MTHU065904|ICPC2ICD10ENG|sarcoma; immunoblastic|9684/3
C0079746|T191|LLT|10053574|MDR|Immunoblastic lymphoma|9684/3
C0079746|T191|PT|10053574|MDR|Immunoblastic lymphoma|9684/3
C0079746|T191|LLT|10062944|MDR|Immunoblastic sarcoma|9684/3
C3472614|T191|LLT|10065039|MDR|Plasmablastic lymphoma|9684/3
C3472614|T191|PT|10065039|MDR|Plasmablastic lymphoma|9684/3
C0079746|T191|PT|357679|MEDCIN|Diffuse non-Hodgkin's lymphoma, immunoblastic|9684/3
C0079746|T191|PT|92522|MEDCIN|large cell immunoblastic lymphoma|9684/3
C0079746|T191|SY|357679|MEDCIN|malignant neoplasm lymphoma diffuse non-hodgkin's, immunoblastic|9684/3
C3472614|T191|PT|391490|MEDCIN|Plasmablastic lymphoma|9684/3
C0079746|T191|PM|D016400|MSH|Diffuse Immunoblastic Lymphosarcoma|9684/3
C0079746|T191|PM|D016400|MSH|Diffuse Immunoblastic Lymphosarcomas|9684/3
C0079746|T191|PM|D016400|MSH|Immunoblastic Large Cell Lymphoma|9684/3
C0079746|T191|DEV|D016400|MSH|IMMUNOBLASTIC LARGE LYMPHOMA|9684/3
C0079746|T191|ET|D016400|MSH|Immunoblastic Large-Cell Lymphoma|9684/3
C0079746|T191|PM|D016400|MSH|Immunoblastic Large-Cell Lymphomas|9684/3
C0079746|T191|PM|D016400|MSH|Immunoblastic Lymphoma, Large-Cell|9684/3
C0079746|T191|PM|D016400|MSH|Immunoblastic Lymphomas, Large-Cell|9684/3
C0079746|T191|ET|D016400|MSH|Immunoblastic Lymphosarcoma, Diffuse|9684/3
C0079746|T191|PM|D016400|MSH|Immunoblastic Lymphosarcomas, Diffuse|9684/3
C0079746|T191|PM|D016400|MSH|Immunoblastic Sarcoma|9684/3
C0079746|T191|PM|D016400|MSH|Immunoblastic Sarcomas|9684/3
C0079746|T191|ET|D016400|MSH|Immunoblastoma|9684/3
C0079746|T191|PM|D016400|MSH|Immunoblastomas|9684/3
C0079746|T191|PM|D016400|MSH|Large Cell Immunoblastic Lymphoma|9684/3
C0079746|T191|DEV|D016400|MSH|LARGE IMMUNOBLASTIC LYMPHOMA|9684/3
C0079746|T191|ET|D016400|MSH|Large-Cell Immunoblastic Lymphoma|9684/3
C0079746|T191|PM|D016400|MSH|Large-Cell Immunoblastic Lymphomas|9684/3
C0079746|T191|PM|D016400|MSH|Large-Cell Lymphoma, Immunoblastic|9684/3
C0079746|T191|PM|D016400|MSH|Large-Cell Lymphomas, Immunoblastic|9684/3
C0079746|T191|DEV|D016400|MSH|LYMPHOMA IMMUNOBLASTIC LARGE|9684/3
C0079746|T191|DEV|D016400|MSH|LYMPHOMA LARGE IMMUNOBLASTIC|9684/3
C0079746|T191|PM|D016400|MSH|Lymphoma, Immunoblastic Large-Cell|9684/3
C0079746|T191|ET|D016400|MSH|Lymphoma, Immunoblastic, Large Cell|9684/3
C0079746|T191|ET|D016400|MSH|Lymphoma, Immunoblastic, Large-Cell|9684/3
C0079746|T191|ET|D016400|MSH|Lymphoma, Large Cell, Immunoblastic|9684/3
C0079746|T191|PM|D016400|MSH|Lymphoma, Large-Cell Immunoblastic|9684/3
C0079746|T191|MH|D016400|MSH|Lymphoma, Large-Cell, Immunoblastic|9684/3
C3472614|T191|PM|D000069293|MSH|Lymphoma, Plasmablastic|9684/3
C0079746|T191|PM|D016400|MSH|Lymphomas, Immunoblastic Large-Cell|9684/3
C0079746|T191|PM|D016400|MSH|Lymphomas, Large-Cell Immunoblastic|9684/3
C3472614|T191|PM|D000069293|MSH|Lymphomas, Plasmablastic|9684/3
C0079746|T191|PM|D016400|MSH|Lymphosarcoma, Diffuse Immunoblastic|9684/3
C0079746|T191|PM|D016400|MSH|Lymphosarcomas, Diffuse Immunoblastic|9684/3
C3472614|T191|PM|D000069293|MSH|Plasmablastic Diffuse Large B cell Lymphoma|9684/3
C3472614|T191|ET|D000069293|MSH|Plasmablastic Diffuse Large B-cell Lymphoma|9684/3
C3472614|T191|MH|D000069293|MSH|Plasmablastic Lymphoma|9684/3
C3472614|T191|PM|D000069293|MSH|Plasmablastic Lymphomas|9684/3
C3472614|T191|PM|D000069293|MSH|Plasmablasts Diffuse Large B cell Lymphoma|9684/3
C3472614|T191|ET|D000069293|MSH|Plasmablasts Diffuse Large B-cell Lymphoma|9684/3
C0079746|T191|ET|D016400|MSH|Sarcoma, Immunoblastic|9684/3
C0079746|T191|PM|D016400|MSH|Sarcomas, Immunoblastic|9684/3
C0079746|T191|PN|NOCODE|MTH|Immunoblastic Large-Cell Lymphoma|9684/3
C3472614|T191|PN|NOCODE|MTH|Plasmablastic lymphoma|9684/3
C0079746|T191|PT|C3461|NCI|Immunoblastic Lymphoma|9684/3
C3472614|T191|AB|C7224|NCI|PBL|9684/3
C3472614|T191|PT|C7224|NCI|Plasmablastic Lymphoma|9684/3
C0079746|T191|PT|C3461|NCI_CDISC|LYMPHOMA, IMMUNOBLASTIC, MALIGNANT|9684/3
C0079746|T191|DN|C3461|NCI_CTRP|Immunoblastic Lymphoma|9684/3
C0079746|T191|AB|XE2bV|RCD|Immunobl mal lymph - larg cell|9684/3
C0079746|T191|SY|XE2bV|RCD|Immunoblastic malignant lymphoma - large cell|9684/3
C0079746|T191|SY|XE2bV|RCD|Immunoblastic sarcoma|9684/3
C0079746|T191|AB|XE2bV|RCD|Mal lymphoma - immunoblastic|9684/3
C0079746|T191|PT|XE2bV|RCD|Malignant lymphoma - immunoblastic|9684/3
C0079746|T191|AB|BBg8.|RCDSY|Malig lymph, immunoblastic|9684/3
C0079746|T191|PT|BBg8.|RCDSY|Malignant lymphoma, immunoblastic type|9684/3
C0079746|T191|SY|109966003|SNOMEDCT_US|Diffuse non-Hodgkin lymphoma, immunoblastic|9684/3
C0079746|T191|SY|109966003|SNOMEDCT_US|Diffuse non-Hodgkin's lymphoma, immunoblastic|9684/3
C0079746|T191|SY|109966003|SNOMEDCT_US|Immunoblastic malignant lymphoma - large cell|9684/3
C0079746|T191|IS|78010001|SNOMEDCT_US|Immunoblastic sarcoma|9684/3
C0079746|T191|SY|109966003|SNOMEDCT_US|Lymphoma, immunoblastic, high grade|9684/3
C0079746|T191|SY|109966003|SNOMEDCT_US|Malignant lymphoma - immunoblastic|9684/3
C3472626|T191|PT|450958009|SNOMEDCT_US|Malignant lymphoma, diffuse large B-cell, immunoblastic|9684/3
C0079746|T191|OAS|78010001|SNOMEDCT_US|Malignant lymphoma, immunoblastic|9684/3
C0079746|T191|IS|78010001|SNOMEDCT_US|Malignant lymphoma, immunoblastic, NOS|9684/3
C0079746|T191|OAP|78010001|SNOMEDCT_US|Malignant lymphoma, large B-cell, diffuse, immunoblastic|9684/3
C0079746|T191|OAS|78010001|SNOMEDCT_US|Malignant lymphoma, large cell, immunoblastic|9684/3
C0079746|T191|OAS|78010001|SNOMEDCT_US|Plasmablastic lymphoma|9684/3
C3472614|T191|PT|450909005|SNOMEDCT_US|Plasmablastic lymphoma|9684/3
C3472614|T191|PT|724648008|SNOMEDCT_US|Plasmablastic lymphoma|9684/3
C0006413|T191|ET|0000004630|AOD|Burkitt's lymphoma|9687/3
C0006413|T191|PT|0007040|CCPSS|LYMPHOMA BURKITT|9687/3
C0006413|T191|SY|0000002229|CHV|burkitt lymphoma|9687/3
C0006413|T191|SY|0000002229|CHV|burkitt lymphomas|9687/3
C0006413|T191|SY|0000002229|CHV|burkitt tumor|9687/3
C0006413|T191|PT|0000002229|CHV|burkitt's lymphoma|9687/3
C0006413|T191|SY|0000002229|CHV|burkitt's non-hodgkin's lymphoma|9687/3
C0006413|T191|SY|0000002229|CHV|burkitt's tumor|9687/3
C0006413|T191|SY|0000002229|CHV|burkitts lymphoma|9687/3
C0006413|T191|SY|0000002229|CHV|burkitts tumor|9687/3
C0343640|T191|ET|2004-6947|CSP|African lymphoma|9687/3
C0006413|T191|PT|2004-6947|CSP|Burkitt's lymphoma|9687/3
C0006413|T191|SY|2004-6947|CSP|Burkitt's tumor|9687/3
C0343640|T191|SY|NOCODE|DXP|AFRICAN LYMPHOMA|9687/3
C0006413|T191|DI|U001121|DXP|LYMPHOMA, BURKITT|9687/3
C0006413|T191|PT|HP:0030080|HPO|Burkitt lymphoma|9687/3
C0006413|T191|PS|C83.7|ICD10|Burkitt's tumour|9687/3
C0006413|T191|PX|C83.7|ICD10|Burkitt's tumour non-Hodgkin's lymphoma|9687/3
C0006413|T191|PS|C83.7|ICD10AE|Burkitt's tumor|9687/3
C0006413|T191|PX|C83.7|ICD10AE|Burkitt's tumor non-Hodgkin's lymphoma|9687/3
C1629504|T047|ET|C83.7|ICD10CM|Atypical Burkitt lymphoma|9687/3
C0006413|T191|AB|C83.7|ICD10CM|Burkitt lymphoma|9687/3
C0006413|T191|HT|C83.7|ICD10CM|Burkitt lymphoma|9687/3
C0006413|T191|AB|C83.70|ICD10CM|Burkitt lymphoma, unspecified site|9687/3
C0006413|T191|PT|C83.70|ICD10CM|Burkitt lymphoma, unspecified site|9687/3
C0006413|T191|HT|200.2|ICD9CM|Burkitt's tumor or lymphoma|9687/3
C0006413|T191|PT|MTHU013216|ICPC2ICD10ENG|Burkitt; lymphoma|9687/3
C0006413|T191|PT|MTHU013221|ICPC2ICD10ENG|Burkitt; tumor|9687/3
C0006413|T191|PT|MTHU046740|ICPC2ICD10ENG|lymphoma; Burkitt|9687/3
C0006413|T191|PT|MTHU046845|ICPC2ICD10ENG|lymphoma; undifferentiated cell, Burkitt's type|9687/3
C0006413|T191|PT|MTHU077034|ICPC2ICD10ENG|tumor; Burkitt|9687/3
C0006413|T191|PT|U000718|LCH|Burkitt's lymphoma|9687/3
C0006413|T191|PT|sh85018105|LCH_NW|Burkitt's lymphoma|9687/3
C0006413|T191|LA|LA26526-6|LNC|Burkitt lymphoma, NOS|9687/3
C0006413|T191|LLT|10006595|MDR|Burkitt's lymphoma|9687/3
C0006413|T191|PT|10006595|MDR|Burkitt's lymphoma|9687/3
C0006413|T191|LLT|10006597|MDR|Burkitt's lymphoma NOS|9687/3
C0006413|T191|HT|10006596|MDR|Burkitt's lymphomas|9687/3
C0006413|T191|LLT|10006604|MDR|Burkitt's tumor|9687/3
C0006413|T191|LLT|10006605|MDR|Burkitt's tumor or lymphoma|9687/3
C0006413|T191|LLT|10006627|MDR|Burkitt's tumour|9687/3
C0006413|T191|LLT|10073809|MDR|Burkitt's tumour or lymphoma|9687/3
C0343640|T191|PT|339724|MEDCIN|African Burkitt's lymphoma|9687/3
C0006413|T191|SY|31690|MEDCIN|Burkitt lymphoma|9687/3
C0343640|T191|SY|339724|MEDCIN|burkitt lymphoma - african|9687/3
C0006413|T191|PT|31690|MEDCIN|Burkitt's lymphoma|9687/3
C0343640|T191|PEP|D002051|MSH|African Lymphoma|9687/3
C0006413|T191|MH|D002051|MSH|Burkitt Lymphoma|9687/3
C0006413|T191|ET|D002051|MSH|Burkitt Tumor|9687/3
C0006413|T191|ET|D002051|MSH|Burkitt's Lymphoma|9687/3
C0006413|T191|ET|D002051|MSH|Burkitt's Tumor|9687/3
C0006413|T191|PM|D002051|MSH|Burkitts Lymphoma|9687/3
C0006413|T191|PM|D002051|MSH|Burkitts Tumor|9687/3
C0343640|T191|PM|D002051|MSH|Lymphoma, African|9687/3
C0006413|T191|PEP|D002051|MSH|Lymphoma, Burkitt|9687/3
C0006413|T191|PM|D002051|MSH|Lymphoma, Burkitt's|9687/3
C0006413|T191|PM|D002051|MSH|Tumor, Burkitt|9687/3
C0006413|T191|PM|D002051|MSH|Tumor, Burkitt's|9687/3
C0343640|T191|PN|NOCODE|MTH|African Burkitt's lymphoma|9687/3
C0006413|T191|PN|NOCODE|MTH|Burkitt Lymphoma|9687/3
C0006413|T191|ET|200.2|MTHICD9|Malignant lymphoma, Burkitt's type|9687/3
C0343640|T191|SY|C27122|NCI|African Burkitt Lymphoma|9687/3
C0343640|T191|SY|C27122|NCI|African Burkitt's Lymphoma|9687/3
C4330613|T191|SY|C131911|NCI|B-Cell Lymphoma with 11q Aberration Resembling Burkitt Lymphoma|9687/3
C0006413|T191|PT|C2912|NCI|Burkitt Lymphoma|9687/3
C0006413|T191|SY|TCGA|NCI|Burkitt Lymphoma|9687/3
C4330613|T191|PT|C131911|NCI|Burkitt-Like Lymphoma with 11q Aberration|9687/3
C0006413|T191|SY|C2912|NCI|Burkitt's Lymphoma|9687/3
C0343640|T191|PT|C27122|NCI|Endemic Burkitt Lymphoma|9687/3
C0343640|T191|SY|C27122|NCI|Endemic Burkitt's Lymphoma|9687/3
C1334158|T191|SY|C27915|NCI|Immunodeficiency Associated Burkitt Lymphoma|9687/3
C1334158|T191|SY|C27915|NCI|Immunodeficiency Associated Burkitt's Lymphoma|9687/3
C1334158|T191|SY|C27915|NCI|Immunodeficiency Related Burkitt Lymphoma|9687/3
C1334158|T191|SY|C27915|NCI|Immunodeficiency Related Burkitt's Lymphoma|9687/3
C1334158|T191|SY|C27915|NCI|Immunodeficiency-Associated Burkitt Lymphoma|9687/3
C1334158|T191|SY|C27915|NCI|Immunodeficiency-Associated Burkitt's Lymphoma|9687/3
C1334158|T191|PT|C27915|NCI|Immunodeficiency-Related Burkitt Lymphoma|9687/3
C1334158|T191|SY|C27915|NCI|Immunodeficiency-Related Burkitt's Lymphoma|9687/3
C4330613|T191|SY|C131911|NCI|MYC-Negative B-Cell Lymphoma with 11q Aberration Resembling Burkitt Lymphoma|9687/3
C4330613|T191|SY|C131911|NCI|MYC-Negative High-Grade B-Cell Lymphoma with 11q Aberration Resembling Burkitt Lymphoma|9687/3
C0006413|T191|SY|C2912|NCI|Small Non-Cleaved Cell Lymphoma, Burkitt's Type|9687/3
C1336077|T191|PT|C27914|NCI|Sporadic Burkitt Lymphoma|9687/3
C1336077|T191|SY|C27914|NCI|Sporadic Burkitt's Lymphoma|9687/3
C0006413|T191|PT|C2912|NCI_CPTAC|Burkitt Lymphoma|9687/3
C0006413|T191|DN|C2912|NCI_CTRP|Burkitt Lymphoma|9687/3
C4330613|T191|DN|C131911|NCI_CTRP|Burkitt-Like Lymphoma with 11q Aberration|9687/3
C0006413|T191|PT|CDR0000045203|NCI_NCI-GLOSS|Burkitt's lymphoma|9687/3
C0006413|T191|LV|CDR0000039258|PDQ|Burkitt Lymphoma|9687/3
C0006413|T191|SY|CDR0000039258|PDQ|Burkitt's Lymphoma|9687/3
C0006413|T191|SY|CDR0000039258|PDQ|Burkitt's tumor|9687/3
C0006413|T191|PT|CDR0000039258|PDQ|childhood Burkitt lymphoma|9687/3
C0006413|T191|SY|CDR0000039258|PDQ|lymphoma, Burkitt's|9687/3
C0006413|T191|SY|CDR0000039258|PDQ|NHL, Burkitt's|9687/3
C0006413|T191|SY|CDR0000039258|PDQ|non-Hodgkin's lymphoma, Burkitt's|9687/3
C0006413|T191|SY|CDR0000039258|PDQ|Small Non-Cleaved Cell Lymphoma, Burkitt's Type|9687/3
C0343640|T191|PT|X70LK|RCD|African Burkitt's lymphoma|9687/3
C0006413|T191|SY|B602.|RCD|BL - Burkitt's lymphoma|9687/3
C0006413|T191|AB|B602.|RCD|Burk typ lymphom-smll noncleav|9687/3
C0006413|T191|SY|Xa0SD|RCD|Burkitt's leukaemia|9687/3
C0006413|T191|OA|B6020|RCD|Burkitt's lymph - unspec. site|9687/3
C0006413|T191|PT|B602.|RCD|Burkitt's lymphoma|9687/3
C0006413|T191|OP|B602z|RCD|Burkitt's lymphoma NOS|9687/3
C0006413|T191|OP|B6020|RCD|Burkitt's lymphoma of unspecified site|9687/3
C0006413|T191|SY|B602.|RCD|Burkitt's tumour|9687/3
C0006413|T191|AB|B602.|RCD|Burkitt's type lymphoma-undiff|9687/3
C0006413|T191|SY|B602.|RCD|Burkitt's type malignant lymphoma - small non-cleaved|9687/3
C0006413|T191|SY|B602.|RCD|Burkitt's type malignant lymphoma - undifferentiated|9687/3
C0006413|T191|SY|Xa0SD|RCDAE|Burkitt's leukemia|9687/3
C0006413|T191|SY|B602.|RCDAE|Burkitt's tumor|9687/3
C0006413|T191|OP|BBq0.|RCDSA|Burkitt's tumor|9687/3
C0006413|T191|OP|BBqz.|RCDSA|Burkitt's tumor NOS|9687/3
C0006413|T191|OP|BBq..|RCDSA|Burkitt's tumors|9687/3
C0006413|T191|OP|BBq0.|RCDSY|Burkitt's tumour|9687/3
C0006413|T191|OP|BBqz.|RCDSY|Burkitt's tumour NOS|9687/3
C0006413|T191|OP|BBq..|RCDSY|Burkitt's tumours|9687/3
C0343640|T191|SY|240531002|SNOMEDCT_US|African Burkitt lymphoma|9687/3
C0343640|T191|PT|240531002|SNOMEDCT_US|African Burkitt's lymphoma|9687/3
C1629504|T047|SY|419879004|SNOMEDCT_US|Atypical Burkitt lymphoma|9687/3
C1629504|T047|PT|419879004|SNOMEDCT_US|Atypical Burkitt's lymphoma|9687/3
C0006413|T191|SY|118617000|SNOMEDCT_US|BL - Burkitt's lymphoma|9687/3
C0006413|T191|SY|118617000|SNOMEDCT_US|Burkitt lymphoma|9687/3
C0006413|T191|PT|77381001|SNOMEDCT_US|Burkitt lymphoma|9687/3
C0006413|T191|PTGB|397400006|SNOMEDCT_US|Burkitt lymphoma/leukaemia|9687/3
C0006413|T191|PT|397400006|SNOMEDCT_US|Burkitt lymphoma/leukemia|9687/3
C4330613|T191|PT|783220004|SNOMEDCT_US|Burkitt-like lymphoma with 11q aberration|9687/3
C0006413|T191|SY|118617000|SNOMEDCT_US|Burkitt's lymphoma|9687/3
C0006413|T191|SY|77381001|SNOMEDCT_US|Burkitt's lymphoma|9687/3
C0006413|T191|OAP|154581008|SNOMEDCT_US|Burkitt's lymphoma|9687/3
C0006413|T191|OF|154581008|SNOMEDCT_US|Burkitt's lymphoma|9687/3
C0006413|T191|SY|118617000|SNOMEDCT_US|Burkitt's lymphoma - disorder|9687/3
C0006413|T191|OAP|188518008|SNOMEDCT_US|Burkitt's lymphoma NOS|9687/3
C0006413|T191|OAP|188509006|SNOMEDCT_US|Burkitt's lymphoma of unspecified site|9687/3
C0006413|T191|IS|77381001|SNOMEDCT_US|Burkitt's lymphoma, NOS|9687/3
C0006413|T191|SY|118617000|SNOMEDCT_US|Burkitt's tumor|9687/3
C0006413|T191|IS|77381001|SNOMEDCT_US|Burkitt's tumor|9687/3
C0006413|T191|SYGB|118617000|SNOMEDCT_US|Burkitt's tumour|9687/3
C0006413|T191|SY|118617000|SNOMEDCT_US|Burkitt's type malignant lymphoma - small non-cleaved|9687/3
C0006413|T191|SY|118617000|SNOMEDCT_US|Burkitt's type malignant lymphoma - undifferentiated|9687/3
C0343640|T191|SY|419770008|SNOMEDCT_US|Endemic Burkitt lymphoma|9687/3
C0343640|T191|PT|419770008|SNOMEDCT_US|Endemic Burkitt's lymphoma|9687/3
C1334158|T191|SY|419094004|SNOMEDCT_US|Immunodeficiency-associated Burkitt lymphoma|9687/3
C1334158|T191|PT|419094004|SNOMEDCT_US|Immunodeficiency-associated Burkitt's lymphoma|9687/3
C0006413|T191|SY|77381001|SNOMEDCT_US|Malignant lymphoma, small noncleaved, Burkitt's, diffuse|9687/3
C0006413|T191|IS|77381001|SNOMEDCT_US|Malignant lymphoma, undifferentiated, Burkitt's type|9687/3
C1336077|T191|SY|420063007|SNOMEDCT_US|Non-endemic Burkitt's lymphoma|9687/3
C1336077|T191|SY|420063007|SNOMEDCT_US|Sporadic Burkitt lymphoma|9687/3
C1336077|T191|PT|420063007|SNOMEDCT_US|Sporadic Burkitt's lymphoma|9687/3
C1321547|T191|LLT|10080211|MDR|T-cell/histiocyte-rich large B-cell lymphoma|9688/3
C1321547|T191|SY|C9496|NCI|T-Cell Rich/Histiocyte-Rich Large B-Cell Lymphoma|9688/3
C1321547|T191|SY|C9496|NCI|T-Cell/Histiocyte Rich Lymphoma|9688/3
C1321547|T191|PT|C9496|NCI|T-Cell/Histiocyte-Rich Large B-Cell Lymphoma|9688/3
C1321547|T191|SY|C9496|NCI|THRLBCL|9688/3
C1321547|T191|DN|C9496|NCI_CTRP|T-Cell/Histiocyte-Rich Large B-Cell Lymphoma|9688/3
C1321547|T191|IS|46732000|SNOMEDCT_US|Histiocyte-rich large B-cell lymphoma|9688/3
C1321547|T191|SY|450959001|SNOMEDCT_US|Histiocyte-rich large B-cell lymphoma|9688/3
C1321547|T191|PT|724645006|SNOMEDCT_US|T-cell histiocyte rich large B-cell lymphoma|9688/3
C1321547|T191|SY|724645006|SNOMEDCT_US|T-cell hystiocyte rich large B-cell lymphoma|9688/3
C1321547|T191|IS|46732000|SNOMEDCT_US|T-cell rich large B-cell lymphoma|9688/3
C1321547|T191|SY|450959001|SNOMEDCT_US|T-cell rich large B-cell lymphoma|9688/3
C1321547|T191|IS|46732000|SNOMEDCT_US|T-cell rich/histiocyte-rich large B-cell lymphoma|9688/3
C1321547|T191|SY|450959001|SNOMEDCT_US|T-cell rich/histiocyte-rich large B-cell lymphoma|9688/3
C1321547|T191|PT|450959001|SNOMEDCT_US|T-cell/histiocyte rich large B-cell lymphoma|9688/3
C0349632|T191|SY|0000031272|CHV|lymphoma splenic marginal zone|9689/3
C0349632|T191|SY|0000031272|CHV|marginal zone splenic lymphoma|9689/3
C0349632|T191|PT|0000031272|CHV|splenic marginal zone lymphoma|9689/3
C0349632|T191|ET|C83.0|ICD10CM|Splenic marginal zone lymphoma|9689/3
C0349632|T191|AB|200.37|ICD9CM|Margin zone lymph spleen|9689/3
C0349632|T191|PT|200.37|ICD9CM|Marginal zone lymphoma, spleen|9689/3
C0349632|T191|LLT|10062113|MDR|Splenic marginal zone lymphoma|9689/3
C0349632|T191|PT|10062113|MDR|Splenic marginal zone lymphoma|9689/3
C0349632|T191|LLT|10041651|MDR|Splenic marginal zone lymphoma NOS|9689/3
C0349632|T191|HT|10041650|MDR|Splenic marginal zone lymphomas|9689/3
C0349632|T191|SY|354827|MEDCIN|leukemia lymphocytic chronic splenic with villous lymphocytes|9689/3
C0349632|T191|PT|230964|MEDCIN|marginal zone B-cell lymphoma of spleen|9689/3
C0349632|T191|PT|230975|MEDCIN|marginal zone lymphoma of spleen|9689/3
C0349632|T191|PT|354827|MEDCIN|Splenic lymphoma with villous lymphocytes|9689/3
C0349632|T191|PN|NOCODE|MTH|Splenic Marginal Zone B-Cell Lymphoma|9689/3
C0349632|T191|ET|200.37|MTHICD9|Marginal zone lymphoma involving spleen|9689/3
C0349632|T191|ET|200.3|MTHICD9|Splenic marginal zone B-cell lymphoma|9689/3
C0349632|T191|SY|C4663|NCI|Marginal Zone Lymphoma of Spleen|9689/3
C0349632|T191|SY|C4663|NCI|Marginal Zone Lymphoma of the Spleen|9689/3
C0349632|T191|AB|C4663|NCI|SLVL|9689/3
C0349632|T191|AB|C4663|NCI|SMZL|9689/3
C0349632|T191|SY|C4663|NCI|Splenic Lymphoma with Circulating Villous Lymphocytes|9689/3
C0349632|T191|SY|C4663|NCI|Splenic Marginal Zone B-Cell Lymphoma|9689/3
C0349632|T191|SY|C4663|NCI|Splenic Marginal Zone B-Cell Lymphoma with Villous Lymphocytes|9689/3
C0349632|T191|SY|TCGA|NCI|Splenic Marginal Zone Lymphoma|9689/3
C0349632|T191|PT|C4663|NCI|Splenic Marginal Zone Lymphoma|9689/3
C0349632|T191|SY|C4663|NCI|Splenic Marginal Zone Lymphoma with Villous Lymphocytes|9689/3
C0349632|T191|DN|C4663|NCI_CTRP|Splenic Marginal Zone Lymphoma|9689/3
C0349632|T191|SY|CDR0000372809|PDQ|marginal zone lymphoma of spleen|9689/3
C0349632|T191|SY|CDR0000372809|PDQ|marginal zone lymphoma of the spleen|9689/3
C0349632|T191|AB|CDR0000372809|PDQ|SMZL|9689/3
C0349632|T191|SY|CDR0000372809|PDQ|splenic marginal zone B-cell lymphoma|9689/3
C0349632|T191|PT|CDR0000372809|PDQ|splenic marginal zone lymphoma|9689/3
C0349632|T191|AB|Xa0Rp|RCD|Splen lymphom with vill lympho|9689/3
C0349632|T191|PT|Xa0Rp|RCD|Splenic lymphoma with villous lymphocytes|9689/3
C0349632|T191|PT|116691000119101|SNOMEDCT_US|Marginal zone lymphoma of spleen|9689/3
C0349632|T191|PT|277551008|SNOMEDCT_US|Splenic lymphoma with villous lymphocytes|9689/3
C0349632|T191|SY|128802003|SNOMEDCT_US|Splenic lymphoma with villous lymphocytes|9689/3
C0349632|T191|PT|763666008|SNOMEDCT_US|Splenic marginal zone B-cell lymphoma|9689/3
C0349632|T191|PT|128802003|SNOMEDCT_US|Splenic marginal zone B-cell lymphoma|9689/3
C0349632|T191|SY|128802003|SNOMEDCT_US|Splenic marginal zone lymphoma|9689/3
C0024301|T191|PT|0000007618|CHV|follicular lymphoma|9690/3
C0024301|T191|SY|0000007618|CHV|follicular lymphomas|9690/3
C0024301|T191|SY|0000007618|CHV|giant follicular lymphoma|9690/3
C0024301|T191|SY|0000007618|CHV|lymphoma follicular|9690/3
C0024301|T191|SY|0000007618|CHV|lymphosarcoma follicular|9690/3
C0024301|T191|SY|0000007618|CHV|nodular lymphoma|9690/3
C0024301|T191|ET|4001-0094|CSP|follicular lymphoma|9690/3
C0024301|T191|PT|C82.9|ICD10|Follicular non-Hodgkin's lymphoma, unspecified|9690/3
C0024301|T191|HT|C82|ICD10CM|Follicular lymphoma|9690/3
C0024301|T191|AB|C82|ICD10CM|Follicular lymphoma|9690/3
C0024301|T191|AB|C82.9|ICD10CM|Follicular lymphoma, unspecified|9690/3
C0024301|T191|HT|C82.9|ICD10CM|Follicular lymphoma, unspecified|9690/3
C0024301|T191|HT|202.0|ICD9CM|Nodular lymphoma|9690/3
C0024301|T191|PT|MTHU012702|ICPC2ICD10ENG|Brill-Symmers|9690/3
C0024301|T191|PT|MTHU029202|ICPC2ICD10ENG|follicular; germinoblastoma|9690/3
C0024301|T191|PT|MTHU029212|ICPC2ICD10ENG|follicular; lymphosarcoma|9690/3
C0024301|T191|PT|MTHU031394|ICPC2ICD10ENG|germinoblastoma; follicular|9690/3
C0024301|T191|PT|MTHU046695|ICPC2ICD10ENG|lymphocytic; lymphoma, nodular|9690/3
C0024301|T191|PT|MTHU046770|ICPC2ICD10ENG|lymphoma; follicular|9690/3
C0024301|T191|PT|MTHU046818|ICPC2ICD10ENG|lymphoma; lymphocytic, nodular|9690/3
C0024301|T191|PT|MTHU046833|ICPC2ICD10ENG|lymphoma; nodular|9690/3
C0024301|T191|PT|MTHU046837|ICPC2ICD10ENG|lymphoma; nodular, lymphocytic|9690/3
C0024301|T191|PT|MTHU046878|ICPC2ICD10ENG|lymphosarcoma; follicular|9690/3
C0024301|T191|PT|MTHU053410|ICPC2ICD10ENG|nodular; lymphoma|9690/3
C0024301|T191|PT|MTHU053414|ICPC2ICD10ENG|nodular; lymphoma, lymphocytic|9690/3
C0024301|T191|LLT|10029478|MDR|Nodular lymphoma|9690/3
C2698750|T191|LLT|10080376|MDR|Paediatric-type follicular lymphoma|9690/3
C2698750|T191|LLT|10080207|MDR|Pediatric-type follicular lymphoma|9690/3
C0024301|T191|PT|355312|MEDCIN|Follicular low grade B-cell lymphoma|9690/3
C0024301|T191|PT|335952|MEDCIN|follicular lymphoma|9690/3
C0024301|T191|PT|357184|MEDCIN|follicular malignant lymphoma - centroblastic-centrocytic|9690/3
C0024301|T191|PT|273324|MEDCIN|giant follicular lymphosarcoma|9690/3
C0024301|T191|SY|355312|MEDCIN|malignant neoplasm lymphoma b-cell low grade follicular|9690/3
C0024301|T191|SY|357184|MEDCIN|malignant neoplasm lymphoma follicular - centroblastic-centrocytic|9690/3
C0024301|T191|SY|335952|MEDCIN|malignant neoplasm nodular lymphoma follicular|9690/3
C0024301|T191|SY|31696|MEDCIN|nodular lymphoma|9690/3
C0024301|T191|PT|273325|MEDCIN|nodular lymphosarcoma|9690/3
C0024301|T191|PT|31696|MEDCIN|nodular malignant lymphoma|9690/3
C0024301|T191|DEV|D008224|MSH|BRILL SYMMERS DIS|9690/3
C0024301|T191|PM|D008224|MSH|Brill Symmers Disease|9690/3
C0024301|T191|ET|D008224|MSH|Brill-Symmers Disease|9690/3
C0024301|T191|PM|D008224|MSH|Disease, Brill-Symmers|9690/3
C0024301|T191|DEV|D008224|MSH|FOLLIC LYMPHOMA|9690/3
C0024301|T191|DEV|D008224|MSH|FOLLIC LYMPHOMA GIANT|9690/3
C0024301|T191|ET|D008224|MSH|Follicular Lymphoma|9690/3
C0024301|T191|ET|D008224|MSH|Follicular Lymphoma, Giant|9690/3
C0024301|T191|PM|D008224|MSH|Follicular Lymphomas|9690/3
C0024301|T191|PM|D008224|MSH|Follicular Lymphomas, Giant|9690/3
C0024301|T191|DEV|D008224|MSH|GIANT FOLLIC LYMPHOMA|9690/3
C0024301|T191|ET|D008224|MSH|Giant Follicular Lymphoma|9690/3
C0024301|T191|PM|D008224|MSH|Giant Follicular Lymphomas|9690/3
C0024301|T191|DEV|D008224|MSH|LYMPHOMA FOLLIC|9690/3
C0024301|T191|DEV|D008224|MSH|LYMPHOMA GIANT FOLLIC|9690/3
C0024301|T191|MH|D008224|MSH|Lymphoma, Follicular|9690/3
C0024301|T191|ET|D008224|MSH|Lymphoma, Giant Follicular|9690/3
C0024301|T191|ET|D008224|MSH|Lymphoma, Nodular|9690/3
C0024301|T191|PM|D008224|MSH|Lymphomas, Follicular|9690/3
C0024301|T191|PM|D008224|MSH|Lymphomas, Giant Follicular|9690/3
C0024301|T191|PM|D008224|MSH|Lymphomas, Nodular|9690/3
C0024301|T191|PM|D008224|MSH|Nodular Lymphoma|9690/3
C0024301|T191|PM|D008224|MSH|Nodular Lymphomas|9690/3
C0024301|T191|PN|NOCODE|MTH|Lymphoma, Follicular|9690/3
C0024301|T191|ET|202.0|MTHICD9|Brill-Symmers disease|9690/3
C0024301|T191|ET|202.0|MTHICD9|Follicular lymphoma|9690/3
C0024301|T191|ET|202.0|MTHICD9|Follicular lymphosarcoma|9690/3
C0024301|T191|ET|202.0|MTHICD9|Giant follicular lymphoma|9690/3
C0024301|T191|ET|202.0|MTHICD9|Giant follicular lymphosarcoma|9690/3
C0024301|T191|ET|202.0|MTHICD9|Nodular lymphocytic lymphoma|9690/3
C0024301|T191|ET|202.0|MTHICD9|Nodular lymphosarcoma|9690/3
C2698750|T191|OP|C80297|NCI|Childhood Follicular Lymphoma|9690/3
C0024301|T191|SY|C3209|NCI|Follicle Center Lymphoma|9690/3
C0024301|T191|PT|C3209|NCI|Follicular Lymphoma|9690/3
C0024301|T191|SY|TCGA|NCI|Follicular Lymphoma|9690/3
C0024301|T191|SY|C3209|NCI|Follicular Non-Hodgkin Lymphoma|9690/3
C0024301|T191|SY|C3209|NCI|Follicular Non-Hodgkin's Lymphoma|9690/3
C2698750|T191|OP|C80297|NCI|Pediatric Follicular Lymphoma|9690/3
C2698750|T191|PT|C80297|NCI|Pediatric-Type Follicular Lymphoma|9690/3
C0024301|T191|SY|C3209|NCI_CDISC|Follicle Center Lymphoma|9690/3
C0024301|T191|SY|C3209|NCI_CDISC|Follicular Centre Cell Lymphoma|9690/3
C0024301|T191|SY|C3209|NCI_CDISC|Follicular Non-Hodgkin Lymphoma|9690/3
C0024301|T191|SY|C3209|NCI_CDISC|Follicular Non-Hodgkin's Lymphoma|9690/3
C0024301|T191|SY|C3209|NCI_CDISC|Lymphoma, Follicular Centre Cell|9690/3
C0024301|T191|PT|C3209|NCI_CDISC|LYMPHOMA, FOLLICULAR, MALIGNANT|9690/3
C0024301|T191|PT|C3209|NCI_CPTAC|Follicular Lymphoma|9690/3
C0024301|T191|PT|10016896|NCI_CTEP-SDC|Follicular lymphoma|9690/3
C0024301|T191|DN|C3209|NCI_CTRP|Follicular Lymphoma|9690/3
C0024301|T191|PT|CDR0000428287|NCI_NCI-GLOSS|follicular lymphoma|9690/3
C2698750|T191|PT|C80297|NCI_NICHD|Childhood Follicular Lymphoma|9690/3
C2698750|T191|SY|C80297|NCI_NICHD|Pediatric Follicular Lymphoma|9690/3
C0024301|T191|SY|CDR0000795359|PDQ|follicle center lymphoma|9690/3
C0024301|T191|PT|CDR0000795359|PDQ|follicular lymphoma|9690/3
C0024301|T191|SY|CDR0000795359|PDQ|follicular non-Hodgkin lymphoma|9690/3
C0024301|T191|SY|CDR0000795359|PDQ|follicular non-Hodgkin's lymphoma|9690/3
C0024301|T191|IS|Xa9FF|RCD|Brill - Symmers' disease|9690/3
C0024301|T191|AB|Xa0T4|RCD|Foll low grade B-cell lymphom|9690/3
C0024301|T191|PT|Xa0T4|RCD|Follicular low grade B-cell lymphoma|9690/3
C0024301|T191|IS|Xa9FF|RCD|Follicular lymphosarcoma|9690/3
C0024301|T191|AB|XaBLw|RCD|Follicular non-Hodgkin's lymph|9690/3
C0024301|T191|PT|XaBLw|RCD|Follicular non-Hodgkin's lymphoma|9690/3
C0024301|T191|SY|XaBBf|RCD|Germinoblastoma, follicular|9690/3
C0024301|T191|IS|Xa9FF|RCD|Giant follicular lymphoma|9690/3
C0024301|T191|AB|XaBBf|RCD|M lyoma,centrbl-centrcyt,foll|9690/3
C0024301|T191|PT|XaBBf|RCD|Malignant lymphoma, centroblastic-centrocytic, follicular|9690/3
C0024301|T191|OP|Xa9FF|RCD|Malignant lymphoma, nodular|9690/3
C0024301|T191|OP|XE1vp|RCD|Nodular lymphoma|9690/3
C0024301|T191|OP|B620z|RCD|Nodular lymphoma NOS|9690/3
C0024301|T191|OP|B6200|RCD|Nodular lymphoma of unspecified site|9690/3
C0024301|T191|OA|B6200|RCD|Nodular lymphoma-unspec. site|9690/3
C0024301|T191|IS|Xa9FF|RCD|Nodular lymphosarcoma|9690/3
C0024301|T191|SY|Xa0T4|RCD|Nodular malignant lymphoma|9690/3
C0024301|T191|AB|BBk2.|RCDSY|Mal.lym,centr-blas/cyt,foll|9690/3
C0024301|T191|OA|XE1wf|RCDSY|Malig.lymphoma, nodular NOS|9690/3
C0024301|T191|PT|BBk2.|RCDSY|Malignant lymphoma, centroblastic-centrocytic, follicular|9690/3
C0024301|T191|OP|XE1wf|RCDSY|Malignant lymphoma, nodular NOS|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Brill - Symmers' disease|9690/3
C0024301|T191|PT|277618009|SNOMEDCT_US|Follicular low grade B-cell lymphoma|9690/3
C0024301|T191|PT|55150002|SNOMEDCT_US|Follicular lymphoma|9690/3
C0024301|T191|OAS|188681004|SNOMEDCT_US|Follicular lymphoma NOS|9690/3
C1301454|T191|PT|397467006|SNOMEDCT_US|Follicular lymphoma, cutaneous follicle center sub-type|9690/3
C1301454|T191|PTGB|397467006|SNOMEDCT_US|Follicular lymphoma, cutaneous follicle centre sub-type|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Follicular lymphosarcoma|9690/3
C0024301|T191|SY|308121000|SNOMEDCT_US|Follicular non-Hodgkin lymphoma|9690/3
C0024301|T191|OAS|188681004|SNOMEDCT_US|Follicular non-Hodgkin's lymphoma|9690/3
C0024301|T191|PT|308121000|SNOMEDCT_US|Follicular non-Hodgkin's lymphoma|9690/3
C0024301|T191|SY|307637005|SNOMEDCT_US|Germinoblastoma, follicular|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Giant follicular lymphoma|9690/3
C0024301|T191|OAP|46324005|SNOMEDCT_US|Malignant lymphoma, centroblastic-centrocytic, follicular|9690/3
C0024301|T191|PT|307637005|SNOMEDCT_US|Malignant lymphoma, centroblastic-centrocytic, follicular|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Malignant lymphoma, centroblastic-centrocytic, follicular|9690/3
C0024301|T191|IS|46324005|SNOMEDCT_US|Malignant lymphoma, centroblastic-centrocytic, follicular -RETIRED-|9690/3
C0024301|T191|OF|46324005|SNOMEDCT_US|Malignant lymphoma, centroblastic-centrocytic, follicular -RETIRED-|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Malignant lymphoma, follicle center|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Malignant lymphoma, follicle center, follicular|9690/3
C0024301|T191|SYGB|55150002|SNOMEDCT_US|Malignant lymphoma, follicle centre|9690/3
C0024301|T191|SYGB|55150002|SNOMEDCT_US|Malignant lymphoma, follicle centre, follicular|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Malignant lymphoma, follicular|9690/3
C0024301|T191|IS|55150002|SNOMEDCT_US|Malignant lymphoma, follicular, NOS|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Malignant lymphoma, lymphocytic, nodular|9690/3
C0024301|T191|IS|55150002|SNOMEDCT_US|Malignant lymphoma, lymphocytic, nodular, NOS|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Malignant lymphoma, nodular|9690/3
C0024301|T191|IS|55150002|SNOMEDCT_US|Malignant lymphoma, nodular, NOS|9690/3
C0024301|T191|PT|269476000|SNOMEDCT_US|Nodular lymphoma|9690/3
C0024301|T191|OAP|188617008|SNOMEDCT_US|Nodular lymphoma NOS|9690/3
C0024301|T191|OAP|188608008|SNOMEDCT_US|Nodular lymphoma of unspecified site|9690/3
C0024301|T191|SY|55150002|SNOMEDCT_US|Nodular lymphosarcoma|9690/3
C0024301|T191|SY|277618009|SNOMEDCT_US|Nodular malignant lymphoma|9690/3
C2698750|T191|PTGB|736322001|SNOMEDCT_US|Paediatric follicular lymphoma|9690/3
C2698750|T191|PTGB|733917002|SNOMEDCT_US|Paediatric follicular lymphoma|9690/3
C2698750|T191|PT|736322001|SNOMEDCT_US|Pediatric follicular lymphoma|9690/3
C2698750|T191|PT|733917002|SNOMEDCT_US|Pediatric follicular lymphoma|9690/3
C0024301|T191|OAS|188607003|SNOMEDCT_US|Reticulosarcoma - follicular or nodular|9690/3
C0079758|T191|PT|0000015227|CHV|follicular mixed cell lymphoma|9691/3
C0079758|T191|PS|C82.1|ICD10|Mixed small cleaved and large cell, follicular|9691/3
C0079758|T191|PX|C82.1|ICD10|Mixed small cleaved and large cell, follicular non-Hodgkin's lymphoma|9691/3
C0079758|T191|AB|C82.1|ICD10CM|Follicular lymphoma grade II|9691/3
C0079758|T191|HT|C82.1|ICD10CM|Follicular lymphoma grade II|9691/3
C0079758|T191|PT|MTHU029206|ICPC2ICD10ENG|follicular; lymphoma, mixed cell type|9691/3
C0079758|T191|PT|MTHU029210|ICPC2ICD10ENG|follicular; lymphoma, small cell, cleaved, and large cell|9691/3
C0079758|T191|PT|MTHU029213|ICPC2ICD10ENG|follicular; lymphosarcoma, mixed cell type|9691/3
C0079758|T191|PT|MTHU029214|ICPC2ICD10ENG|follicular; reticulolymphosarcoma|9691/3
C0079758|T191|PT|MTHU046773|ICPC2ICD10ENG|lymphoma; follicular, mixed cell type|9691/3
C0079758|T191|PT|MTHU046779|ICPC2ICD10ENG|lymphoma; follicular, small cell, cleaved, and large cell|9691/3
C0079758|T191|PT|MTHU046790|ICPC2ICD10ENG|lymphoma; mixed cell type, follicular|9691/3
C0079758|T191|PT|MTHU046835|ICPC2ICD10ENG|lymphoma; nodular, mixed lymphocytic-histiocytic|9691/3
C0079758|T191|PT|MTHU046879|ICPC2ICD10ENG|lymphosarcoma; follicular, mixed cell type|9691/3
C0079758|T191|PT|MTHU053412|ICPC2ICD10ENG|nodular; lymphoma, mixed lymphocytic-histiocytic|9691/3
C0079758|T191|PT|MTHU053419|ICPC2ICD10ENG|nodular; reticulolymphosarcoma|9691/3
C0079758|T191|PT|MTHU064358|ICPC2ICD10ENG|reticulolymphosarcoma; follicular|9691/3
C0079758|T191|PT|MTHU064359|ICPC2ICD10ENG|reticulolymphosarcoma; nodular|9691/3
C0079758|T191|PT|357183|MEDCIN|Follicular malignant lymphoma - mixed cell type|9691/3
C0079758|T191|PT|357970|MEDCIN|follicular non-Hodgkin's lymphoma, mixed small cleaved and large cell|9691/3
C0079758|T191|PT|357968|MEDCIN|Follicular non-Hodgkin's lymphoma, mixed small cleaved cell and large cell|9691/3
C0079758|T191|SY|357968|MEDCIN|malig lymphoma follicular, non-hodgkin's mixed small cleaved cell and large cell|9691/3
C0079758|T191|SY|357970|MEDCIN|malignant lymphoma follicular, non-hodgkin's mixed small cleaved and large cell|9691/3
C0079758|T191|SY|357183|MEDCIN|malignant neoplasm lymphoma b-cell low grade follicular mixed cell type|9691/3
C0079758|T191|DEV|D008224|MSH|FOLLIC MIXED LYMPHOMA|9691/3
C0079758|T191|PM|D008224|MSH|Follicular Mixed Cell Lymphoma|9691/3
C0079758|T191|ET|D008224|MSH|Follicular Mixed-Cell Lymphoma|9691/3
C0079758|T191|PM|D008224|MSH|Follicular Mixed-Cell Lymphomas|9691/3
C0079758|T191|DEV|D008224|MSH|LYMPHOMA FOLLIC MIXED|9691/3
C0079758|T191|DEV|D008224|MSH|LYMPHOMA FOLLIC MIXED LYMPHOCYTIC HISTIOCYTIC|9691/3
C0079758|T191|DEV|D008224|MSH|LYMPHOMA FOLLIC MIXED SMALL LARGE LYMPHOID|9691/3
C0079758|T191|DEV|D008224|MSH|LYMPHOMA FOLLIC SMALL LARGE CLEAVED|9691/3
C0079758|T191|DEV|D008224|MSH|LYMPHOMA MIXED FOLLIC|9691/3
C0079758|T191|DEV|D008224|MSH|LYMPHOMA NODULAR MIXED SMALL LARGE|9691/3
C0079758|T191|PM|D008224|MSH|Lymphoma, Follicular Mixed-Cell|9691/3
C0079758|T191|ET|D008224|MSH|Lymphoma, Follicular, Mixed Cell|9691/3
C0079758|T191|ET|D008224|MSH|Lymphoma, Follicular, Mixed Lymphocytic-Histiocytic|9691/3
C0079758|T191|ET|D008224|MSH|Lymphoma, Follicular, Mixed Small and Large Lymphoid|9691/3
C0079758|T191|ET|D008224|MSH|Lymphoma, Follicular, Small and Large Cleaved Cell|9691/3
C0079758|T191|ET|D008224|MSH|Lymphoma, Follicular, Small and Large Cleaved-Cell|9691/3
C0079758|T191|PEP|D008224|MSH|Lymphoma, Mixed-Cell, Follicular|9691/3
C0079758|T191|ET|D008224|MSH|Lymphoma, Nodular, Mixed Lymphocytic Histiocytic|9691/3
C0079758|T191|ET|D008224|MSH|Lymphoma, Nodular, Mixed Lymphocytic-Histiocytic|9691/3
C0079758|T191|ET|D008224|MSH|Lymphoma, Nodular, Mixed Small and Large Cell|9691/3
C0079758|T191|PM|D008224|MSH|Lymphomas, Follicular Mixed-Cell|9691/3
C0079758|T191|PM|D008224|MSH|Mixed Cell Lymphoma, Follicular|9691/3
C0079758|T191|DEV|D008224|MSH|MIXED LYMPHOMA FOLLIC|9691/3
C0079758|T191|ET|D008224|MSH|Mixed-Cell Lymphoma, Follicular|9691/3
C0079758|T191|PM|D008224|MSH|Mixed-Cell Lymphomas, Follicular|9691/3
C0079758|T191|PN|NOCODE|MTH|Lymphoma, Mixed-Cell, Follicular|9691/3
C0079758|T191|SY|C8968|NCI|Follicular Mixed Cell Lymphoma|9691/3
C0079758|T191|SY|C8968|NCI|Follicular Mixed Lymphocytic-Histiocytic Lymphoma|9691/3
C0079758|T191|PT|C8968|NCI|Grade 2 Follicular Lymphoma|9691/3
C0079758|T191|SY|TCGA|NCI|Grade 2 Follicular Lymphoma|9691/3
C0079758|T191|SY|C8968|NCI|Grade II Follicular Lymphoma|9691/3
C0079758|T191|SY|C8968|NCI|Grade II Follicular Mixed Cell Lymphoma|9691/3
C0079758|T191|SY|C8968|NCI|Nodular Mixed Lymphoma|9691/3
C0079758|T191|PT|C8968|NCI_CPTAC|Grade 2 Follicular Lymphoma|9691/3
C0079758|T191|DN|C8968|NCI_CTRP|Grade 2 Follicular Lymphoma|9691/3
C0079758|T191|PT|CDR0000349454|NCI_NCI-GLOSS|follicular mixed cell lymphoma|9691/3
C0079758|T191|PT|CDR0000430862|NCI_NCI-GLOSS|grade 2 follicular lymphoma|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|FM lymphoma|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|follicular mixed cell lymphoma|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|Follicular Mixed Lymphocytic-Histiocytic Lymphoma|9691/3
C0079758|T191|PT|CDR0000038359|PDQ|grade 2 follicular lymphoma|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|Grade II Follicular Lymphoma|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|grade II follicular mixed cell lymphoma|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|lymphoma, follicular mixed cell|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|lymphoma, nodular mixed|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|mixed cell lymphoma, follicular|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|NM lymphoma|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|NML|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|nodular MC lymphoma|9691/3
C0079758|T191|SY|CDR0000038359|PDQ|nodular mixed lymphoma|9691/3
C0079758|T191|AB|Xa0TA|RCD|Fol mal lymph-mix small+large|9691/3
C0079758|T191|OA|B6271|RCD|Fol non-H mix sm cl/lg cel lym|9691/3
C0079758|T191|AB|Xa0TA|RCD|Foll malig lymphom - mix cell|9691/3
C0079758|T191|AB|Xa0TA|RCD|Follicular malig lymphoma - mix small cleaved and large cell|9691/3
C0079758|T191|PT|Xa0TA|RCD|Follicular malignant lymphoma - mixed cell type|9691/3
C0079758|T191|SY|Xa0TA|RCD|Follicular malignant lymphoma - mixed small cleaved and large cell|9691/3
C0079758|T191|OA|B6271|RCD|Follicular non-Hodg mixed sml cleavd & lge cell lymphoma|9691/3
C0079758|T191|OP|B6271|RCD|Follicular non-Hodgkin's mixed small cleaved and large cell lymphoma|9691/3
C0079758|T191|AB|XaBBd|RCD|M lyoma,lymphcyt-histcyt,nod|9691/3
C0079758|T191|PT|XaBBd|RCD|Malignant lymphoma, mixed lymphocytic-histiocytic, nodular|9691/3
C0079758|T191|AB|XaBBd|RCD|Reticulolymphosarc,follicular|9691/3
C0079758|T191|SY|XaBBd|RCD|Reticulolymphosarcoma, follicular|9691/3
C0079758|T191|SY|XaBBd|RCD|Reticulolymphosarcoma, nodular|9691/3
C0079758|T191|AB|BBk1.|RCDSY|Malig lymphoma, mixed lymphocytic-histiocytic, nodular|9691/3
C0079758|T191|AB|BBk1.|RCDSY|Malig.lymph,lymph/hist,nod.|9691/3
C0079758|T191|PT|BBk1.|RCDSY|Malignant lymphoma, mixed lymphocytic-histiocytic, nodular|9691/3
C0079758|T191|SY|109971005|SNOMEDCT_US|Follicular lymphoma grade 2|9691/3
C1301456|T191|PT|397469009|SNOMEDCT_US|Follicular lymphoma, diffuse follicle center cell sub-type, grade 2|9691/3
C1301456|T191|PTGB|397469009|SNOMEDCT_US|Follicular lymphoma, diffuse follicle centre cell sub-type, grade 2|9691/3
C0079758|T191|PT|55020008|SNOMEDCT_US|Follicular lymphoma, grade 2|9691/3
C0079758|T191|PT|277624003|SNOMEDCT_US|Follicular malignant lymphoma - mixed cell type|9691/3
C0079758|T191|SY|277624003|SNOMEDCT_US|Follicular malignant lymphoma - mixed small cleaved and large cell|9691/3
C1301456|T191|SY|702977001|SNOMEDCT_US|Follicular non-Hodgkin lymphoma diffuse follicle center cell sub-type grade 2|9691/3
C1301456|T191|SYGB|702977001|SNOMEDCT_US|Follicular non-Hodgkin lymphoma diffuse follicle centre cell sub-type grade 2|9691/3
C0079758|T191|SY|109971005|SNOMEDCT_US|Follicular non-Hodgkin lymphoma, mixed small cleaved cell and large cell|9691/3
C0079758|T191|SY|188672005|SNOMEDCT_US|Follicular non-Hodgkin mixed small cleaved and large cell lymphoma|9691/3
C1301456|T191|PT|702977001|SNOMEDCT_US|Follicular non-Hodgkin's lymphoma diffuse follicle center cell sub-type grade 2|9691/3
C1301456|T191|PTGB|702977001|SNOMEDCT_US|Follicular non-Hodgkin's lymphoma diffuse follicle centre cell sub-type grade 2|9691/3
C0079758|T191|SY|109971005|SNOMEDCT_US|Follicular non-Hodgkin's lymphoma, mixed small cleaved cell and large cell|9691/3
C0079758|T191|PT|188672005|SNOMEDCT_US|Follicular non-Hodgkin's mixed small cleaved and large cell lymphoma|9691/3
C0079758|T191|SY|55020008|SNOMEDCT_US|Malignant lymphoma, mixed cell type, follicular|9691/3
C0079758|T191|SY|55020008|SNOMEDCT_US|Malignant lymphoma, mixed cell type, nodular|9691/3
C0079758|T191|PT|307636001|SNOMEDCT_US|Malignant lymphoma, mixed lymphocytic-histiocytic, nodular|9691/3
C0079758|T191|SY|55020008|SNOMEDCT_US|Malignant lymphoma, mixed lymphocytic-histiocytic, nodular|9691/3
C0079758|T191|SY|55020008|SNOMEDCT_US|Malignant lymphoma, mixed small cleaved and large cell, follicular|9691/3
C0079758|T191|SY|307636001|SNOMEDCT_US|Reticulolymphosarcoma, follicular|9691/3
C0079758|T191|SY|307636001|SNOMEDCT_US|Reticulolymphosarcoma, nodular|9691/3
C1956130|T191|AB|C82.0|ICD10CM|Follicular lymphoma grade I|9695/3
C1956130|T191|HT|C82.0|ICD10CM|Follicular lymphoma grade I|9695/3
C1956130|T191|ET|D008224|MSH|Follicular Lymphoma, Grade 1|9695/3
C1956130|T191|PEP|D008224|MSH|Lymphoma, Follicular, Grade 1|9695/3
C1956130|T191|PN|NOCODE|MTH|Lymphoma, Follicular, Grade 1|9695/3
C1956130|T191|SY|C3465|NCI|Follicular Small Cleaved Cell Lymphoma|9695/3
C1956130|T191|PT|C3465|NCI|Grade 1 Follicular Lymphoma|9695/3
C1956130|T191|SY|TCGA|NCI|Grade 1 Follicular Lymphoma|9695/3
C1956130|T191|SY|C3465|NCI|Grade I Follicular Lymphoma|9695/3
C1956130|T191|SY|C3465|NCI|Grade I Follicular Small Cleaved Cell Lymphoma|9695/3
C1956130|T191|OP|C3465|NCI|Poorly Differentiated Nodular Lymphocytic Lymphoma|9695/3
C1956130|T191|PT|C3465|NCI_CPTAC|Grade 1 Follicular Lymphoma|9695/3
C1956130|T191|DN|C3465|NCI_CTRP|Grade 1 Follicular Lymphoma|9695/3
C1956130|T191|PT|CDR0000430861|NCI_NCI-GLOSS|grade 1 follicular lymphoma|9695/3
C1956130|T191|SY|CDR0000038316|PDQ|FSC lymphoma|9695/3
C1956130|T191|PT|CDR0000038316|PDQ|grade 1 follicular lymphoma|9695/3
C1956130|T191|SY|CDR0000038316|PDQ|Grade I Follicular Lymphoma|9695/3
C1956130|T191|SY|CDR0000038316|PDQ|grade I follicular small cleaved cell lymphoma|9695/3
C1956130|T191|IS|CDR0000038316|PDQ|Poorly Differentiated Nodular Lymphocytic Lymphoma|9695/3
C1301455|T191|PT|397468001|SNOMEDCT_US|Follicular lymphoma, diffuse follicle center sub-type, grade 1|9695/3
C1301455|T191|PTGB|397468001|SNOMEDCT_US|Follicular lymphoma, diffuse follicle centre sub-type, grade 1|9695/3
C1956130|T191|PT|46744002|SNOMEDCT_US|Follicular lymphoma, grade 1|9695/3
C1301455|T191|SY|702786004|SNOMEDCT_US|Follicular non-Hodgkin lymphoma diffuse follicle center sub-type grade 1|9695/3
C1301455|T191|SYGB|702786004|SNOMEDCT_US|Follicular non-Hodgkin lymphoma diffuse follicle centre sub-type grade 1|9695/3
C1301455|T191|PT|702786004|SNOMEDCT_US|Follicular non-Hodgkin's lymphoma diffuse follicle center sub-type grade 1|9695/3
C1301455|T191|PTGB|702786004|SNOMEDCT_US|Follicular non-Hodgkin's lymphoma diffuse follicle centre sub-type grade 1|9695/3
C0079745|T191|SY|0000034151|CHV|follicular grade 3 lymphoma|9698/3
C0079745|T191|SY|0000015223|CHV|follicular large cell lymphoma|9698/3
C0079745|T191|SY|0000034151|CHV|follicular lymphoma grade 3|9698/3
C0079745|T191|PT|0000034151|CHV|follicular, centroblastic malignant lymphoma|9698/3
C0079745|T191|PT|0000015223|CHV|large cell follicular lymphoma|9698/3
C0079745|T191|PS|C82.2|ICD10|Large cell, follicular|9698/3
C1333846|T191|AB|C82.3|ICD10CM|Follicular lymphoma grade IIIa|9698/3
C1333846|T191|HT|C82.3|ICD10CM|Follicular lymphoma grade IIIa|9698/3
C0079745|T191|PT|MTHU046836|ICPC2ICD10ENG|lymphoma; nodular, histiocytic|9698/3
C0079745|T191|PT|MTHU053413|ICPC2ICD10ENG|nodular; lymphoma, histiocytic|9698/3
C0079745|T191|PT|357226|MEDCIN|follicular malignant lymphoma - large cell|9698/3
C0079745|T191|PT|357185|MEDCIN|malignant follicular lymphoma - centroblastic|9698/3
C0079745|T191|SY|357226|MEDCIN|malignant follicular lymphoma - large cell|9698/3
C0079745|T191|SY|357185|MEDCIN|malignant neoplasm lymphoma follicular - centroblastic|9698/3
C0079745|T191|SY|357226|MEDCIN|malignant neoplasm lymphoma follicular - large cell|9698/3
C0079745|T191|DEV|D008224|MSH|FOLLIC LARGE LYMPHOMA|9698/3
C0079745|T191|PM|D008224|MSH|Follicular Large Cell Lymphoma|9698/3
C0079745|T191|ET|D008224|MSH|Follicular Large-Cell Lymphoma|9698/3
C0079745|T191|PM|D008224|MSH|Follicular Large-Cell Lymphomas|9698/3
C1956131|T191|ET|D008224|MSH|Follicular Lymphoma, Grade 3|9698/3
C0079745|T191|ET|D008224|MSH|Histiocytic Lymphoma, Nodular|9698/3
C0079745|T191|PM|D008224|MSH|Histiocytic Lymphomas, Nodular|9698/3
C0079745|T191|PM|D008224|MSH|Large Cell Lymphoma, Follicular|9698/3
C0079745|T191|ET|D008224|MSH|Large Lymphoid Lymphoma, Nodular|9698/3
C0079745|T191|DEV|D008224|MSH|LARGE LYMPHOMA FOLLIC|9698/3
C0079745|T191|ET|D008224|MSH|Large-Cell Lymphoma, Follicular|9698/3
C0079745|T191|PM|D008224|MSH|Large-Cell Lymphomas, Follicular|9698/3
C0079745|T191|DEV|D008224|MSH|LYMPHOMA FOLLIC LARGE|9698/3
C0079745|T191|DEV|D008224|MSH|LYMPHOMA LARGE FOLLIC|9698/3
C0079745|T191|DEV|D008224|MSH|LYMPHOMA NODULAR LARGE FOLLIC CENTER|9698/3
C0079745|T191|PM|D008224|MSH|Lymphoma, Follicular Large Cell|9698/3
C0079745|T191|ET|D008224|MSH|Lymphoma, Follicular Large-Cell|9698/3
C1956131|T191|PEP|D008224|MSH|Lymphoma, Follicular, Grade 3|9698/3
C0079745|T191|ET|D008224|MSH|Lymphoma, Histiocytic, Nodular|9698/3
C0079745|T191|ET|D008224|MSH|Lymphoma, Large Cell, Follicular|9698/3
C0079745|T191|ET|D008224|MSH|Lymphoma, Large Lymphoid, Nodular|9698/3
C0079745|T191|PEP|D008224|MSH|Lymphoma, Large-Cell, Follicular|9698/3
C0079745|T191|PM|D008224|MSH|Lymphoma, Nodular Histiocytic|9698/3
C0079745|T191|ET|D008224|MSH|Lymphoma, Nodular, Large Follicular Center Cell|9698/3
C0079745|T191|ET|D008224|MSH|Lymphoma, Nodular, Large Follicular Center-Cell|9698/3
C0079745|T191|PM|D008224|MSH|Lymphomas, Follicular Large-Cell|9698/3
C0079745|T191|PM|D008224|MSH|Lymphomas, Nodular Histiocytic|9698/3
C0079745|T191|PM|D008224|MSH|Nodular Histiocytic Lymphoma|9698/3
C0079745|T191|PM|D008224|MSH|Nodular Histiocytic Lymphomas|9698/3
C0079745|T191|DEV|D008224|MSH|NODULAR LARGE FOLLIC CENTER LYMPHOMA|9698/3
C0079745|T191|PM|D008224|MSH|Nodular Large Follicular Center Cell Lymphoma|9698/3
C0079745|T191|ET|D008224|MSH|Nodular Large Follicular Center-Cell Lymphoma|9698/3
C1956131|T191|PN|NOCODE|MTH|Lymphoma, Follicular, Grade 3|9698/3
C0079745|T191|PN|U002379|MTH|Lymphoma, Large-Cell, Follicular|9698/3
C0079745|T191|ET|202.0|MTHICD9|Large cell follicular lymphoma|9698/3
C0079745|T191|ET|200.0|MTHICD9|Lymphoma histiocytic nodular|9698/3
C0079745|T191|ET|200.0|MTHICD9|Malignant lymphoma histiocytic nodular|9698/3
C0079745|T191|SY|C3460|NCI|Follicular Large Cell Lymphoma|9698/3
C0079745|T191|OP|C3460|NCI|Follicular Lymphoma, Predominantly Large Cell|9698/3
C0079745|T191|PT|C3460|NCI|Grade 3 Follicular Lymphoma|9698/3
C0079745|T191|SY|TCGA|NCI|Grade 3 Follicular Lymphoma|9698/3
C1333846|T191|PT|C7191|NCI|Grade 3a Follicular Lymphoma|9698/3
C1333849|T191|PT|C7192|NCI|Grade 3b Follicular Lymphoma|9698/3
C0079745|T191|SY|C3460|NCI|Grade III Follicular Large Cell Lymphoma|9698/3
C0079745|T191|SY|C3460|NCI|Grade III Follicular Lymphoma|9698/3
C0079745|T191|OP|C8994|NCI|Malignant Lymphoma Centroblastic, Follicular|9698/3
C0079745|T191|PT|C8994|NCI|Malignant Lymphoma Centroblastic, Follicular|9698/3
C0079745|T191|OP|C3460|NCI|Nodular Histiocytic Lymphoma|9698/3
C0079745|T191|PT|C3460|NCI_CPTAC|Grade 3 Follicular Lymphoma|9698/3
C1333846|T191|PT|C7191|NCI_CPTAC|Grade 3a Follicular Lymphoma|9698/3
C0079745|T191|DN|C3460|NCI_CTRP|Grade 3 Follicular Lymphoma|9698/3
C0079745|T191|PT|CDR0000044238|NCI_NCI-GLOSS|follicular large cell lymphoma|9698/3
C0079745|T191|PT|CDR0000430863|NCI_NCI-GLOSS|grade 3 follicular lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|FL lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|follicular large cell lymphoma|9698/3
C0079745|T191|PT|CDR0000038381|PDQ|grade 3 follicular lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|grade III follicular large cell lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|grade III follicular lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|histiocytic nodular lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|large cell follicular lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|lymphoma, follicular large cell|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|lymphoma, nodular histiocytic|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|NH lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|NHL|9698/3
C0079745|T191|IS|CDR0000038381|PDQ|nodular histiocytic lymphoma|9698/3
C0079745|T191|SY|CDR0000038381|PDQ|nodular histiocytic lymphoma|9698/3
C0079745|T191|AB|Xa0TX|RCD|Foll malig lymphoma-large cell|9698/3
C0079745|T191|PT|Xa0TX|RCD|Follicular malignant lymphoma - large cell|9698/3
C0079745|T191|AB|XaBBp|RCD|Germinoblastic sarc, follicul|9698/3
C0079745|T191|SY|XaBBp|RCD|Germinoblastic sarcoma, follicular|9698/3
C0079745|T191|AB|Xa0TX|RCD|Malig lymphom-histiocyt, nodul|9698/3
C0079745|T191|AB|Xa0TX|RCD|Malig lymphom-noncleav, follic|9698/3
C0079745|T191|AB|XaBBp|RCD|Malig lyoma,centroblast,foll|9698/3
C0079745|T191|SY|Xa0TX|RCD|Malignant lymphoma - histiocytic, nodular|9698/3
C0079745|T191|SY|Xa0TX|RCD|Malignant lymphoma - non-cleaved, follicular|9698/3
C0079745|T191|PT|XaBBp|RCD|Malignant lymphoma, centroblastic type, follicular|9698/3
C0079745|T191|AB|BBk7.|RCDSY|Mal.lymp,centroblastic,foll|9698/3
C0079745|T191|PT|BBk7.|RCDSY|Malignant lymphoma, centroblastic type, follicular|9698/3
C1956131|T191|PT|40411000|SNOMEDCT_US|Follicular lymphoma, grade 3|9698/3
C0079745|T191|OAP|188673000|SNOMEDCT_US|Follicular malignant lymphoma - large cell|9698/3
C0079745|T191|OAP|277641001|SNOMEDCT_US|Follicular malignant lymphoma - large cell|9698/3
C0079745|T191|OF|188673000|SNOMEDCT_US|Follicular malignant lymphoma - large cell|9698/3
C0079745|T191|SY|307647008|SNOMEDCT_US|Germinoblastic sarcoma, follicular|9698/3
C0079745|T191|OAS|277641001|SNOMEDCT_US|Malignant lymphoma - histiocytic, nodular|9698/3
C0079745|T191|OAS|277641001|SNOMEDCT_US|Malignant lymphoma - non-cleaved, follicular|9698/3
C0079745|T191|PT|307647008|SNOMEDCT_US|Malignant lymphoma, centroblastic type, follicular|9698/3
C0079745|T191|OAP|80358008|SNOMEDCT_US|Malignant lymphoma, centroblastic, follicular|9698/3
C0079745|T191|SY|40411000|SNOMEDCT_US|Malignant lymphoma, centroblastic, follicular|9698/3
C0079745|T191|IS|80358008|SNOMEDCT_US|Malignant lymphoma, centroblastic, follicular -RETIRED-|9698/3
C0079745|T191|OF|80358008|SNOMEDCT_US|Malignant lymphoma, centroblastic, follicular -RETIRED-|9698/3
C0079745|T191|SY|40411000|SNOMEDCT_US|Malignant lymphoma, histiocytic, nodular|9698/3
C0079745|T191|SY|40411000|SNOMEDCT_US|Malignant lymphoma, large cell, follicular|9698/3
C0079745|T191|IS|40411000|SNOMEDCT_US|Malignant lymphoma, large cell, follicular, NOS|9698/3
C0079745|T191|SY|40411000|SNOMEDCT_US|Malignant lymphoma, large cell, noncleaved, follicular|9698/3
C0079745|T191|SY|40411000|SNOMEDCT_US|Malignant lymphoma, large cleaved cell, follicular|9698/3
C0079745|T191|SY|40411000|SNOMEDCT_US|Malignant lymphoma, noncleaved, follicular|9698/3
C0079745|T191|IS|40411000|SNOMEDCT_US|Malignant lymphoma, noncleaved, follicular, NOS|9698/3
C0242647|T191|SY|0000024900|CHV|malt lymphoma|9699/3
C0242647|T191|PT|0000036642|CHV|maltoma|9699/3
C0242647|T191|SY|0000036642|CHV|maltomas|9699/3
C0242647|T191|SY|0000024900|CHV|marginal zone b cell lymphoma|9699/3
C0242647|T191|SY|0000024900|CHV|marginal zone b-cell lymphoma|9699/3
C0242647|T191|SY|0000024900|CHV|marginal zone lymphoma|9699/3
C0242647|T191|SY|0000024900|CHV|nodal marginal zone lymphoma|9699/3
C0242647|T191|AB|C88.4|ICD10CM|Extrnod mrgnl zn B-cell lymph of mucosa-assoc lymphoid tiss|9699/3
C0855139|T191|ET|C83.0|ICD10CM|Nodal marginal zone lymphoma|9699/3
C1367654|T191|HT|200.3|ICD9CM|Marginal zone lymphoma|9699/3
C0855139|T191|PT|MTHU009822|ICPC2ICD10ENG|B-cell; lymphoma, monocytoid|9699/3
C0855139|T191|PT|MTHU046739|ICPC2ICD10ENG|lymphoma; B-cell, monocytoid|9699/3
C0855139|T191|PT|MTHU046827|ICPC2ICD10ENG|lymphoma; monocytoid B-cell|9699/3
C0855139|T191|PT|MTHU050297|ICPC2ICD10ENG|monocytoid B-cell; lymphoma|9699/3
C0242647|T191|LLT|10060707|MDR|MALT lymphoma|9699/3
C1367654|T191|LLT|10076596|MDR|Marginal zone lymphoma|9699/3
C1367654|T191|PT|10076596|MDR|Marginal zone lymphoma|9699/3
C0855139|T191|LLT|10029460|MDR|Nodal marginal zone B-cell lymphoma|9699/3
C0855139|T191|PT|10029460|MDR|Nodal marginal zone B-cell lymphoma|9699/3
C0855139|T191|LLT|10029462|MDR|Nodal marginal zone B-cell lymphoma NOS|9699/3
C0855139|T191|HT|10029461|MDR|Nodal marginal zone B-cell lymphomas|9699/3
C0242647|T191|PT|338555|MEDCIN|extranodal marginal zone B-cell lymphoma of mucosa associated lymphoid tissue|9699/3
C0855139|T191|SY|355314|MEDCIN|malignant neoplasm lymphoma b-cell low grade diffuse monocytoid|9699/3
C1275321|T191|SY|357442|MEDCIN|malignant neoplasm lymphoma b-cell primary cutaneous marginal zone|9699/3
C1367654|T191|PT|271575|MEDCIN|marginal zone B-cell lymphoma|9699/3
C0242647|T191|SY|355326|MEDCIN|marginal zone b-cell lymphoma mucosa-associated|9699/3
C0242647|T191|SY|338555|MEDCIN|marginal zone b-cell lymphoma of mucosa associated lymphoid tissue extranodal|9699/3
C0242647|T191|PT|272058|MEDCIN|marginal zone B-cell lymphoma of reticuloendothelial system|9699/3
C1367654|T191|PT|312615|MEDCIN|marginal zone lymphoma|9699/3
C0855139|T191|PT|355314|MEDCIN|Monocytoid B-cell lymphoma|9699/3
C0242647|T191|PT|355326|MEDCIN|Mucosa-associated lymphoma|9699/3
C0855139|T191|PT|312618|MEDCIN|nodal marginal zone B-cell lymphoma|9699/3
C1275321|T191|PT|357442|MEDCIN|Primary cutaneous marginal zone B-cell lymphoma|9699/3
C0242647|T191|DEV|D018442|MSH|LYMPHOMA MALT|9699/3
C0242647|T191|DEV|D018442|MSH|LYMPHOMA MUCOSA ASSOC LYMPHOID TISSUE|9699/3
C0242647|T191|PM|D018442|MSH|Lymphoma of Mucosa Associated Lymphoid Tissue|9699/3
C0242647|T191|ET|D018442|MSH|Lymphoma of Mucosa-Associated Lymphoid Tissue|9699/3
C0242647|T191|MH|D018442|MSH|Lymphoma, B-Cell, Marginal Zone|9699/3
C0242647|T191|PM|D018442|MSH|Lymphoma, MALT|9699/3
C0242647|T191|PM|D018442|MSH|Lymphoma, Mucosa Associated Lymphoid Tissue|9699/3
C0242647|T191|ET|D018442|MSH|Lymphoma, Mucosa-Associated Lymphoid Tissue|9699/3
C0242647|T191|PM|D018442|MSH|Lymphomas, MALT|9699/3
C0242647|T191|ET|D018442|MSH|MALT Lymphoma|9699/3
C0242647|T191|PM|D018442|MSH|MALT Lymphomas|9699/3
C0242647|T191|PM|D018442|MSH|Marginal Zone B Cell Lymphoma|9699/3
C0242647|T191|ET|D018442|MSH|Marginal Zone B-Cell Lymphoma|9699/3
C0242647|T191|DEV|D018442|MSH|MUCOSA ASSOC LYMPHOID TISSUE LYMPHOMA|9699/3
C0242647|T191|PM|D018442|MSH|Mucosa Associated Lymphoid Tissue Lymphoma|9699/3
C0242647|T191|ET|D018442|MSH|Mucosa-Associated Lymphoid Tissue Lymphoma|9699/3
C1367654|T191|PN|NOCODE|MTH|Marginal Zone B-Cell Lymphoma|9699/3
C0855139|T191|PN|NOCODE|MTH|Monocytoid B-cell lymphoma|9699/3
C0242647|T191|PN|NOCODE|MTH|Mucosa-Associated Lymphoid Tissue Lymphoma|9699/3
C0855139|T191|ET|200.3|MTHICD9|Nodal marginal zone B-cell lymphoma|9699/3
C2698751|T191|SY|C80299|NCI|Childhood Nodal Marginal Zone Lymphoma|9699/3
C0242647|T191|SY|C3898|NCI|Extranodal Marginal Zone B-Cell Lymphoma of Mucosa-Associated Lymphoid Tissue|9699/3
C0242647|T191|SY|TCGA|NCI|Extranodal Marginal Zone Lymphoma of Mucosa-Associated Lymphoid Tissue|9699/3
C0242647|T191|PT|C3898|NCI|Extranodal Marginal Zone Lymphoma of Mucosa-Associated Lymphoid Tissue|9699/3
C0242647|T191|OP|C3898|NCI|Immunocytoma|9699/3
C0242647|T191|SY|C3898|NCI|MALT Lymphoma|9699/3
C0242647|T191|SY|C3898|NCI|MALToma|9699/3
C1367654|T191|SY|C4341|NCI|Marginal Zone B-Cell Lymphoma|9699/3
C1367654|T191|PT|C4341|NCI|Marginal Zone Lymphoma|9699/3
C0855139|T191|SY|C8863|NCI|Monocytoid B-Cell Lymphoma|9699/3
C0242647|T191|SY|C3898|NCI|Mucosa-Associated Lymphoid Tissue Lymphoma|9699/3
C1367654|T191|AB|C4341|NCI|MZBCL|9699/3
C1367654|T191|AB|C4341|NCI|MZL|9699/3
C0855139|T191|SY|C8863|NCI|Nodal Marginal Zone B-Cell Lymphoma|9699/3
C0855139|T191|SY|TCGA|NCI|Nodal Marginal Zone Lymphoma|9699/3
C0855139|T191|PT|C8863|NCI|Nodal Marginal Zone Lymphoma|9699/3
C2698751|T191|PT|C80299|NCI|Pediatric Nodal Marginal Zone Lymphoma|9699/3
C0242647|T191|PT|C3898|NCI_CPTAC|Extranodal Marginal Zone Lymphoma of Mucosa-Associated Lymphoid Tissue|9699/3
C1367654|T191|PT|C4341|NCI_CPTAC|Marginal Zone Lymphoma|9699/3
C0242647|T191|SY|10015822|NCI_CTEP-SDC|MALT-lymphoma|9699/3
C0855139|T191|SY|10029462|NCI_CTEP-SDC|Nodal marginal zone B-cell lymph.|9699/3
C0855139|T191|PT|10029462|NCI_CTEP-SDC|Nodal marginal zone B-cell lymphoma|9699/3
C0242647|T191|DN|C3898|NCI_CTRP|Extranodal Marginal Zone Lymphoma of Mucosa-Associated Lymphoid Tissue|9699/3
C1367654|T191|DN|C4341|NCI_CTRP|Marginal Zone Lymphoma|9699/3
C0855139|T191|DN|C8863|NCI_CTRP|Nodal Marginal Zone Lymphoma|9699/3
C0242647|T191|PT|CDR0000045774|NCI_NCI-GLOSS|MALT lymphoma|9699/3
C1367654|T191|PT|CDR0000562554|NCI_NCI-GLOSS|marginal zone B-cell lymphoma|9699/3
C1367654|T191|PT|CDR0000543124|NCI_NCI-GLOSS|marginal zone lymphoma|9699/3
C0242647|T191|PT|CDR0000044437|NCI_NCI-GLOSS|mucosa-associated lymphoid tissue lymphoma|9699/3
C1367654|T191|PT|CDR0000562555|NCI_NCI-GLOSS|MZL|9699/3
C2698751|T191|PT|C80299|NCI_NICHD|Childhood Nodal Marginal Zone Lymphoma|9699/3
C2698751|T191|SY|C80299|NCI_NICHD|Pediatric Nodal Marginal Zone Lymphoma|9699/3
C0242647|T191|PT|CDR0000372812|PDQ|extranodal marginal zone B-cell lymphoma of mucosa-associated lymphoid tissue|9699/3
C0242647|T191|IS|CDR0000372812|PDQ|immunocytoma|9699/3
C0242647|T191|SY|CDR0000042230|PDQ|lymphoid tissue, mucosa-associated|9699/3
C0242647|T191|AB|CDR0000042230|PDQ|MALT|9699/3
C0242647|T191|SY|CDR0000372812|PDQ|MALT lymphoma|9699/3
C0242647|T191|SY|CDR0000372812|PDQ|MALToma|9699/3
C1367654|T191|SY|CDR0000371894|PDQ|marginal zone B-cell lymphoma|9699/3
C1367654|T191|ET|CDR0000371894|PDQ|Marginal zone lymphoma|9699/3
C1367654|T191|PT|CDR0000371894|PDQ|marginal zone lymphoma|9699/3
C0855139|T191|SY|CDR0000372811|PDQ|monocytoid B-cell lymphoma|9699/3
C0242647|T191|OP|CDR0000042230|PDQ|mucosa-associated lymphoid tissue|9699/3
C0242647|T191|SY|CDR0000372812|PDQ|mucosa-associated lymphoid tissue lymphoma|9699/3
C1367654|T191|AB|CDR0000371894|PDQ|MZBCL|9699/3
C1367654|T191|AB|CDR0000371894|PDQ|MZL|9699/3
C0855139|T191|PT|CDR0000372811|PDQ|nodal marginal zone B-cell lymphoma|9699/3
C0242647|T191|SY|Xa0T8|RCD|Maltoma|9699/3
C0855139|T191|PT|Xa0T9|RCD|Monocytoid B-cell lymphoma|9699/3
C0242647|T191|PT|Xa0T8|RCD|Mucosa-associated lymphoma|9699/3
C0855139|T191|OP|BBv0.|RCDSY|Monocytoid B-cell lymphoma|9699/3
C0855139|T191|OP|BBm9.|RCDSY|Monocytoid B-cell lymphoma|9699/3
C0242647|T191|PT|397350003|SNOMEDCT_US|Extranodal marginal zone B-cell lymphoma of mucosa-associated lymphoid tissue|9699/3
C0242647|T191|SY|445269007|SNOMEDCT_US|Extranodal marginal zone B-cell lymphoma of mucosa-associated lymphoid tissue|9699/3
C0242647|T191|SY|128803008|SNOMEDCT_US|MALT lymphoma|9699/3
C0242647|T191|SY|277622004|SNOMEDCT_US|Maltoma|9699/3
C1367654|T191|PT|128803008|SNOMEDCT_US|Marginal zone B-cell lymphoma|9699/3
C1367654|T191|OAP|103683000|SNOMEDCT_US|Marginal zone lymphoma|9699/3
C1367654|T191|SY|128803008|SNOMEDCT_US|Marginal zone lymphoma|9699/3
C1367654|T191|PT|447100004|SNOMEDCT_US|Marginal zone lymphoma|9699/3
C1367654|T191|IS|103683000|SNOMEDCT_US|Marginal zone lymphoma -RETIRED-|9699/3
C1367654|T191|OF|103683000|SNOMEDCT_US|Marginal zone lymphoma -RETIRED-|9699/3
C1367654|T191|IS|103683000|SNOMEDCT_US|Marginal zone lymphoma, NOS|9699/3
C0855139|T191|PT|277623009|SNOMEDCT_US|Monocytoid B-cell lymphoma|9699/3
C0855139|T191|SY|128803008|SNOMEDCT_US|Monocytoid B-cell lymphoma|9699/3
C0855139|T191|OAP|13204007|SNOMEDCT_US|Monocytoid B-cell lymphoma|9699/3
C0855139|T191|IS|13204007|SNOMEDCT_US|Monocytoid B-cell lymphoma -RETIRED-|9699/3
C0855139|T191|OF|13204007|SNOMEDCT_US|Monocytoid B-cell lymphoma -RETIRED-|9699/3
C0242647|T191|PT|277622004|SNOMEDCT_US|Mucosa-associated lymphoma|9699/3
C0242647|T191|SY|128803008|SNOMEDCT_US|Mucosal-associated lymphoid tissue lymphoma|9699/3
C0855139|T191|PT|726721002|SNOMEDCT_US|Nodal marginal zone B-cell lymphoma|9699/3
C0855139|T191|PT|397349003|SNOMEDCT_US|Nodal marginal zone B-cell lymphoma|9699/3
C0242647|T191|SY|128803008|SNOMEDCT_US|Nodal marginal zone lymphoma|9699/3
C2698751|T191|PTGB|733860007|SNOMEDCT_US|Paediatric nodal marginal zone lymphoma|9699/3
C2698751|T191|PT|733860007|SNOMEDCT_US|Pediatric nodal marginal zone lymphoma|9699/3
C1275321|T191|PT|420028002|SNOMEDCT_US|Primary cutaneous marginal zone B-cell lymphoma|9699/3
C1275321|T191|PT|404140004|SNOMEDCT_US|Primary cutaneous marginal zone B-cell lymphoma|9699/3
C1275321|T191|SY|404140004|SNOMEDCT_US|SALT type B-cell lymphoma|9699/3
C1275321|T191|SY|404140004|SNOMEDCT_US|Skin-associated lymphoid tissue type B-cell lymphoma|9699/3
C0026948|T191|PT|0045940|CCPSS|MYCOSIS FUNGOIDES|9700/3
C0026948|T191|SY|0000008397|CHV|mf|9700/3
C0026948|T191|PT|0000008397|CHV|mycosis fungoides|9700/3
C0026948|T191|PT|U000454|COSTAR|MYCOSIS FUNGOIDES|9700/3
C0026948|T191|PT|2004-7126|CSP|mycosis fungoides lymphoma|9700/3
C0026948|T191|SY|NOCODE|DXP|GRANULOMA, FUNGOIDES|9700/3
C0026948|T191|DI|U001231|DXP|MYCOSIS FUNGOIDES|9700/3
C0026948|T191|PT|C84.0|ICD10|Mycosis fungoides|9700/3
C0026948|T191|HT|C84.0|ICD10CM|Mycosis fungoides|9700/3
C0026948|T191|AB|C84.0|ICD10CM|Mycosis fungoides|9700/3
C0026948|T191|PT|C84.00|ICD10CM|Mycosis fungoides, unspecified site|9700/3
C0026948|T191|AB|C84.00|ICD10CM|Mycosis fungoides, unspecified site|9700/3
C0026948|T191|HT|202.1|ICD9CM|Mycosis fungoides|9700/3
C0026948|T191|PT|MTHU050796|ICPC2ICD10ENG|Mycosis fungoides|9700/3
C0026948|T191|PT|U003084|LCH|Mycosis fungoides|9700/3
C0026948|T191|PT|sh85089199|LCH_NW|Mycosis fungoides|9700/3
C0026948|T191|HT|10028484|MDR|Mycoses fungoides|9700/3
C0026948|T191|LLT|10028483|MDR|Mycosis fungoides|9700/3
C0026948|T191|LLT|10028500|MDR|Mycosis fungoides NOS|9700/3
C1627767|T047|PT|350537|MEDCIN|Follicular mucinosis type mycosis fungoides|9700/3
C0026948|T191|PT|31604|MEDCIN|mycosis fungoides|9700/3
C1367970|T191|PT|350548|MEDCIN|Pagetoid reticulosis|9700/3
C1367970|T191|PM|D056267|MSH|Disease, Woringer Kolopp|9700/3
C1367970|T191|PM|D056267|MSH|Disease, Woringer-Kolopp|9700/3
C1367970|T191|PM|D056267|MSH|Kolopp Disease, Woringer|9700/3
C0026948|T191|MH|D009182|MSH|Mycosis Fungoides|9700/3
C1367970|T191|PM|D056267|MSH|Pagetoid Reticuloses|9700/3
C1367970|T191|MH|D056267|MSH|Pagetoid Reticulosis|9700/3
C1367970|T191|PM|D056267|MSH|Reticuloses, Pagetoid|9700/3
C1367970|T191|PM|D056267|MSH|Reticulosis, Pagetoid|9700/3
C1367970|T191|ET|D056267|MSH|Woringer Kolopp Disease|9700/3
C1367970|T191|ET|D056267|MSH|Woringer-Kolopp Disease|9700/3
C0026948|T191|PN|U002093|MTH|Mycosis Fungoides|9700/3
C1367970|T191|PN|NOCODE|MTH|Pagetoid reticulosis|9700/3
C1627767|T047|SY|C35685|NCI|Follicular Mycosis Fungoides|9700/3
C1627767|T047|PT|C35685|NCI|Folliculotropic Mycosis Fungoides|9700/3
C0026948|T191|AB|C3246|NCI|MF|9700/3
C0026948|T191|PT|C3246|NCI|Mycosis Fungoides|9700/3
C0026948|T191|SY|TCGA|NCI|Mycosis Fungoides|9700/3
C1627767|T047|SY|C35685|NCI|Mycosis Fungoides-Associated Follicular Mucinosis|9700/3
C1367970|T191|PT|C35794|NCI|Pagetoid Reticulosis|9700/3
C0026948|T191|PT|C3246|NCI_CPTAC|Mycosis Fungoides|9700/3
C0026948|T191|SY|10028500|NCI_CTEP-SDC|CTCL/ Mycosis fungoides|9700/3
C0026948|T191|PT|10028500|NCI_CTEP-SDC|Cutaneous T-cell lymphoma/Mycosis fungoides|9700/3
C0026948|T191|DN|C3246|NCI_CTRP|Mycosis Fungoides|9700/3
C0026948|T191|PT|CDR0000045794|NCI_NCI-GLOSS|mycosis fungoides|9700/3
C0026948|T191|SY|CDR0000043725|PDQ|mycosis fungoides|9700/3
C0026948|T191|SY|B621.|RCD|MF - Mycosis fungoides|9700/3
C0026948|T191|PT|B621.|RCD|Mycosis fungoides|9700/3
C0026948|T191|OP|B621z|RCD|Mycosis fungoides NOS|9700/3
C0026948|T191|OP|B6210|RCD|Mycosis fungoides of unspecified site|9700/3
C0026948|T191|OA|B6210|RCD|Mycosis fungoides-unspec. site|9700/3
C0026948|T191|PT|BBl..|RCDSY|Mycosis fungoides|9700/3
C0026948|T191|OP|BBlz.|RCDSY|Mycosis fungoides NOS|9700/3
C1627767|T047|PT|404109006|SNOMEDCT_US|Follicular mucinosis type mycosis fungoides|9700/3
C1627767|T047|PT|418628003|SNOMEDCT_US|Follicular mycosis fungoides|9700/3
C1627767|T047|SY|404109006|SNOMEDCT_US|Folliculotropic mycosis fungoides|9700/3
C0026948|T191|SY|118618005|SNOMEDCT_US|MF - Mycosis fungoides|9700/3
C0026948|T191|SY|118618005|SNOMEDCT_US|Mycosis fungoides|9700/3
C0026948|T191|PT|90120004|SNOMEDCT_US|Mycosis fungoides|9700/3
C0026948|T191|OAP|188628007|SNOMEDCT_US|Mycosis fungoides NOS|9700/3
C0026948|T191|OAP|188618003|SNOMEDCT_US|Mycosis fungoides of unspecified site|9700/3
C1367970|T191|PT|404119000|SNOMEDCT_US|Pagetoid reticulosis|9700/3
C1367970|T191|PT|419386004|SNOMEDCT_US|Pagetoid reticulosis|9700/3
C1367970|T191|SY|90120004|SNOMEDCT_US|Pagetoid reticulosis|9700/3
C0026948|T191|IT|1110|WHO|MYCOSIS FUNGOIDES|9700/3
C0036920|T191|PT|0000011288|CHV|sezary syndrome|9701/3
C0036920|T191|SY|0000011288|CHV|sezary's disease|9701/3
C0036920|T191|SY|0000011288|CHV|sezary's syndrome|9701/3
C0036920|T191|PT|NOCODE|COSTAR|Sezary Syndrome|9701/3
C0036920|T191|ET|2004-7126|CSP|Sezary syndrome|9701/3
C0036920|T191|SY|NOCODE|DXP|RETICULOSIS SYNDROME, SEZARY|9701/3
C0036920|T191|DI|U001733|DXP|SEZARY SYNDROME|9701/3
C0036920|T191|PT|C84.1|ICD10|Sezary's disease|9701/3
C0036920|T191|AB|C84.1|ICD10CM|Sezary disease|9701/3
C0036920|T191|HT|C84.1|ICD10CM|Sézary disease|9701/3
C0036920|T191|AB|C84.10|ICD10CM|Sezary disease, unspecified site|9701/3
C0036920|T191|PT|C84.10|ICD10CM|Sézary disease, unspecified site|9701/3
C0036920|T191|HT|202.2|ICD9CM|Sezary's disease|9701/3
C0036920|T191|PT|MTHU064372|ICPC2ICD10ENG|reticulosis; Sézary|9701/3
C0036920|T191|PT|MTHU067628|ICPC2ICD10ENG|Sézary|9701/3
C0036920|T191|PT|MTHU067629|ICPC2ICD10ENG|Sézary; reticulosis|9701/3
C0036920|T191|LLT|10040493|MDR|Sezary syndrome|9701/3
C0036920|T191|LLT|10040500|MDR|Sezary's disease|9701/3
C0036920|T191|LLT|10040516|MDR|Sezary's syndrome|9701/3
C0036920|T191|PT|31605|MEDCIN|Sezary syndrome|9701/3
C0036920|T191|ET|D012751|MSH|Erythroderma, Sezary|9701/3
C0036920|T191|PM|D012751|MSH|Lymphoma, Sezary's|9701/3
C0036920|T191|PM|D012751|MSH|Sezary Erythroderma|9701/3
C0036920|T191|PM|D012751|MSH|Sezary Lymphoma|9701/3
C0036920|T191|MH|D012751|MSH|Sezary Syndrome|9701/3
C0036920|T191|ET|D012751|MSH|Sezary's Lymphoma|9701/3
C0036920|T191|PM|D012751|MSH|Sezarys Lymphoma|9701/3
C0036920|T191|PM|D012751|MSH|Syndrome, Sezary|9701/3
C0036920|T191|PN|U002240|MTH|Sezary Syndrome|9701/3
C0036920|T191|PT|C3366|NCI|Sezary Syndrome|9701/3
C0036920|T191|SY|TCGA|NCI|Sezary Syndrome|9701/3
C0036920|T191|SY|C3366|NCI|Sézary Syndrome|9701/3
C0036920|T191|SY|C3366|NCI|Sezary's Disease|9701/3
C0036920|T191|PT|C3366|NCI_CPTAC|Sezary Syndrome|9701/3
C0036920|T191|SY|10011677|NCI_CTEP-SDC|CTCL / Sezary syndrome|9701/3
C0036920|T191|PT|10011677|NCI_CTEP-SDC|Cutaneous T-cell lymphoma/Sezary syndrome|9701/3
C0036920|T191|DN|C3366|NCI_CTRP|Sezary Syndrome|9701/3
C0036920|T191|PT|CDR0000045878|NCI_NCI-GLOSS|Sezary syndrome|9701/3
C0036920|T191|SY|CDR0000043725|PDQ|Sezary syndrome|9701/3
C0036920|T191|ET|CDR0000043725|PDQ|Sezary syndrome|9701/3
C0036920|T191|PT|B622.|RCD|Sezary's disease|9701/3
C0036920|T191|OP|B622z|RCD|Sezary's disease NOS|9701/3
C0036920|T191|OP|B6220|RCD|Sezary's disease of unspecified site|9701/3
C0036920|T191|OA|B6220|RCD|Sezary's disease-unspec. site|9701/3
C0036920|T191|OP|BBl1.|RCDSY|Sezary's disease|9701/3
C0036920|T191|SY|4950009|SNOMEDCT_US|Sézary disease|9701/3
C0036920|T191|SY|118611004|SNOMEDCT_US|Sézary disease|9701/3
C0036920|T191|PT|4950009|SNOMEDCT_US|Sezary syndrome|9701/3
C0036920|T191|SY|118611004|SNOMEDCT_US|Sezary's disease|9701/3
C0036920|T191|SY|4950009|SNOMEDCT_US|Sezary's disease|9701/3
C0036920|T191|IS|188638002|SNOMEDCT_US|Sezary's disease NOS|9701/3
C0036920|T191|OAP|188638002|SNOMEDCT_US|Sézary's disease NOS|9701/3
C0036920|T191|OAP|188629004|SNOMEDCT_US|Sézary's disease of unspecified site|9701/3
C0036920|T191|OAS|188629004|SNOMEDCT_US|Sezary's disease of unspecified site|9701/3
C0036920|T191|IS|4950009|SNOMEDCT_US|Sezary's syndrome|9701/3
C0036920|T191|SY|4950009|SNOMEDCT_US|Sézary's syndrome|9701/3
C0079774|T191|SY|0000015231|CHV|cell lymphomas peripheral t|9702/3
C0079774|T191|SY|0000015231|CHV|peripheral t cell lymphoma|9702/3
C0079774|T191|SY|0000015231|CHV|peripheral t-cell lymphoma|9702/3
C0079774|T191|PT|C84.4|ICD10|Peripheral T-cell lymphoma|9702/3
C1332078|T191|AB|C84.7|ICD10CM|Anaplastic large cell lymphoma, ALK-negative|9702/3
C1332078|T191|HT|C84.7|ICD10CM|Anaplastic large cell lymphoma, ALK-negative|9702/3
C0079774|T191|AB|C84|ICD10CM|Mature T/NK-cell lymphomas|9702/3
C0079774|T191|HT|C84|ICD10CM|Mature T/NK-cell lymphomas|9702/3
C0079774|T191|AB|C84.9|ICD10CM|Mature T/NK-cell lymphomas, unspecified|9702/3
C0079774|T191|HT|C84.9|ICD10CM|Mature T/NK-cell lymphomas, unspecified|9702/3
C0079774|T191|HT|202.7|ICD9CM|Peripheral T-cell lymphoma|9702/3
C0079774|T191|PT|MTHU046846|ICPC2ICD10ENG|lymphoma; peripheral T-cell|9702/3
C0079774|T191|PT|MTHU046859|ICPC2ICD10ENG|lymphoma; T-cell, peripheral|9702/3
C0079774|T191|PT|MTHU058747|ICPC2ICD10ENG|peripheral; T-cell lymphoma|9702/3
C0079774|T191|PT|MTHU073542|ICPC2ICD10ENG|T-cell; lymphoma, peripheral|9702/3
C0079774|T191|LLT|10034623|MDR|Peripheral T-cell lymphoma unspecified|9702/3
C0079774|T191|PT|10034623|MDR|Peripheral T-cell lymphoma unspecified|9702/3
C0079774|T191|LLT|10034624|MDR|Peripheral T-cell lymphoma unspecified NOS|9702/3
C1332078|T191|PT|333226|MEDCIN|ALK-negative anaplastic large cell lymphoma|9702/3
C1332078|T191|SY|333226|MEDCIN|lymphoma anaplastic large cell ALK-negative|9702/3
C0079774|T191|SY|338146|MEDCIN|malignant neoplasm lymphoma mature nk/t-cell|9702/3
C0079774|T191|PT|338146|MEDCIN|mature NK/T-cell lymphoma|9702/3
C0079774|T191|PT|312907|MEDCIN|mature T-cell lymphoma|9702/3
C0079774|T191|PM|D016411|MSH|Lymphoma, Peripheral T-Cell|9702/3
C0079774|T191|ET|D016411|MSH|Lymphoma, T Cell, Peripheral|9702/3
C0079774|T191|MH|D016411|MSH|Lymphoma, T-Cell, Peripheral|9702/3
C0079774|T191|PM|D016411|MSH|Lymphomas, Peripheral T-Cell|9702/3
C0079774|T191|PM|D016411|MSH|Peripheral T Cell Lymphoma|9702/3
C0079774|T191|ET|D016411|MSH|Peripheral T-Cell Lymphoma|9702/3
C0079774|T191|PM|D016411|MSH|Peripheral T-Cell Lymphomas|9702/3
C0079774|T191|PM|D016411|MSH|T Cell Lymphoma, Peripheral|9702/3
C0079774|T191|ET|D016411|MSH|T-Cell Lymphoma, Peripheral|9702/3
C0079774|T191|PM|D016411|MSH|T-Cell Lymphomas, Peripheral|9702/3
C0079774|T191|PN|NOCODE|MTH|Peripheral T-Cell Lymphoma|9702/3
C1332078|T191|AB|C37194|NCI|ALCL, ALK-|9702/3
C1332078|T191|SY|C37194|NCI|ALK-Negative Anaplastic Large Cell Lymphoma|9702/3
C1332078|T191|PT|C37194|NCI|Anaplastic Large Cell Lymphoma, ALK-Negative|9702/3
C2700204|T191|PT|C80375|NCI|Follicular T-Cell Lymphoma|9702/3
C2700204|T191|SY|C80375|NCI|Follicular Variant Peripheral T-Cell Lymphoma|9702/3
C2700204|T191|AB|C80375|NCI|FTCL|9702/3
C0079774|T191|SY|C3468|NCI|Mature T-and NK-Cell Lymphoma|9702/3
C0079774|T191|SY|C3468|NCI|Mature T-Cell and NK-Cell Lymphoma|9702/3
C0079774|T191|PT|C3468|NCI|Mature T-Cell and NK-Cell Non-Hodgkin Lymphoma|9702/3
C0079774|T191|SY|C3468|NCI|Mature T-Cell and NK-Cell Non-Hodgkin's Lymphoma|9702/3
C0079774|T191|SY|C3468|NCI|Mature T-Cell Non-Hodgkin's Lymphoma|9702/3
C4528209|T191|SY|C139011|NCI|Nodal Peripheral T-Cell Lymphoma with T Follicular Helper Phenotype|9702/3
C4528209|T191|PT|C139011|NCI|Nodal Peripheral T-Cell Lymphoma with TFH Phenotype|9702/3
C4528209|T191|SY|C139011|NCI|Nodal PTCL with T Follicular Helper Phenotype|9702/3
C4528209|T191|SY|C139011|NCI|Nodal PTCL with TFH Phenotype|9702/3
C0079774|T191|SY|C3468|NCI|Peripheral T-Cell Lymphoma|9702/3
C0079774|T191|SY|C4340|NCI|Peripheral T-Cell Lymphoma, NOS|9702/3
C0079774|T191|PT|C4340|NCI|Peripheral T-Cell Lymphoma, Not Otherwise Specified|9702/3
C0079774|T191|SY|TCGA|NCI|Peripheral T-Cell Lymphoma, Not Otherwise Specified|9702/3
C0079774|T191|AB|C3468|NCI|PTCL|9702/3
C1332078|T191|PT|C37194|NCI_CPTAC|Anaplastic Large Cell Lymphoma, ALK-Negative|9702/3
C0079774|T191|PT|C3468|NCI_CPTAC|Mature T-Cell and NK-Cell Non-Hodgkin Lymphoma|9702/3
C0079774|T191|PT|C4340|NCI_CPTAC|Peripheral T-Cell Lymphoma, Not Otherwise Specified|9702/3
C0079774|T191|PT|10034624|NCI_CTEP-SDC|Peripheral T-cell lymphoma, NOS|9702/3
C0079774|T191|DN|C3468|NCI_CTRP|Mature T-Cell and NK-Cell Non-Hodgkin Lymphoma|9702/3
C0079774|T191|PT|CDR0000393800|NCI_NCI-GLOSS|mature T-cell lymphoma|9702/3
C0079774|T191|PT|CDR0000405873|NCI_NCI-GLOSS|peripheral T-cell lymphoma|9702/3
C0079774|T191|SY|CDR0000641396|PDQ|peripheral T-cell lymphoma, NOS|9702/3
C0079774|T191|PT|CDR0000641396|PDQ|peripheral T-cell lymphoma, not otherwise specified|9702/3
C0079774|T191|PT|Xa0Th|RCD|Peripheral T-cell lymphoma|9702/3
C0079774|T191|OA|BBm5.|RCDSY|Peripheral T-cell lymphoma|9702/3
C0079774|T191|OP|BBm5.|RCDSY|Peripheral T-cell lymphoma NOS|9702/3
C1332078|T191|PT|448212009|SNOMEDCT_US|Anaplastic large cell lymphoma, ALK negative|9702/3
C1332078|T191|SY|448212009|SNOMEDCT_US|Anaplastic lymphoma kinase negative anaplastic large cell lymphoma|9702/3
C2700204|T191|PT|784551004|SNOMEDCT_US|Follicular T-cell lymphoma|9702/3
C1282453|T191|PT|314927000|SNOMEDCT_US|High grade T-cell lymphoma morphology|9702/3
C1282456|T191|PT|314930007|SNOMEDCT_US|Low grade T-cell lymphoma morphology|9702/3
C0079774|T191|SY|3172003|SNOMEDCT_US|Mature T-cell lymphoma|9702/3
C4528209|T191|PT|784296005|SNOMEDCT_US|Nodal peripheral T-cell lymphoma with T follicular helper phenotype|9702/3
C0079774|T191|PT|3172003|SNOMEDCT_US|Peripheral T-cell lymphoma|9702/3
C0079774|T191|OAP|188688005|SNOMEDCT_US|Peripheral T-cell lymphoma|9702/3
C0079774|T191|SY|109977009|SNOMEDCT_US|Peripheral T-cell lymphoma|9702/3
C0079774|T191|OF|188688005|SNOMEDCT_US|Peripheral T-cell lymphoma|9702/3
C0079774|T191|SY|3172003|SNOMEDCT_US|Peripheral T-cell lymphoma unspecified|9702/3
C0079774|T191|SY|3172003|SNOMEDCT_US|Peripheral T-cell lymphoma, no ICD-O subtype|9702/3
C0079774|T191|SY|3172003|SNOMEDCT_US|Peripheral T-cell lymphoma, no International Classification of Diseases for Oncology subtype|9702/3
C0079774|T191|IS|3172003|SNOMEDCT_US|Peripheral T-cell lymphoma, NOS|9702/3
C1282452|T191|PT|314926009|SNOMEDCT_US|T-cell lymphoma morphology|9702/3
C0020981|T191|SY|0000006589|CHV|aild|9705/3
C0020981|T191|SY|0000006589|CHV|angioblastic lymphadenopathy|9705/3
C0020981|T191|PT|0000006589|CHV|angioimmunoblastic lymphadenopathy|9705/3
C0020981|T191|SY|0000006589|CHV|angioimmunoblastic lymphoma|9705/3
C0020981|T191|SY|0000006589|CHV|immunoblastic lymphadenopathy|9705/3
C0020981|T191|DI|U001112|DXP|LYMPHADENOPATHY, ANGIOIMMUNOBLASTIC, WITH DYSPROTEINEMIA|9705/3
C0020981|T191|SY|NOCODE|DXP|LYMPHADENOPATHY, IMMUNOBLASTIC|9705/3
C0020981|T191|PT|C86.5|ICD10CM|Angioimmunoblastic T-cell lymphoma|9705/3
C0020981|T191|AB|C86.5|ICD10CM|Angioimmunoblastic T-cell lymphoma|9705/3
C0020981|T191|PT|MTHU006365|ICPC2ICD10ENG|angioimmunoblastic; lymphadenopathy|9705/3
C0020981|T191|PT|MTHU006366|ICPC2ICD10ENG|angioimmunoblastic; lymphoma|9705/3
C0020981|T191|PT|MTHU046565|ICPC2ICD10ENG|lymphadenopathy; angioimmunoblastic|9705/3
C0020981|T191|PT|MTHU046737|ICPC2ICD10ENG|lymphoma; angioimmunoblastic|9705/3
C0020981|T191|LLT|10080248|MDR|Angioimmunoblastic lymphadenopathy|9705/3
C0020981|T191|LLT|10079289|MDR|Angioimmunoblastic lymphadenopathy with dysproteinaemia|9705/3
C0020981|T191|LLT|10079282|MDR|Angioimmunoblastic lymphadenopathy with dysproteinemia|9705/3
C0020981|T191|LLT|10002449|MDR|Angioimmunoblastic T-cell lymphoma|9705/3
C0020981|T191|PT|10002449|MDR|Angioimmunoblastic T-cell lymphoma|9705/3
C0020981|T191|LLT|10002451|MDR|Angioimmunoblastic T-cell lymphoma NOS|9705/3
C0020981|T191|HT|10002450|MDR|Angioimmunoblastic T-cell lymphomas|9705/3
C0020981|T191|SY|31466|MEDCIN|AILD|9705/3
C0020981|T191|PT|31466|MEDCIN|angioimmunoblastic T-cell lymphoma|9705/3
C0020981|T191|SY|33782|MEDCIN|immunoblastic lymphadenopathy|9705/3
C0020981|T191|PT|33782|MEDCIN|malignant immunoblastic lymphadenopathy|9705/3
C0020981|T191|PM|D007119|MSH|Angioimmunoblastic Lymphadenopathies|9705/3
C0020981|T191|ET|D007119|MSH|Angioimmunoblastic Lymphadenopathy|9705/3
C0020981|T191|PM|D007119|MSH|Immunoblastic Lymphadenopathies|9705/3
C0020981|T191|MH|D007119|MSH|Immunoblastic Lymphadenopathy|9705/3
C0020981|T191|PM|D007119|MSH|Lymphadenopathies, Angioimmunoblastic|9705/3
C0020981|T191|PM|D007119|MSH|Lymphadenopathies, Immunoblastic|9705/3
C0020981|T191|PM|D007119|MSH|Lymphadenopathy, Angioimmunoblastic|9705/3
C0020981|T191|ET|D007119|MSH|Lymphadenopathy, Immunoblastic|9705/3
C0020981|T191|PN|NOCODE|MTH|Angioimmunoblastic Lymphadenopathy|9705/3
C0020981|T191|AB|C7528|NCI|AILD|9705/3
C0020981|T191|AB|C7528|NCI|AILT|9705/3
C0020981|T191|OP|C7528|NCI|Angioimmunoblastic Lymphadenopathy|9705/3
C0020981|T191|SY|C7528|NCI|Angioimmunoblastic Lymphadenopathy Type T-Cell Lymphoma|9705/3
C0020981|T191|OP|C7528|NCI|Angioimmunoblastic Lymphadenopathy with Dysproteinemia|9705/3
C0020981|T191|PT|C7528|NCI|Angioimmunoblastic T-Cell Lymphoma|9705/3
C0020981|T191|SY|TCGA|NCI|Angioimmunoblastic T-Cell Lymphoma|9705/3
C0020981|T191|PT|C7528|NCI_CPTAC|Angioimmunoblastic T-Cell Lymphoma|9705/3
C0020981|T191|DN|C7528|NCI_CTRP|Angioimmunoblastic T-Cell Lymphoma|9705/3
C0020981|T191|PT|CDR0000346464|NCI_NCI-GLOSS|angioimmunoblastic T-cell lymphoma|9705/3
C0020981|T191|AB|CDR0000042765|PDQ|AILD|9705/3
C0020981|T191|AB|CDR0000042765|PDQ|AILT|9705/3
C0020981|T191|IS|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy|9705/3
C0020981|T191|SY|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy|9705/3
C0020981|T191|SY|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy type T-cell lymphoma|9705/3
C0020981|T191|IS|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy with dysproteinemia|9705/3
C0020981|T191|SY|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy with dysproteinemia|9705/3
C0020981|T191|PT|CDR0000042765|PDQ|angioimmunoblastic T-cell lymphoma|9705/3
C0020981|T191|PT|Q0300328|QMR|ANGIOIMMUNOBLASTIC LYMPHADENOPATHY|9705/3
C0020981|T191|AB|Xa0Tk|RCD|Angioim lymphadenopy+dysprot|9705/3
C0020981|T191|PT|Xa0Tk|RCD|Angioimmunoblastic lymphadenopathy with dysproteinaemia|9705/3
C0020981|T191|SY|Xa0Tk|RCD|Angioimmunoblastic lymphoma|9705/3
C0020981|T191|PT|Xa0Tk|RCDAE|Angioimmunoblastic lymphadenopathy with dysproteinemia|9705/3
C0020981|T191|OA|BBm8.|RCDSY|Angioimmunoblas lymphadenop|9705/3
C0020981|T191|OP|BBm8.|RCDSY|Angioimmunoblastic lymphadenopathy|9705/3
C0020981|T191|OAS|127216000|SNOMEDCT_US|AILD|9705/3
C0020981|T191|PT|52097008|SNOMEDCT_US|Angioimmunoblastic lymphadenopathy|9705/3
C0020981|T191|OAP|127216000|SNOMEDCT_US|Angioimmunoblastic lymphadenopathy with dysproteinaemia|9705/3
C0020981|T191|OAP|127216000|SNOMEDCT_US|Angioimmunoblastic lymphadenopathy with dysproteinemia|9705/3
C0020981|T191|SY|835009|SNOMEDCT_US|Angioimmunoblastic lymphoma|9705/3
C0020981|T191|PT|835009|SNOMEDCT_US|Angioimmunoblastic T-cell lymphoma|9705/3
C0020981|T191|PT|413537009|SNOMEDCT_US|Angioimmunoblastic T-cell lymphoma|9705/3
C0522624|T191|AB|C86.3|ICD10CM|Subcutaneous panniculitis-like T-cell lymphoma|9708/3
C0522624|T191|PT|C86.3|ICD10CM|Subcutaneous panniculitis-like T-cell lymphoma|9708/3
C0522624|T191|SY|338549|MEDCIN|lymphoma mature t-cell subcutaneous panniculitis-like|9708/3
C0522624|T191|PT|338549|MEDCIN|subcutaneous panniculitis-like T-cell lymphoma|9708/3
C0522624|T191|NM|C537503|MSH|Subcutaneous panniculitis-like T-cell lymphoma|9708/3
C0522624|T191|PN|NOCODE|MTH|Subcutaneous panniculitis-like T-cell lymphoma|9708/3
C0522624|T191|AB|C6918|NCI|SPTCL|9708/3
C0522624|T191|PT|C6918|NCI|Subcutaneous Panniculitis-Like T-Cell Lymphoma|9708/3
C0522624|T191|SY|TCGA|NCI|Subcutaneous Panniculitis-Like T-Cell Lymphoma|9708/3
C0522624|T191|SY|C6918|NCI|Subcutaneous Panniculitis-Like T-Cell Lymphoma, Alpha/Beta Type|9708/3
C0522624|T191|SY|404133000|SNOMEDCT_US|Subcutaneous panniculitic cutaneous T-cell lymphoma|9708/3
C0522624|T191|SY|103682005|SNOMEDCT_US|Subcutaneous panniculitic T-cell lymphoma|9708/3
C0522624|T191|PT|404133000|SNOMEDCT_US|Subcutaneous panniculitis-like T-cell lymphoma|9708/3
C0522624|T191|PT|103682005|SNOMEDCT_US|Subcutaneous panniculitis-like T-cell lymphoma|9708/3
C0079773|T191|SY|0000015230|CHV|cells cutaneous lymphomas t|9709/3
C0079773|T191|SY|0000015230|CHV|cutaneous t cell lymphoma|9709/3
C0079773|T191|PT|0000015230|CHV|cutaneous t-cell lymphoma|9709/3
C0079773|T191|SY|0000015230|CHV|t cell cutaneous lymphoma|9709/3
C0079773|T191|ET|2004-7126|CSP|cutaneous T cell lymphoma|9709/3
C0079773|T191|PT|HP:0012192|HPO|Cutaneous T-cell lymphoma|9709/3
C0079773|T191|PT|10011677|MDR|Cutaneous T-cell lymphoma|9709/3
C0079773|T191|LLT|10011677|MDR|Cutaneous T-cell lymphoma|9709/3
C0079773|T191|PT|351484|MEDCIN|Primary cutaneous T-cell lymphoma|9709/3
C0079773|T191|SY|351484|MEDCIN|skin malignant lymphoma mature t-cell cutaneous primary|9709/3
C0079773|T191|PM|D016410|MSH|Cutaneous T Cell Lymphoma|9709/3
C0079773|T191|ET|D016410|MSH|Cutaneous T-Cell Lymphoma|9709/3
C0079773|T191|PM|D016410|MSH|Cutaneous T-Cell Lymphomas|9709/3
C0079773|T191|PM|D016410|MSH|Lymphoma, Cutaneous T-Cell|9709/3
C0079773|T191|ET|D016410|MSH|Lymphoma, T Cell, Cutaneous|9709/3
C0079773|T191|MH|D016410|MSH|Lymphoma, T-Cell, Cutaneous|9709/3
C0079773|T191|PM|D016410|MSH|Lymphomas, Cutaneous T-Cell|9709/3
C0079773|T191|PM|D016410|MSH|T Cell Lymphoma, Cutaneous|9709/3
C0079773|T191|ET|D016410|MSH|T-Cell Lymphoma, Cutaneous|9709/3
C0079773|T191|PM|D016410|MSH|T-Cell Lymphomas, Cutaneous|9709/3
C0079773|T191|PN|NOCODE|MTH|Lymphoma, T-Cell, Cutaneous|9709/3
C0079773|T191|AB|C3467|NCI|CTCL|9709/3
C0079773|T191|SY|C3467|NCI|Cutaneous T Cell Lymphoma|9709/3
C0079773|T191|SY|C3467|NCI|Cutaneous T-Cell Non-Hodgkin Lymphoma|9709/3
C0079773|T191|SY|C3467|NCI|Cutaneous T-Cell Non-Hodgkin's Lymphoma|9709/3
C0079773|T191|AB|C3467|NCI|PCTCL|9709/3
C4528220|T191|PT|C139023|NCI|Primary Cutaneous Acral CD8-Positive T-Cell Lymphoma|9709/3
C4518232|T191|SY|C45339|NCI|Primary Cutaneous Aggressive Epidermotropic CD8-Positive T-Cell Lymphoma|9709/3
C4528627|T191|PT|C45366|NCI|Primary Cutaneous CD4-Positive Small/Medium T-Cell Lymphoproliferative Disorder|9709/3
C4528627|T191|SY|C45366|NCI|Primary Cutaneous CD4-Positive Small/Medium-Sized Pleomorphic T-Cell Lymphoproliferative Disorder|9709/3
C4528627|T191|SY|C45366|NCI|Primary Cutaneous CD4-Positive Small/Medium-Sized T-Cell Lymphoproliferative Disorder|9709/3
C4518232|T191|PT|C45339|NCI|Primary Cutaneous CD8-Positive Aggressive Epidermotropic Cytotoxic T-Cell Lymphoma|9709/3
C4518232|T191|SY|C45339|NCI|Primary Cutaneous CD8-Positive Aggressive Epidermotropic T-Cell Lymphoma|9709/3
C0079773|T191|PT|C3467|NCI|Primary Cutaneous T-Cell Non-Hodgkin Lymphoma|9709/3
C0079773|T191|SY|C3467|NCI|Primary Cutaneous T-Cell Non-Hodgkin's Lymphoma|9709/3
C0079773|T191|SY|C3467|NCI|Skin T-Cell Non-Hodgkin's Lymphoma|9709/3
C0079773|T191|SY|C3467|NCI|T-Cell Non-Hodgkin's Lymphoma of Skin|9709/3
C0079773|T191|SY|C3467|NCI|T-Cell Non-Hodgkin's Lymphoma of the Skin|9709/3
C0079773|T191|PT|C3467|NCI_CPTAC|Primary Cutaneous T-Cell Non-Hodgkin Lymphoma|9709/3
C0079773|T191|DN|C3467|NCI_CTRP|Cutaneous T-Cell Non-Hodgkin Lymphoma|9709/3
C0079773|T191|PT|CDR0000046771|NCI_NCI-GLOSS|cutaneous T-cell lymphoma|9709/3
C0079773|T191|AB|CDR0000043725|PDQ|CTCL|9709/3
C0079773|T191|SY|CDR0000043725|PDQ|cutaneous T-cell lymphoma|9709/3
C0079773|T191|PSC|CDR0000043725|PDQ|cutaneous T-cell non-Hodgkin lymphoma|9709/3
C0079773|T191|SY|CDR0000043725|PDQ|lymphoma, cutaneous T-cell|9709/3
C0079773|T191|SY|CDR0000043725|PDQ|T cell lymphoma, cutaneous|9709/3
C0079773|T191|SY|CDR0000043725|PDQ|T-cell lymphoma, cutaneous|9709/3
C0079773|T191|PT|R0121577|QMR|CUTANEOUS T-CELL LYMPHOMA|9709/3
C0079773|T191|AB|X78hl|RCD|CTCL - Cutan T-cell lymphoma|9709/3
C0079773|T191|SY|X78hl|RCD|CTCL - Cutaneous T-cell lymphoma|9709/3
C0079773|T191|SY|X78hl|RCD|Cutaneous T-cell lymphoma|9709/3
C4518232|T191|SY|765136002|SNOMEDCT_US|Berti lymphoma|9709/3
C0079773|T191|OAS|255099004|SNOMEDCT_US|CTCL - Cutaneous T-cell lymphoma|9709/3
C0079773|T191|SY|400122007|SNOMEDCT_US|CTCL - Cutaneous T-cell lymphoma|9709/3
C0079773|T191|PT|28054005|SNOMEDCT_US|Cutaneous T-cell lymphoma|9709/3
C0079773|T191|OAS|255099004|SNOMEDCT_US|Cutaneous T-cell lymphoma|9709/3
C0079773|T191|SY|400122007|SNOMEDCT_US|Cutaneous T-cell lymphoma|9709/3
C0079773|T191|SY|28054005|SNOMEDCT_US|Cutaneous T-cell lymphoma, no ICD-O subtype|9709/3
C0079773|T191|SY|28054005|SNOMEDCT_US|Cutaneous T-cell lymphoma, no International Classification of Diseases for Oncology subtype|9709/3
C1690583|T191|OAS|419563005|SNOMEDCT_US|Cutaneous T-cell lymphoma, pleomorphic small/medium-sized|9709/3
C4528627|T191|SY|788674000|SNOMEDCT_US|PCSM-TCL- primary cutaneous CD4 positive small/medium T-cell lymphoproliferative disorder|9709/3
C4528220|T191|PT|787198005|SNOMEDCT_US|Primary cutaneous acral CD8 positive T-cell lymphoma|9709/3
C4528627|T191|PT|788674000|SNOMEDCT_US|Primary cutaneous CD4 positive small/medium T-cell lymphoproliferative disorder|9709/3
C4528627|T191|PT|788570002|SNOMEDCT_US|Primary cutaneous CD4-positive small/medium T-cell lymphoproliferative disorder|9709/3
C4518232|T191|PT|765136002|SNOMEDCT_US|Primary cutaneous CD8 positive aggressive epidermotropic cytotoxic T-cell lymphoma|9709/3
C4518232|T191|PT|733895005|SNOMEDCT_US|Primary cutaneous CD8 positive aggressive epidermotropic cytotoxic T-cell lymphoma|9709/3
C4518232|T191|SY|765136002|SNOMEDCT_US|Primary cutaneous epidermotropic cytotoxic CD8 positive T-cell lymphoma|9709/3
C1640806|T191|PT|419018000|SNOMEDCT_US|Primary cutaneous large T-cell lymphoma - category|9709/3
C0079773|T191|PT|400122007|SNOMEDCT_US|Primary cutaneous T-cell lymphoma|9709/3
C1634515|T191|PT|419283005|SNOMEDCT_US|Primary cutaneous T-cell lymphoma - category|9709/3
C1690583|T191|OAP|419563005|SNOMEDCT_US|Primary cutaneous T-cell lymphoma, pleomorphic small/medium-sized|9709/3
C0334660|T191|SY|0000030017|CHV|angioendotheliomatosis|9712/3
C0334660|T191|PT|0000030017|CHV|intravascular lymphomatosis|9712/3
C0334660|T191|ET|C83.8|ICD10CM|Intravascular large B-cell lymphoma|9712/3
C0334660|T191|PT|MTHU006358|ICPC2ICD10ENG|angioendotheliomatosis|9712/3
C0334660|T191|LLT|10069643|MDR|Intravascular large B-cell lymphoma|9712/3
C0334660|T191|PT|355310|MEDCIN|Angioendotheliomatosis|9712/3
C0334660|T191|SY|355310|MEDCIN|malignant neoplasm lymphoma b-cell high grade diffuse angioendotheliomatosis|9712/3
C0334660|T191|PN|NOCODE|MTH|Angioendotheliomatosis|9712/3
C0334660|T191|SY|C4342|NCI|Angiotropic Large Cell Lymphoma|9712/3
C0334660|T191|SY|C4342|NCI|Angiotropic Lymphoma|9712/3
C0334660|T191|SY|C4342|NCI|Intravascular B-Cell Lymphoma|9712/3
C0334660|T191|PT|C4342|NCI|Intravascular Large B-Cell Lymphoma|9712/3
C0334660|T191|SY|C4342|NCI|Malignant Angioendotheliomatosis|9712/3
C0334660|T191|PT|X78hp|RCD|Angioendotheliomatosis|9712/3
C0334660|T191|SY|X78hp|RCD|Intravascular lymphomatosis|9712/3
C0334660|T191|AB|X78hp|RCD|Malignant angioendotheliomatos|9712/3
C0334660|T191|SY|X78hp|RCD|Malignant angioendotheliomatosis|9712/3
C0334660|T191|OP|BBv1.|RCDSY|Angioendotheliomatosis|9712/3
C0334660|T191|OP|BBmJ.|RCDSY|Angioendotheliomatosis|9712/3
C0334660|T191|PT|255102004|SNOMEDCT_US|Angioendotheliomatosis|9712/3
C0334660|T191|OAP|17158006|SNOMEDCT_US|Angioendotheliomatosis|9712/3
C0334660|T191|SY|46732000|SNOMEDCT_US|Angioendotheliomatosis|9712/3
C0334660|T191|IS|17158006|SNOMEDCT_US|Angioendotheliomatosis -RETIRED-|9712/3
C0334660|T191|OF|17158006|SNOMEDCT_US|Angioendotheliomatosis -RETIRED-|9712/3
C0334660|T191|SY|46732000|SNOMEDCT_US|Angiotropic lymphoma|9712/3
C0334660|T191|SY|46732000|SNOMEDCT_US|Intravascular B-cell lymphoma|9712/3
C0334660|T191|PT|399648005|SNOMEDCT_US|Intravascular large B-cell lymphoma|9712/3
C0334660|T191|SY|46732000|SNOMEDCT_US|Intravascular large B-cell lymphoma|9712/3
C0334660|T191|SY|255102004|SNOMEDCT_US|Intravascular lymphomatosis|9712/3
C0334660|T191|SY|255102004|SNOMEDCT_US|Malignant angioendotheliomatosis|9712/3
C0206180|T191|PT|0000020845|CHV|anaplastic large cell lymphoma|9714/3
C0206180|T191|SY|0000020845|CHV|ki 1 lymphoma|9714/3
C0206180|T191|SY|0000020845|CHV|ki-1 lymphoma|9714/3
C0206180|T191|SY|0000020845|CHV|large cell anaplastic lymphoma|9714/3
C0206180|T191|PT|HP:0012193|HPO|Anaplastic large-cell lymphoma|9714/3
C1332079|T191|HT|C84.6|ICD10CM|Anaplastic large cell lymphoma, ALK-positive|9714/3
C1332079|T191|AB|C84.6|ICD10CM|Anaplastic large cell lymphoma, ALK-positive|9714/3
C0206180|T191|ET|C84.6|ICD10CM|Anaplastic large cell lymphoma, CD30-positive|9714/3
C0206180|T191|HT|200.6|ICD9CM|Anaplastic large cell lymphoma|9714/3
C0206180|T191|LLT|10073478|MDR|Anaplastic large-cell lymphoma|9714/3
C0206180|T191|PT|10073478|MDR|Anaplastic large-cell lymphoma|9714/3
C1332079|T191|PT|333216|MEDCIN|alk-positive anaplastic large cell lymphoma|9714/3
C0206180|T191|PT|312891|MEDCIN|anaplastic large cell lymphoma|9714/3
C1332079|T191|SY|333216|MEDCIN|lymphoma anaplastic large cell alk-positive|9714/3
C0206180|T191|PM|D017728|MSH|Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|ET|D017728|MSH|Anaplastic Large-Cell Lymphoma|9714/3
C0206180|T191|PM|D017728|MSH|Anaplastic Large-Cell Lymphomas|9714/3
C0206180|T191|DSV|D017728|MSH|CD 030 POSITIVE ANAPLASTIC LARGE CELL LYMPHOMA|9714/3
C0206180|T191|PM|D017728|MSH|CD30 Positive Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|ET|D017728|MSH|CD30-Positive Anaplastic Large-Cell Lymphoma|9714/3
C0206180|T191|PM|D017728|MSH|CD30+ Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|ET|D017728|MSH|CD30+ Anaplastic Large-Cell Lymphoma|9714/3
C0206180|T191|PM|D017728|MSH|Ki 1 Lymphoma|9714/3
C0206180|T191|ET|D017728|MSH|Ki-1 Lymphoma|9714/3
C0206180|T191|PM|D017728|MSH|Ki-1 Lymphomas|9714/3
C0206180|T191|PM|D017728|MSH|Large-Cell Lymphoma, Anaplastic|9714/3
C0206180|T191|PM|D017728|MSH|Large-Cell Lymphomas, Anaplastic|9714/3
C0206180|T191|DSV|D017728|MSH|LYMPHOMA LARGE CELL KI 01|9714/3
C0206180|T191|PM|D017728|MSH|Lymphoma, Anaplastic Large-Cell|9714/3
C0206180|T191|PM|D017728|MSH|Lymphoma, Ki-1|9714/3
C0206180|T191|MH|D017728|MSH|Lymphoma, Large-Cell, Anaplastic|9714/3
C0206180|T191|ET|D017728|MSH|Lymphoma, Large-Cell, Ki-1|9714/3
C0206180|T191|PM|D017728|MSH|Lymphomas, Anaplastic Large-Cell|9714/3
C0206180|T191|PM|D017728|MSH|Lymphomas, Ki-1|9714/3
C0206180|T191|PM|D017728|MSH|Systemic Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|ET|D017728|MSH|Systemic Anaplastic Large-Cell Lymphoma|9714/3
C0206180|T191|PN|NOCODE|MTH|Ki-1+ Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|AB|C3720|NCI|ALCL|9714/3
C1332079|T191|AB|C37193|NCI|ALCL, ALK+|9714/3
C1332079|T191|SY|C37193|NCI|ALK-Positive Anaplastic Large Cell Lymphoma|9714/3
C1332079|T191|SY|C37193|NCI|ALKoma|9714/3
C0206180|T191|SY|TCGA|NCI|Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|PT|C3720|NCI|Anaplastic Large Cell Lymphoma|9714/3
C1332079|T191|PT|C37193|NCI|Anaplastic Large Cell Lymphoma, ALK-Positive|9714/3
C0206180|T191|SY|C3720|NCI|CD30 Positive Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|OP|C3720|NCI|Ki-1 Lymphoma|9714/3
C0206180|T191|OP|C3720|NCI|Ki-1+ ALCL|9714/3
C0206180|T191|OP|C3720|NCI|Ki-1+ Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|PT|C3720|NCI_CPTAC|Anaplastic Large Cell Lymphoma|9714/3
C1332079|T191|PT|C37193|NCI_CPTAC|Anaplastic Large Cell Lymphoma, ALK-Positive|9714/3
C0206180|T191|DN|C3720|NCI_CTRP|Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|SY|3264|NCI_FDA|ALCL|9714/3
C0206180|T191|PT|3264|NCI_FDA|Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|PT|CDR0000575433|NCI_NCI-GLOSS|ALCL|9714/3
C0206180|T191|PT|CDR0000045552|NCI_NCI-GLOSS|anaplastic large cell lymphoma|9714/3
C0206180|T191|AB|CDR0000042785|PDQ|ALCL|9714/3
C0206180|T191|PT|CDR0000042785|PDQ|anaplastic large cell lymphoma|9714/3
C0206180|T191|SY|CDR0000042785|PDQ|CD30 Positive Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|IS|CDR0000042785|PDQ|Ki-1 Lymphoma|9714/3
C0206180|T191|SY|CDR0000042785|PDQ|Ki-1+ ALCL|9714/3
C0206180|T191|SY|CDR0000042785|PDQ|Ki-1+ Anaplastic Large Cell Lymphoma|9714/3
C0206180|T191|SY|CDR0000042785|PDQ|lymphoma, anaplastic large cell|9714/3
C0206180|T191|PT|Xa0TS|RCD|Large cell anaplastic lymphoma|9714/3
C0206180|T191|SY|53237008|SNOMEDCT_US|Anaplastic large cell lymphoma|9714/3
C0206180|T191|SY|53237008|SNOMEDCT_US|Anaplastic large cell lymphoma, CD30+|9714/3
C0206180|T191|PT|53237008|SNOMEDCT_US|Anaplastic large cell lymphoma, T cell and Null cell type|9714/3
C1531540|T191|SY|413527004|SNOMEDCT_US|Anaplastic large cell lymphoma, T- and null cell primary systemic types|9714/3
C1531540|T191|PT|703626001|SNOMEDCT_US|Anaplastic large cell lymphoma, T/Null cell, primary systemic type|9714/3
C1531540|T191|PT|413527004|SNOMEDCT_US|Anaplastic large cell lymphoma, T/Null cell, primary systemic type|9714/3
C4518436|T191|PT|738770003|SNOMEDCT_US|Anaplastic lymphoma kinase positive anaplastic large cell lymphoma|9714/3
C4518436|T191|PT|734044003|SNOMEDCT_US|Anaplastic lymphoma kinase positive anaplastic large cell lymphoma|9714/3
C0206180|T191|PT|277637000|SNOMEDCT_US|Large cell anaplastic lymphoma|9714/3
C1333984|T191|AB|C86.1|ICD10CM|Hepatosplenic T-cell lymphoma|9716/3
C1333984|T191|PT|C86.1|ICD10CM|Hepatosplenic T-cell lymphoma|9716/3
C1333984|T191|LLT|10076434|MDR|Hepatosplenic gamma-delta T-cell lymphoma|9716/3
C1333984|T191|LLT|10066957|MDR|Hepatosplenic T-cell lymphoma|9716/3
C1333984|T191|PT|10066957|MDR|Hepatosplenic T-cell lymphoma|9716/3
C0522627|T191|PT|368855|MEDCIN|Hepatosplenic gamma-delta cell lymphoma|9716/3
C1333984|T191|PT|338550|MEDCIN|hepatosplenic T-cell lymphoma|9716/3
C1333984|T191|SY|338550|MEDCIN|malignant neoplasm lymphoma mature t-cell hepatosplenic|9716/3
C0522627|T191|SY|368855|MEDCIN|non-hodgkin's lymphoma hepatosplenic gamma-delta cell|9716/3
C1333984|T191|SY|C8459|NCI|Hepatosplenic Gamma/Delta T-Cell Lymphoma|9716/3
C1333984|T191|PT|C8459|NCI|Hepatosplenic T-Cell Lymphoma|9716/3
C1333984|T191|SY|TCGA|NCI|Hepatosplenic T-Cell Lymphoma|9716/3
C1333984|T191|DN|C8459|NCI_CTRP|Hepatosplenic T-Cell Lymphoma|9716/3
C1333984|T191|SY|CDR0000613812|PDQ|Hepatosplenic Gamma/Delta T-Cell Lymphoma|9716/3
C1333984|T191|PT|CDR0000613812|PDQ|hepatosplenic T-cell lymphoma|9716/3
C0522627|T191|PT|103685007|SNOMEDCT_US|Hepatosplenic gamma-delta cell lymphoma|9716/3
C0522627|T191|PT|699657009|SNOMEDCT_US|Hepatosplenic gamma-delta cell lymphoma|9716/3
C1333984|T191|PT|445406001|SNOMEDCT_US|Hepatosplenic T-cell lymphoma|9716/3
C0456889|T191|ET|C86.2|ICD10CM|Enteropathy associated T-cell lymphoma|9717/3
C0456889|T191|PT|10073481|MDR|Enteropathy-associated T-cell lymphoma|9717/3
C0456889|T191|LLT|10073481|MDR|Enteropathy-associated T-cell lymphoma|9717/3
C4721452|T191|LLT|10022703|MDR|Intestinal T-cell lymphoma|9717/3
C4721452|T191|LLT|10022705|MDR|Intestinal T-cell lymphoma NOS|9717/3
C4721452|T191|HT|10022704|MDR|Intestinal T-cell lymphomas|9717/3
C0456889|T191|SY|271162|MEDCIN|digestive malignant lymphoma intestinal T-cell|9717/3
C0456889|T191|PT|352247|MEDCIN|Enteropathy associated T-cell lymphoma|9717/3
C4721452|T191|PT|271162|MEDCIN|intestinal T-cell lymphoma|9717/3
C0456889|T191|SY|352247|MEDCIN|lymphoma mature t-cell enteropathy associated|9717/3
C0456889|T191|PM|D058527|MSH|Enteropathy Associated T Cell Lymphoma|9717/3
C0456889|T191|MH|D058527|MSH|Enteropathy-Associated T-Cell Lymphoma|9717/3
C0456889|T191|PM|D058527|MSH|Enteropathy-Associated T-Cell Lymphomas|9717/3
C0456889|T191|ET|D058527|MSH|Lymphoma, T-Cell, Enteropathy-Associated|9717/3
C0456889|T191|PM|D058527|MSH|Lymphomas, Enteropathy-Associated T-Cell|9717/3
C0456889|T191|PM|D058527|MSH|T Cell Lymphoma, Enteropathy Associated|9717/3
C0456889|T191|ET|D058527|MSH|T-Cell Lymphoma, Enteropathy-Associated|9717/3
C0456889|T191|PM|D058527|MSH|T-Cell Lymphomas, Enteropathy-Associated|9717/3
C0456889|T191|PN|NOCODE|MTH|Enteropathy-Associated T-Cell Lymphoma|9717/3
C4721452|T191|PN|NOCODE|MTH|Intestinal T-Cell Lymphoma|9717/3
C0456889|T191|SY|C4737|NCI|EATL, Type I|9717/3
C0456889|T191|SY|C4737|NCI|Enteropathy Associated T-Cell Lymphoma|9717/3
C0456889|T191|PT|C4737|NCI|Enteropathy-Associated T-Cell Lymphoma|9717/3
C0456889|T191|SY|TCGA|NCI|Enteropathy-Associated T-Cell Lymphoma|9717/3
C0456889|T191|SY|C4737|NCI|Enteropathy-Associated T-Cell Lymphoma, Type I|9717/3
C0456889|T191|SY|C4737|NCI|Enteropathy-Type T-Cell Lymphoma|9717/3
C4721452|T191|PT|C150495|NCI|Intestinal T-Cell Lymphoma|9717/3
C3272525|T191|AB|C96058|NCI|MEITL|9717/3
C3272525|T191|SY|C96058|NCI|Monomorphic CD56+ Intestinal T-Cell Lymphoma|9717/3
C3272525|T191|PT|C96058|NCI|Monomorphic Epitheliotropic Intestinal T-Cell Lymphoma|9717/3
C3272525|T191|SY|C96058|NCI|Type II EATL|9717/3
C0456889|T191|DN|C4737|NCI_CTRP|Enteropathy-Associated T-Cell Lymphoma|9717/3
C4721452|T191|DN|C150495|NCI_CTRP|Intestinal T-Cell Lymphoma|9717/3
C0456889|T191|AB|Xa0Tu|RCD|EACTL - Ent-ass T-cell lymphom|9717/3
C0456889|T191|SY|Xa0Tu|RCD|EACTL - Enteropathy-associated T-cell lymphoma|9717/3
C0456889|T191|AB|Xa0Tu|RCD|Enterop-assoc T-cell lymphoma|9717/3
C0456889|T191|PT|Xa0Tu|RCD|Enteropathy-associated T-cell lymphoma|9717/3
C0456889|T191|SY|277654008|SNOMEDCT_US|EACTL - Enteropathy-associated T-cell lymphoma|9717/3
C4721452|T191|SY|103686008|SNOMEDCT_US|Enteropathy associated T-cell lymphoma|9717/3
C0456889|T191|PT|277654008|SNOMEDCT_US|Enteropathy-associated T-cell lymphoma|9717/3
C0456889|T191|SY|277654008|SNOMEDCT_US|Enteropathy-type T-cell lymphoma|9717/3
C4721452|T191|SY|103686008|SNOMEDCT_US|Enteropathy-type T-cell lymphoma|9717/3
C4721452|T191|PT|103686008|SNOMEDCT_US|Intestinal T-cell lymphoma|9717/3
C3272525|T191|PT|787036009|SNOMEDCT_US|Monomorphic epitheliotropic intestinal T-cell lymphoma|9717/3
C0206182|T191|PT|0000020847|CHV|lymphomatoid papulosis|9718/1
C0206182|T191|PT|L41.2|ICD10|Lymphomatoid papulosis|9718/1
C0206182|T191|ET|C86.6|ICD10CM|Lymphomatoid papulosis|9718/1
C0206182|T191|PT|MTHU057362|ICPC2ICD10ENG|papulosis; lymphomatoid|9718/1
C0206182|T191|PT|10056670|MDR|Lymphomatoid papulosis|9718/1
C0206182|T191|LLT|10056670|MDR|Lymphomatoid papulosis|9718/1
C0206182|T191|PT|314716|MEDCIN|Lymphomatoid papulosis|9718/1
C0206182|T191|PM|D017731|MSH|Lymphomatoid Papuloses|9718/1
C0206182|T191|MH|D017731|MSH|Lymphomatoid Papulosis|9718/1
C0206182|T191|PM|D017731|MSH|Papuloses, Lymphomatoid|9718/1
C0206182|T191|PM|D017731|MSH|Papulosis, Lymphomatoid|9718/1
C0206182|T191|PN|NOCODE|MTH|Lymphomatoid Papulosis|9718/1
C0206182|T191|PT|C3721|NCI|Lymphomatoid Papulosis|9718/1
C0206182|T191|SY|TCGA|NCI|Lymphomatoid Papulosis|9718/1
C0206182|T191|AB|C3721|NCI|LyP|9718/1
C0206182|T191|PT|X50BR|RCD|Lymphomatoid papulosis|9718/1
C0206182|T191|OAP|200986009|SNOMEDCT_US|Lymphomatoid papulosis|9718/1
C0206182|T191|PT|397353001|SNOMEDCT_US|Lymphomatoid papulosis|9718/1
C0206182|T191|OF|200986009|SNOMEDCT_US|Lymphomatoid papulosis|9718/1
C0206182|T191|PT|31047003|SNOMEDCT_US|Lymphomatoid papulosis|9718/1
C0206182|T191|IS|128804002|SNOMEDCT_US|Lymphomatoid papulosis|9718/1
C1301362|T191|ET|C86.6|ICD10CM|Primary cutaneous anaplastic large cell lymphoma|9718/3
C1301362|T191|ET|C86.6|ICD10CM|Primary cutaneous CD30-positive large T-cell lymphoma|9718/3
C1301362|T191|LLT|10065863|MDR|Anaplastic large-cell lymphoma, primary cutaneous type|9718/3
C1301362|T191|MH|D054446|MSH|Lymphoma, Primary Cutaneous Anaplastic Large Cell|9718/3
C1301362|T191|ET|D054446|MSH|Primary Cutaneous Anaplastic Large Cell Lymphoma|9718/3
C1301362|T191|PM|D054446|MSH|Primary Cutaneous CD30 positive Large T Cell Lymphoma|9718/3
C1301362|T191|ET|D054446|MSH|Primary Cutaneous CD30-positive Large T-Cell Lymphoma|9718/3
C1301362|T191|PN|NOCODE|MTH|Primary Cutaneous Anaplastic Large Cell Lymphoma|9718/3
C1301362|T191|AB|C6860|NCI|C-ALCL|9718/3
C1301362|T191|SY|C6860|NCI|Primary Anaplastic Large Cell Lymphoma of Skin|9718/3
C1301362|T191|SY|C6860|NCI|Primary Anaplastic Large Cell Lymphoma of the Skin|9718/3
C1301362|T191|PT|C6860|NCI|Primary Cutaneous Anaplastic Large Cell Lymphoma|9718/3
C1301362|T191|SY|TCGA|NCI|Primary Cutaneous Anaplastic Large Cell Lymphoma|9718/3
C1301362|T191|SY|C6860|NCI|Primary Cutaneous CD30 Positive Anaplastic Large Cell Lymphoma|9718/3
C1371159|T191|PT|C7195|NCI|Primary Cutaneous CD30-Positive T-Cell Lymphoproliferative Disorder|9718/3
C1301362|T191|AB|C6860|NCI|Primary Cutaneous CD30+ ALCL|9718/3
C1301362|T191|SY|C6860|NCI|Primary Cutaneous CD30+ Anaplastic Large Cell Lymphoma|9718/3
C1371159|T191|SY|C7195|NCI|Primary Cutaneous CD30+ T-Cell Lymphoproliferative Disorder|9718/3
C1301362|T191|SY|10065863|NCI_CTEP-SDC|ALCL, cutaneous|9718/3
C1301362|T191|PT|10065863|NCI_CTEP-SDC|Anaplastic large-cell lymphoma, primary cutaneous type|9718/3
C1301362|T191|SY|397352006|SNOMEDCT_US|Anaplastic large cell lymphoma, T/Null cell, primary cutaneous type|9718/3
C1301362|T191|OAP|413526008|SNOMEDCT_US|Anaplastic large cell lymphoma, T/Null cell, primary cutaneous type|9718/3
C1301362|T191|SY|397352006|SNOMEDCT_US|Cutaneous T-cell lymphoma, large cell, CD30-positive|9718/3
C1301362|T191|SY|773995001|SNOMEDCT_US|pcALCL - primary cutaneous anaplastic large cell lymphoma|9718/3
C1301362|T191|IS|128804002|SNOMEDCT_US|Primary cutaneous anaplastic large cell lymphoma|9718/3
C1301362|T191|PT|773995001|SNOMEDCT_US|Primary cutaneous anaplastic large cell lymphoma|9718/3
C1301362|T191|PT|397352006|SNOMEDCT_US|Primary cutaneous anaplastic large cell lymphoma|9718/3
C1301362|T191|SY|397352006|SNOMEDCT_US|Primary cutaneous anaplastic large T-cell lymphoma, CD30-positive|9718/3
C1301362|T191|SY|128875000|SNOMEDCT_US|Primary cutaneous CD30 antigen positive large T-cell lymphoma|9718/3
C1371159|T191|SY|128804002|SNOMEDCT_US|Primary cutaneous CD30 antigen positive T-cell lymphoproliferative disorder|9718/3
C1301362|T191|PT|128875000|SNOMEDCT_US|Primary cutaneous CD30+ large T-cell lymphoma|9718/3
C1301362|T191|SY|128804002|SNOMEDCT_US|Primary cutaneous CD30+ large T-cell lymphoma|9718/3
C1371159|T191|PT|128804002|SNOMEDCT_US|Primary cutaneous CD30+ T-cell lymphoproliferative disorder|9718/3
C0392788|T191|PT|C86.0|ICD10CM|Extranodal NK/T-cell lymphoma, nasal type|9719/3
C0392788|T191|AB|C86.0|ICD10CM|Extranodal NK/T-cell lymphoma, nasal type|9719/3
C0558916|T191|ET|C84.9|ICD10CM|NK/T cell lymphoma NOS|9719/3
C0392788|T191|PT|MTHU006355|ICPC2ICD10ENG|angiocentric T-cell; lymphoma|9719/3
C0392788|T191|PT|MTHU046736|ICPC2ICD10ENG|lymphoma; angiocentric T-cell|9719/3
C0392788|T191|PT|MTHU046858|ICPC2ICD10ENG|lymphoma; T-cell, angiocentric|9719/3
C0392788|T191|PT|MTHU073541|ICPC2ICD10ENG|T-cell; lymphoma, angiocentric|9719/3
C0392788|T191|LLT|10002411|MDR|Angiocentric lymphoma|9719/3
C0392788|T191|PT|10002411|MDR|Angiocentric lymphoma|9719/3
C0392788|T191|LLT|10002413|MDR|Angiocentric lymphoma NOS|9719/3
C0392788|T191|HT|10002412|MDR|Angiocentric lymphomas|9719/3
C0392788|T191|LLT|10065855|MDR|Extranodal NK/T-cell lymphoma, nasal type|9719/3
C0392788|T191|PT|338145|MEDCIN|extranodal NK/T-cell lymphoma of nasal cavity|9719/3
C0392788|T191|PM|D054391|MSH|Extranodal NK T Cell Lymphoma, Nasal|9719/3
C0392788|T191|PM|D054391|MSH|Extranodal NK T Cell Lymphoma, Nasal and Nasal Type|9719/3
C0392788|T191|PM|D054391|MSH|Extranodal NK T Cell Lymphoma, Nasal Type|9719/3
C0392788|T191|ET|D054391|MSH|Extranodal NK-T-Cell Lymphoma, Nasal|9719/3
C0392788|T191|PEP|D054391|MSH|Extranodal NK-T-Cell Lymphoma, Nasal and Nasal-Type|9719/3
C0392788|T191|ET|D054391|MSH|Extranodal NK-T-Cell Lymphoma, Nasal Type|9719/3
C0558916|T191|PN|NOCODE|MTH|Nasal and nasal-type NK/T-cell lymphoma|9719/3
C0392788|T191|PN|NOCODE|MTH|Nasal Type Extranodal NK/T-Cell Lymphoma|9719/3
C0392788|T191|SY|C4684|NCI|Angiocentric T-Cell Lymphoma|9719/3
C0392788|T191|SY|C4684|NCI|Extranodal NK/T-Cell Lymphoma, Nasal Type|9719/3
C0392788|T191|PT|C4684|NCI|Nasal Type Extranodal NK/T-Cell Lymphoma|9719/3
C0392788|T191|SY|TCGA|NCI|Nasal Type Extranodal NK/T-Cell Lymphoma|9719/3
C0392788|T191|SY|C4684|NCI_CDISC|Angiocentric T-Cell Lymphoma|9719/3
C0392788|T191|PT|C4684|NCI_CDISC|RETICULOSIS, MALIGNANT|9719/3
C0392788|T191|SY|10065855|NCI_CTEP-SDC|Extranodal NK/T lymphoma-nasal|9719/3
C0392788|T191|PT|10065855|NCI_CTEP-SDC|Extranodal NK/T-cell lymphoma, nasal type|9719/3
C0392788|T191|DN|C4684|NCI_CTRP|Nasal Type Extranodal NK/T-Cell Lymphoma|9719/3
C0392788|T191|SY|CDR0000489005|PDQ|angiocentric T-cell lymphoma|9719/3
C0392788|T191|SY|CDR0000489005|PDQ|Nasal Type Extranodal NK/T-Cell Lymphoma|9719/3
C0392788|T191|PT|Xa0To|RCD|Angiocentric T-cell lymphoma|9719/3
C0558916|T191|OP|BBv2.|RCDSY|AngiocentricT-cell lymphoma|9719/3
C0392788|T191|OF|188689002|SNOMEDCT_US|Angiocentric T-cell lymphoma|9719/3
C0392788|T191|SY|414166008|SNOMEDCT_US|Angiocentric T-cell lymphoma|9719/3
C0392788|T191|OAP|66855003|SNOMEDCT_US|Angiocentric T-cell lymphoma|9719/3
C0392788|T191|OAP|188689002|SNOMEDCT_US|Angiocentric T-cell lymphoma|9719/3
C0392788|T191|OAP|277648007|SNOMEDCT_US|Angiocentric T-cell lymphoma|9719/3
C0392788|T191|IS|66855003|SNOMEDCT_US|Angiocentric T-cell lymphoma -RETIRED-|9719/3
C0392788|T191|OF|66855003|SNOMEDCT_US|Angiocentric T-cell lymphoma -RETIRED-|9719/3
C0392788|T191|SY|414166008|SNOMEDCT_US|Extranodal natural killer/T-cell lymphoma, nasal type|9719/3
C0392788|T191|PT|414166008|SNOMEDCT_US|Extranodal NK/T-cell lymphoma, nasal type|9719/3
C0558916|T191|SY|128805001|SNOMEDCT_US|Natural killer-/T-cell lymphoma, nasal and nasal-type|9719/3
C0558916|T191|PT|128805001|SNOMEDCT_US|NK/T-cell lymphoma, nasal and nasal-type|9719/3
C0558916|T191|SY|128805001|SNOMEDCT_US|T/NK-cell lymphoma|9719/3
C0392788|T191|SY|414166008|SNOMEDCT_US|T/NK-cell lymphoma|9719/3
C0558916|T191|SY|128805001|SNOMEDCT_US|T/NK-cell lymphoma, nasal and nasal type|9719/3
C2699747|T191|PT|C80374|NCI|Systemic EBV-Positive T-Cell Lymphoma of Childhood|9724/3
C2699747|T191|OP|C80374|NCI|Systemic EBV-Positive T-Cell Lymphoproliferative Disorder of Childhood|9724/3
C2699747|T191|PT|C80374|NCI_NICHD|Systemic EBV-Positive T-Cell Lymphoproliferative Disease of Childhood|9724/3
C2699747|T191|PT|450906003|SNOMEDCT_US|Systemic EBV positive T-cell lymphoproliferative disease of childhood|9724/3
C2699747|T191|SY|450906003|SNOMEDCT_US|Systemic Epstein Barr virus positive T-cell lymphoproliferative disease of childhood|9724/3
C1708397|T191|PT|368033|MEDCIN|Hydroa vacciniforme-like lymphoma|9725/3
C1708397|T191|OP|C45327|NCI|Hydroa Vacciniforme-Like Cutaneous T-Cell Lymphoma|9725/3
C1708397|T191|OP|C45327|NCI|Hydroa Vacciniforme-Like Lymphoma|9725/3
C1708397|T191|PT|C45327|NCI|Hydroa Vacciniforme-Like Lymphoproliferative Disorder|9725/3
C1708397|T191|SY|C45327|NCI_NICHD|HV-Like Lymphoma|9725/3
C1708397|T191|PT|C45327|NCI_NICHD|Hydroa Vacciniforme-Like Lymphoma|9725/3
C1708397|T191|PT|763719001|SNOMEDCT_US|Hydroa vacciniforme-like lymphoma|9725/3
C1708397|T191|PT|450907007|SNOMEDCT_US|Hydroa vacciniforme-like lymphoma|9725/3
C1708397|T191|PT|789440003|SNOMEDCT_US|Hydroa vacciniforme-like lymphoproliferative disorder|9725/3
C1707547|T191|PT|392177|MEDCIN|Primary cutaneous gamma-delta-positive T-cell lymphoma|9726/3
C1707547|T191|SY|392177|MEDCIN|skin malignant lymphoma mature T-cell cutaneous primary gamma-delta-positive|9726/3
C1707547|T191|SY|C45340|NCI|Cutaneous Gamma/Delta T-Cell Lymphoma|9726/3
C1707547|T191|SY|C45340|NCI|Peripheral Gamma-Delta T-Cell Lymphoma|9726/3
C1707547|T191|PT|C45340|NCI|Primary Cutaneous Gamma-Delta T-Cell Lymphoma|9726/3
C1707547|T191|DN|C45340|NCI_CTRP|Primary Cutaneous Gamma-Delta T-Cell Lymphoma|9726/3
C1707547|T191|PT|450908002|SNOMEDCT_US|Primary cutaneous gamma-delta T-cell lymphoma|9726/3
C1707547|T191|SY|733627006|SNOMEDCT_US|Primary cutaneous gamma-delta T-cell lymphoma|9726/3
C1707547|T191|PT|733627006|SNOMEDCT_US|Primary cutaneous gamma-delta-positive T-cell lymphoma|9726/3
C0079748|T191|PT|0003356|CCPSS|LYMPHOMA LYMPHOBLASTIC|9727/3
C0079748|T191|PT|0000015226|CHV|lymphoblastic lymphoma|9727/3
C0079748|T191|SY|0000015226|CHV|lymphoblastoma|9727/3
C0079748|T191|SY|0000015226|CHV|lymphoma lymphoblastic|9727/3
C1301363|T191|AB|C86.4|ICD10CM|Blastic NK-cell lymphoma|9727/3
C1301363|T191|PT|C86.4|ICD10CM|Blastic NK-cell lymphoma|9727/3
C0079748|T191|ET|C83.5|ICD10CM|Lymphoblastic lymphoma NOS|9727/3
C0079748|T191|PT|MTHU046682|ICPC2ICD10ENG|lymphoblastic; lymphoma|9727/3
C0079748|T191|PT|MTHU046686|ICPC2ICD10ENG|lymphoblastoma|9727/3
C0079748|T191|PT|MTHU046814|ICPC2ICD10ENG|lymphoma; lymphoblastic|9727/3
C0079748|T191|LLT|10065923|MDR|Lymphoblastic lymphoma|9727/3
C1301363|T191|PT|338552|MEDCIN|Blastic NK-cell lymphoma|9727/3
C1301363|T191|PT|357125|MEDCIN|Blastic plasmacytoid dendritic cell neoplasm|9727/3
C1301363|T191|SY|338552|MEDCIN|malignant neoplasm lymphoma nk-cell blastic|9727/3
C1301363|T191|SY|357125|MEDCIN|neoplasm of hematopoietic cell type blastic plasmacytoid dendritic cell|9727/3
C0079748|T191|PN|NOCODE|MTH|Precursor cell lymphoblastic lymphoma|9727/3
C0079748|T191|ET|200.1|MTHICD9|Diffuse lymphoblastic lymphoma|9727/3
C0079748|T191|ET|200.1|MTHICD9|Diffuse lymphoblastic lymphosarcoma|9727/3
C0079748|T191|ET|200.1|MTHICD9|Diffuse lymphoblastic malignant lymphoma|9727/3
C0079748|T191|ET|200.1|MTHICD9|Diffuse lymphoblastoma|9727/3
C0079748|T191|ET|200.1|MTHICD9|Lymphoblastic lymphoma|9727/3
C0079748|T191|ET|200.1|MTHICD9|Lymphoblastic lymphosarcoma|9727/3
C0079748|T191|ET|200.1|MTHICD9|Lymphoblastic malignant lymphoma|9727/3
C0079748|T191|ET|200.1|MTHICD9|Lymphoblastoma|9727/3
C1301363|T191|SY|C7203|NCI|Agranular CD4+ CD56+ Hematodermic Neoplasm/Tumor|9727/3
C1301363|T191|OP|C7203|NCI|Agranular CD4+ Natural Killer Cell Leukemia|9727/3
C1301363|T191|OP|C7203|NCI|Blastic Natural Killer Leukemia/Lymphoma|9727/3
C1301363|T191|OP|C7203|NCI|Blastic NK-Cell Lymphoma|9727/3
C1301363|T191|PT|C7203|NCI|Blastic Plasmacytoid Dendritic Cell Neoplasm|9727/3
C1301363|T191|SY|TCGA|NCI|Blastic Plasmacytoid Dendritic Cell Neoplasm|9727/3
C1301363|T191|AB|C7203|NCI|BPDCN|9727/3
C1301363|T191|SY|C7203|NCI|CD4+/CD56+ Hematodermic Neoplasm|9727/3
C0079748|T191|PT|C9360|NCI|Lymphoblastic Lymphoma|9727/3
C1301363|T191|OP|C7203|NCI|Monomorphic NK-Cell Lymphoma|9727/3
C0079748|T191|SY|C9360|NCI|Precursor Cell Lymphoblastic Lymphoma|9727/3
C0079748|T191|SY|C9360|NCI|Precursor Lymphoblastic Lymphoma|9727/3
C0079748|T191|PT|C9360|NCI_CDISC|LYMPHOMA, LYMPHOBLASTIC, MALIGNANT|9727/3
C0079748|T191|SY|C9360|NCI_CDISC|Precursor Cell Lymphoblastic Lymphoma|9727/3
C0079748|T191|SY|C9360|NCI_CDISC|Precursor Lymphoblastic Lymphoma|9727/3
C0079748|T191|PT|C9360|NCI_CPTAC|Lymphoblastic Lymphoma|9727/3
C1301363|T191|DN|C7203|NCI_CTRP|Blastic Plasmacytoid Dendritic Cell Neoplasm|9727/3
C0079748|T191|DN|C9360|NCI_CTRP|Lymphoblastic Lymphoma|9727/3
C0079748|T191|PT|CDR0000597158|NCI_NCI-GLOSS|lymphoblastic lymphoma|9727/3
C0079748|T191|PT|CDR0000597159|NCI_NCI-GLOSS|precursor lymphoblastic lymphoma|9727/3
C1301363|T191|SY|CDR0000671060|PDQ|blastic NK-cell lymphoma|9727/3
C1301363|T191|PT|CDR0000671060|PDQ|blastic plasmacytoid dendritic cell neoplasm|9727/3
C0079748|T191|SY|Xa0TP|RCD|Lymphoblastic lymphoma|9727/3
C0079748|T191|SY|B6274|RCD|Lymphoblastic lymphosarcoma|9727/3
C0079748|T191|SY|Xa0TP|RCD|Lymphoblastoma|9727/3
C0079748|T191|AB|Xa0TP|RCD|Malig lymphoma - lymphoblastic|9727/3
C0079748|T191|PT|Xa0TP|RCD|Malignant lymphoma - lymphoblastic|9727/3
C0079748|T191|IS|BBgG.|RCDSY|Lymphoblastic lymphoma NOS|9727/3
C1301363|T191|OAP|397354007|SNOMEDCT_US|Blastic NK-cell lymphoma|9727/3
C1301363|T191|PT|445105005|SNOMEDCT_US|Blastic plasmacytoid dendritic cell neoplasm|9727/3
C1301363|T191|PT|445030005|SNOMEDCT_US|Blastic plasmacytoid dendritic cell neoplasm|9727/3
C0079748|T191|SY|109965004|SNOMEDCT_US|Diffuse non-Hodgkin lymphoma, lymphoblastic|9727/3
C0079748|T191|SY|109965004|SNOMEDCT_US|Diffuse non-Hodgkin's lymphoma, lymphoblastic|9727/3
C0079748|T191|SY|109965004|SNOMEDCT_US|Lymphoblastic lymphoma|9727/3
C0079748|T191|SY|109965004|SNOMEDCT_US|Lymphoblastic lymphoma, diffuse|9727/3
C0079748|T191|SY|188675007|SNOMEDCT_US|Lymphoblastic lymphosarcoma|9727/3
C0079748|T191|IS|8175003|SNOMEDCT_US|Lymphoblastoma|9727/3
C0079748|T191|SY|109965004|SNOMEDCT_US|Lymphoblastoma|9727/3
C0079748|T191|SY|109965004|SNOMEDCT_US|Malignant lymphoma - lymphoblastic|9727/3
C0079748|T191|IS|8175003|SNOMEDCT_US|Malignant lymphoma, convoluted cell|9727/3
C0079748|T191|OAP|8175003|SNOMEDCT_US|Malignant lymphoma, lymphoblastic|9727/3
C0079748|T191|SY|128806000|SNOMEDCT_US|Malignant lymphoma, lymphoblastic|9727/3
C0079748|T191|IS|8175003|SNOMEDCT_US|Malignant lymphoma, lymphoblastic -RETIRED-|9727/3
C0079748|T191|OF|8175003|SNOMEDCT_US|Malignant lymphoma, lymphoblastic -RETIRED-|9727/3
C0079748|T191|PT|128806000|SNOMEDCT_US|Precursor cell lymphoblastic lymphoma|9727/3
C0855146|T191|PT|10036523|MDR|Precursor B-lymphoblastic lymphoma|9728/3
C0855146|T191|LLT|10036523|MDR|Precursor B-lymphoblastic lymphoma|9728/3
C0855146|T191|LLT|10036525|MDR|Precursor B-lymphoblastic lymphoma NOS|9728/3
C0855146|T191|HT|10036524|MDR|Precursor B-lymphoblastic lymphomas|9728/3
C0855146|T191|PN|NOCODE|MTH|B Lymphoblastic Lymphoma|9728/3
C1292757|T191|PN|NOCODE|MTH|Precursor B-cell lymphoblastic lymphoma|9728/3
C0855146|T191|PT|C8868|NCI|B Lymphoblastic Lymphoma|9728/3
C0855146|T191|SY|C8868|NCI|B-Lymphoblastic Lymphoma|9728/3
C0855146|T191|SY|C8868|NCI|Precursor B-Lymphoblastic Lymphoma|9728/3
C0855146|T191|SY|10036525|NCI_CTEP-SDC|Precur. B-lymphoblastic lymphoma|9728/3
C0855146|T191|PT|10036525|NCI_CTEP-SDC|Precursor B-lymphoblastic lymphoma|9728/3
C0855146|T191|DN|C8868|NCI_CTRP|B Lymphoblastic Lymphoma|9728/3
C1292757|T191|PT|128807009|SNOMEDCT_US|Precursor B-cell lymphoblastic lymphoma|9728/3
C1292758|T191|SY|356964|MEDCIN|malignant neoplasm precursor t-cell lymphoblastic lymphoma|9729/3
C1292758|T191|PT|356964|MEDCIN|malignant precursor T-cell lymphoblastic lymphoma|9729/3
C1292758|T191|PN|NOCODE|MTH|Precursor T-cell lymphoblastic lymphoma|9729/3
C1292758|T191|SY|C6919|NCI|Precursor T Lymphoblastic Lymphoma|9729/3
C1292758|T191|SY|C6919|NCI|Precursor T-Cell Lymphoblastic Lymphoma|9729/3
C1292758|T191|SY|C6919|NCI|Precursor T-Lymphoblastic Lymphoma|9729/3
C1292758|T191|PT|C6919|NCI|T Lymphoblastic Lymphoma|9729/3
C1292758|T191|SY|C6919|NCI|T-Lymphoblastic Lymphoma|9729/3
C1292758|T191|SY|10036545|NCI_CTEP-SDC|Precur. T-lymphoblastic lymphoma|9729/3
C1292758|T191|PT|10036545|NCI_CTEP-SDC|Precursor T-lymphoblastic lymphoma|9729/3
C1292758|T191|DN|C6919|NCI_CTRP|T Lymphoblastic Lymphoma|9729/3
C1292758|T191|PT|CDR0000509757|NCI_NCI-GLOSS|precursor T-lymphoblastic lymphoma|9729/3
C1292758|T191|PT|CDR0000509758|NCI_NCI-GLOSS|T-lymphoblastic lymphoma|9729/3
C1292758|T191|PT|421246008|SNOMEDCT_US|Precursor T-cell lymphoblastic lymphoma|9729/3
C1292758|T191|PT|128808004|SNOMEDCT_US|Precursor T-cell lymphoblastic lymphoma|9729/3
C0474852|T191|PN|NOCODE|MTH|Plasma cell tumor, benign|9731/0
C0474852|T191|PT|BBn1.|RCD|Plasma cell tumour, benign|9731/0
C0474852|T191|SY|BBn1.|RCD|Plasmacytoma, benign|9731/0
C0474852|T191|PT|BBn1.|RCDAE|Plasma cell tumor, benign|9731/0
C0474852|T191|PT|110460003|SNOMEDCT_US|Plasma cell tumor, benign|9731/0
C0474852|T191|PTGB|110460003|SNOMEDCT_US|Plasma cell tumour, benign|9731/0
C0474852|T191|SY|110460003|SNOMEDCT_US|Plasmacytoma, benign|9731/0
C0032131|T191|PT|0014009|CCPSS|PLASMACYTOMA|9731/3
C0032131|T191|SY|0000009812|CHV|bone plasmacytoma|9731/3
C0032131|T191|SY|0000009812|CHV|plasma cell neoplasms|9731/3
C0032131|T191|SY|0000009812|CHV|plasma cell tumor|9731/3
C0032131|T191|SY|0000009812|CHV|plasma cell tumors|9731/3
C0032131|T191|PT|0000009812|CHV|plasmacytoma|9731/3
C0032131|T191|SY|0000009812|CHV|plasmacytomas|9731/3
C0032131|T191|SY|0000009812|CHV|plasmacytomas solitary|9731/3
C0032131|T191|SY|0000009812|CHV|plasmocytoma|9731/3
C0032131|T191|SY|0000009812|CHV|plasmocytomas|9731/3
C0032131|T191|SY|0000009812|CHV|solitary plasmacytoma|9731/3
C0032131|T191|PT|HP:0011857|HPO|Plasmacytoma|9731/3
C0032131|T191|ET|HP:0006775|HPO|Plasmocytoma|9731/3
C0032131|T191|ET|C90.3|ICD10CM|Plasmacytoma NOS|9731/3
C0032131|T191|ET|C90.3|ICD10CM|Solitary myeloma|9731/3
C0032131|T191|AB|C90.3|ICD10CM|Solitary plasmacytoma|9731/3
C0032131|T191|HT|C90.3|ICD10CM|Solitary plasmacytoma|9731/3
C0032131|T191|ET|C90.30|ICD10CM|Solitary plasmacytoma NOS|9731/3
C0032131|T191|PT|MTHU050354|ICPC2ICD10ENG|monostotic; myeloma|9731/3
C0032131|T191|PT|MTHU050355|ICPC2ICD10ENG|monostotic; myeloma, plasma cell|9731/3
C0032131|T191|PT|MTHU050876|ICPC2ICD10ENG|myeloma; monostotic|9731/3
C0032131|T191|PT|MTHU050877|ICPC2ICD10ENG|myeloma; monostotic, plasma cell|9731/3
C0032131|T191|PT|MTHU050878|ICPC2ICD10ENG|myeloma; solitary|9731/3
C0032131|T191|PT|MTHU059929|ICPC2ICD10ENG|plasma cell; tumor|9731/3
C0032131|T191|PT|MTHU059937|ICPC2ICD10ENG|plasmacytoma|9731/3
C0032131|T191|PT|MTHU068378|ICPC2ICD10ENG|solitary; myeloma|9731/3
C0032131|T191|PT|MTHU077140|ICPC2ICD10ENG|tumor; plasma cell|9731/3
C0032131|T191|PT|U003707|LCH|Plasmacytoma|9731/3
C0032131|T191|PT|sh85103091|LCH_NW|Plasmacytoma|9731/3
C0032131|T191|LLT|10035229|MDR|Plasma cell tumor|9731/3
C0032131|T191|LLT|10073875|MDR|Plasma cell tumour|9731/3
C0032131|T191|LLT|10035484|MDR|Plasmacytoma|9731/3
C0032131|T191|PT|10035484|MDR|Plasmacytoma|9731/3
C0032131|T191|PT|31706|MEDCIN|malignant plasmacytoma|9731/3
C0032131|T191|SY|31706|MEDCIN|plasmacytoma|9731/3
C0032131|T191|ET|332|MEDLINEPLUS|Plasmacytoma|9731/3
C0032131|T191|ET|D010954|MSH|Plasma Cell Tumor|9731/3
C0032131|T191|PM|D010954|MSH|Plasma Cell Tumors|9731/3
C0032131|T191|MH|D010954|MSH|Plasmacytoma|9731/3
C0032131|T191|PM|D010954|MSH|Plasmacytomas|9731/3
C0032131|T191|ET|D010954|MSH|Plasmocytoma|9731/3
C0032131|T191|PM|D010954|MSH|Plasmocytomas|9731/3
C0032131|T191|PM|D010954|MSH|Tumor, Plasma Cell|9731/3
C0032131|T191|PM|D010954|MSH|Tumors, Plasma Cell|9731/3
C0032131|T191|PN|NOCODE|MTH|Plasmacytoma|9731/3
C1532560|T191|PN|NOCODE|MTH|Plasmacytoma - category|9731/3
C0032131|T191|ET|238.6|MTHICD9|Plasmacytoma NOS|9731/3
C0032131|T191|ET|238.6|MTHICD9|Solitary myeloma|9731/3
C0032131|T191|PT|C9349|NCI|Plasmacytoma|9731/3
C0032131|T191|PT|C6932|NCI|Solitary Plasmacytoma|9731/3
C0032131|T191|PT|C9349|NCI_CPTAC|Plasmacytoma|9731/3
C0032131|T191|PT|10035484|NCI_CTEP-SDC|Solitary plasmacytoma|9731/3
C0032131|T191|PT|C9349|NCI_CTRP|Plasmacytoma|9731/3
C0032131|T191|DN|C9349|NCI_CTRP|Plasmacytoma|9731/3
C0032131|T191|PT|CDR0000046231|NCI_NCI-GLOSS|plasmacytoma|9731/3
C0032131|T191|SY|Xa9AA|RCD|Monostotic myeloma|9731/3
C0032131|T191|PT|XM1FQ|RCD|Plasma cell tumour|9731/3
C0032131|T191|PT|Xa9AA|RCD|Plasmacytoma|9731/3
C0032131|T191|OP|XaBLx|RCD|Plasmacytoma NOS|9731/3
C0032131|T191|SY|Xa9AA|RCD|Solitary myeloma|9731/3
C0032131|T191|PT|XM1FQ|RCDAE|Plasma cell tumor|9731/3
C0032131|T191|OP|BBnz.|RCDSA|Plasma cell tumor NOS|9731/3
C0032131|T191|OP|BBn..|RCDSA|Plasma cell tumors|9731/3
C0032131|T191|OP|BBnz.|RCDSY|Plasma cell tumour NOS|9731/3
C0032131|T191|OP|BBn..|RCDSY|Plasma cell tumours|9731/3
C0032131|T191|OP|BBn2.|RCDSY|Plasmacytoma NOS|9731/3
C0032131|T191|OAS|302852008|SNOMEDCT_US|Monostotic myeloma|9731/3
C0032131|T191|OAS|189507001|SNOMEDCT_US|Myeloma - solitary|9731/3
C0032131|T191|OAS|154644004|SNOMEDCT_US|Myeloma, solitary|9731/3
C0032131|T191|OAS|269652000|SNOMEDCT_US|Myeloma, solitary|9731/3
C0032131|T191|OAP|274907000|SNOMEDCT_US|Plasma cell tumor|9731/3
C0032131|T191|SY|10639003|SNOMEDCT_US|Plasma cell tumor|9731/3
C0032131|T191|OAP|274907000|SNOMEDCT_US|Plasma cell tumour|9731/3
C0032131|T191|SYGB|10639003|SNOMEDCT_US|Plasma cell tumour|9731/3
C0032131|T191|OAP|302852008|SNOMEDCT_US|Plasmacytoma|9731/3
C0032131|T191|OAP|188719003|SNOMEDCT_US|Plasmacytoma|9731/3
C0032131|T191|OF|188719003|SNOMEDCT_US|Plasmacytoma|9731/3
C0032131|T191|PT|415112005|SNOMEDCT_US|Plasmacytoma|9731/3
C0032131|T191|PT|10639003|SNOMEDCT_US|Plasmacytoma|9731/3
C1532560|T191|PT|415113000|SNOMEDCT_US|Plasmacytoma - category|9731/3
C0032131|T191|OAS|302852008|SNOMEDCT_US|Plasmacytoma - disorder|9731/3
C0032131|T191|SY|415112005|SNOMEDCT_US|Plasmacytoma - disorder|9731/3
C0032131|T191|OAS|189507001|SNOMEDCT_US|Plasmacytoma NOS|9731/3
C0032131|T191|OF|188720009|SNOMEDCT_US|Plasmacytoma NOS|9731/3
C0032131|T191|OAP|308122007|SNOMEDCT_US|Plasmacytoma NOS|9731/3
C0032131|T191|OAP|188720009|SNOMEDCT_US|Plasmacytoma NOS|9731/3
C0032131|T191|SY|10639003|SNOMEDCT_US|Plasmacytoma of bone|9731/3
C0032131|T191|IS|10639003|SNOMEDCT_US|Plasmacytoma, NOS|9731/3
C0032131|T191|OAS|189507001|SNOMEDCT_US|Solitary myeloma|9731/3
C0032131|T191|OAS|302852008|SNOMEDCT_US|Solitary myeloma|9731/3
C0032131|T191|OAS|269652000|SNOMEDCT_US|Solitary myeloma|9731/3
C0032131|T191|OAS|154644004|SNOMEDCT_US|Solitary myeloma|9731/3
C0032131|T191|SY|10639003|SNOMEDCT_US|Solitary myeloma|9731/3
C0032131|T191|SY|10639003|SNOMEDCT_US|Solitary plasmacytoma|9731/3
C0032131|T191|SY|10639003|SNOMEDCT_US|Solitary plasmacytoma of bone|9731/3
C0026764|T191|ET|0000004636|AOD|multiple myeloma|9732/3
C0026764|T191|PT|0046024|CCPSS|MULTIPLE MYELOMA|9732/3
C0026764|T191|SD|40|CCS|Multiple myeloma|9732/3
C0026764|T191|MD|2.10.4|CCS|Multiple myeloma|9732/3
C0026764|T191|SD|NEO065|CCSR_10|Multiple myeloma|9732/3
C0026764|T191|SY|0000008325|CHV|kahler disease|9732/3
C0026764|T191|SY|0000008325|CHV|kahler's disease|9732/3
C0026764|T191|SY|0000008325|CHV|multiple myeloma|9732/3
C0026764|T191|SY|0000008325|CHV|multiple myelomas|9732/3
C0026764|T191|SY|0000008325|CHV|multiple myelomatosis|9732/3
C0026764|T191|SY|0000008325|CHV|myeloma|9732/3
C0026764|T191|SY|0000008325|CHV|myelomas|9732/3
C0026764|T191|SY|0000008325|CHV|myelomatosis|9732/3
C0026764|T191|SY|0000008325|CHV|plasma cell myeloma|9732/3
C0026764|T191|SY|0000008325|CHV|plasma cell neoplasms|9732/3
C0026764|T191|PT|496|COSTAR|MULTIPLE MYELOMA|9732/3
C0026764|T191|PT|2004-0850|CSP|multiple myeloma|9732/3
C0026764|T191|ET|2004-0850|CSP|myeloma|9732/3
C0026764|T191|ET|2004-0850|CSP|myelomatosis|9732/3
C0026764|T191|ET|2004-0850|CSP|plasma cell myeloma|9732/3
C0026764|T191|GT|MYELOMA|CST|MULTIPLE MYELOMA|9732/3
C0026764|T191|GT|MYELOMA|CST|MULTIPLE MYELOMA MYELOMATOSIS|9732/3
C0026764|T191|PT|MYELOMA|CST|MYELOMA|9732/3
C0026764|T191|GT|MYELOMA|CST|MYELOMATOSIS MULTIPLE|9732/3
C0026764|T191|SY|NOCODE|DXP|KAHLER DISEASE|9732/3
C0026764|T191|SY|NOCODE|DXP|KAHLER-BOZZOLO DISEASE|9732/3
C0026764|T191|DI|U001237|DXP|MYELOMA, MULTIPLE|9732/3
C0026764|T191|ET|HP:0006775|HPO|Kahler's disease|9732/3
C0026764|T191|PT|HP:0006775|HPO|Multiple myeloma|9732/3
C0026764|T191|PT|C90.0|ICD10|Multiple myeloma|9732/3
C0026764|T191|ET|C90.0|ICD10CM|Kahler's disease|9732/3
C0026764|T191|HT|C90.0|ICD10CM|Multiple myeloma|9732/3
C0026764|T191|AB|C90.0|ICD10CM|Multiple myeloma|9732/3
C0026764|T191|ET|C90.00|ICD10CM|Multiple myeloma NOS|9732/3
C0026764|T191|ET|C90.0|ICD10CM|Myelomatosis|9732/3
C0026764|T191|ET|C90.0|ICD10CM|Plasma cell myeloma|9732/3
C0026764|T191|HT|203.0|ICD9CM|Multiple myeloma|9732/3
C0026764|T191|PT|MTHU040779|ICPC2ICD10ENG|Kahler|9732/3
C0026764|T191|PT|MTHU050875|ICPC2ICD10ENG|myeloma|9732/3
C0026764|T191|PT|MTHU050866|ICPC2ICD10ENG|myelomata; multiple|9732/3
C0026764|T191|PT|MTHU050867|ICPC2ICD10ENG|myelomatosis|9732/3
C0026764|T191|PTN|B74015|ICPC2P|multiple myeloma|9732/3
C0026764|T191|PT|B74015|ICPC2P|Myeloma;multiple|9732/3
C0026764|T191|PT|U003053|LCH|Multiple myeloma|9732/3
C0026764|T191|PT|sh85088367|LCH_NW|Multiple myeloma|9732/3
C0026764|T191|LA|LA26799-9|LNC|Plasma cell neoplasm|9732/3
C0026764|T191|LLT|10028228|MDR|Multiple myeloma|9732/3
C0026764|T191|OL|10028232|MDR|Multiple myeloma myelomatosis|9732/3
C0026764|T191|LLT|10028566|MDR|Myeloma|9732/3
C0026764|T191|LLT|10028568|MDR|Myelomatosis|9732/3
C0026764|T191|LLT|10028569|MDR|Myelomatosis multiple|9732/3
C0026764|T191|LLT|10034613|MDR|Peripheral plasma cell myeloma|9732/3
C0026764|T191|LLT|10035226|MDR|Plasma cell myeloma|9732/3
C0026764|T191|PT|10035226|MDR|Plasma cell myeloma|9732/3
C0026764|T191|HT|10074470|MDR|Plasma cell myelomas|9732/3
C0026764|T191|PT|31705|MEDCIN|multiple myeloma|9732/3
C0026764|T191|PT|332|MEDLINEPLUS|Multiple Myeloma|9732/3
C0026764|T191|SY|332|MEDLINEPLUS|Plasma-cell myeloma|9732/3
C0026764|T191|ET|332|MEDLINEPLUS|Plasma-cell Myeloma|9732/3
C0026764|T191|PM|D009101|MSH|Cell Myeloma, Plasma|9732/3
C0026764|T191|PM|D009101|MSH|Cell Myelomas, Plasma|9732/3
C0026764|T191|PM|D009101|MSH|Disease, Kahler|9732/3
C0026764|T191|ET|D009101|MSH|Kahler Disease|9732/3
C0026764|T191|MH|D009101|MSH|Multiple Myeloma|9732/3
C0026764|T191|PM|D009101|MSH|Multiple Myelomas|9732/3
C0026764|T191|PM|D009101|MSH|Myeloma Multiple|9732/3
C0026764|T191|ET|D009101|MSH|Myeloma-Multiple|9732/3
C0026764|T191|PM|D009101|MSH|Myeloma-Multiples|9732/3
C0026764|T191|ET|D009101|MSH|Myeloma, Multiple|9732/3
C0026764|T191|PM|D009101|MSH|Myeloma, Plasma Cell|9732/3
C0026764|T191|ET|D009101|MSH|Myeloma, Plasma-Cell|9732/3
C0026764|T191|PM|D009101|MSH|Myelomas, Multiple|9732/3
C0026764|T191|PM|D009101|MSH|Myelomas, Plasma Cell|9732/3
C0026764|T191|PM|D009101|MSH|Myelomas, Plasma-Cell|9732/3
C0026764|T191|PM|D009101|MSH|Myelomatoses|9732/3
C0026764|T191|ET|D009101|MSH|Myelomatosis|9732/3
C0026764|T191|ET|D009101|MSH|Plasma Cell Myeloma|9732/3
C0026764|T191|PM|D009101|MSH|Plasma Cell Myelomas|9732/3
C0026764|T191|PM|D009101|MSH|Plasma-Cell Myeloma|9732/3
C0026764|T191|PM|D009101|MSH|Plasma-Cell Myelomas|9732/3
C0026764|T191|PN|NOCODE|MTH|Multiple Myeloma|9732/3
C0026764|T191|ET|203.0|MTHICD9|Kahler's disease|9732/3
C0026764|T191|ET|203.0|MTHICD9|Myelomatosis|9732/3
C0026764|T191|SY|C3242|NCI|Multiple Myeloma|9732/3
C0026764|T191|SY|C3242|NCI|Myeloma|9732/3
C0026764|T191|PT|C3242|NCI|Plasma Cell Myeloma|9732/3
C0026764|T191|SY|TCGA|NCI|Plasma Cell Myeloma|9732/3
C0026764|T191|SY|C3242|NCI_CDISC|Multiple Myeloma|9732/3
C0026764|T191|SY|C3242|NCI_CDISC|Myeloma|9732/3
C0026764|T191|PT|C3242|NCI_CDISC|MYELOMA, PLASMA CELL, MALIGNANT|9732/3
C0026764|T191|SY|C3242|NCI_CPTAC|Multiple Myeloma|9732/3
C0026764|T191|PT|C3242|NCI_CPTAC|Plasma Cell Myeloma|9732/3
C0026764|T191|PT|10028566|NCI_CTEP-SDC|Myeloma, NOS|9732/3
C0026764|T191|PT|C3242|NCI_CTRP|Multiple Myeloma|9732/3
C0026764|T191|DN|C3242|NCI_CTRP|Multiple Myeloma/Plasma Cell Myeloma|9732/3
C0026764|T191|SY|C3242|NCI_CTRP|Plasma Cell Myeloma|9732/3
C0026764|T191|PT|CDR0000411381|NCI_NCI-GLOSS|Kahler disease|9732/3
C0026764|T191|PT|CDR0000045793|NCI_NCI-GLOSS|multiple myeloma|9732/3
C0026764|T191|PT|CDR0000045795|NCI_NCI-GLOSS|myeloma|9732/3
C0026764|T191|PT|CDR0000411383|NCI_NCI-GLOSS|myelomatosis|9732/3
C0026764|T191|PT|CDR0000411384|NCI_NCI-GLOSS|plasma cell myeloma|9732/3
C0026764|T191|SY|CDR0000037974|PDQ|multiple myeloma|9732/3
C0026764|T191|SY|CDR0000040068|PDQ|multiple myeloma|9732/3
C0026764|T191|PT|CDR0000042947|PDQ|multiple myeloma|9732/3
C0026764|T191|ET|CDR0000037974|PDQ|Multiple myeloma / Plasma cell neoplasm|9732/3
C0026764|T191|PT|CDR0000037974|PDQ|multiple myeloma and other plasma cell neoplasms|9732/3
C0026764|T191|SY|CDR0000042947|PDQ|Myeloma|9732/3
C0026764|T191|SY|CDR0000042947|PDQ|myeloma, multiple|9732/3
C0026764|T191|SY|CDR0000040068|PDQ|myeloma, plasma cell|9732/3
C0026764|T191|SY|CDR0000037974|PDQ|myeloma, plasma cell|9732/3
C0026764|T191|SY|CDR0000040068|PDQ|neoplasm, plasma cell|9732/3
C0026764|T191|SY|CDR0000037974|PDQ|neoplasm, plasma cell|9732/3
C0026764|T191|SY|CDR0000040068|PDQ|plasma cell myeloma|9732/3
C0026764|T191|SY|CDR0000037974|PDQ|plasma cell myeloma|9732/3
C0026764|T191|SY|CDR0000042947|PDQ|Plasma Cell Myeloma|9732/3
C0026764|T191|PT|CDR0000040068|PDQ|plasma cell neoplasm|9732/3
C0026764|T191|SY|CDR0000037974|PDQ|plasma cell neoplasms|9732/3
C0026764|T191|PT|R0121721|QMR|PLASMA CELL MYELOMA|9732/3
C0026764|T191|SY|B630.|RCD|Kahler's disease|9732/3
C0026764|T191|SY|B630.|RCD|Multiple myeloma|9732/3
C0026764|T191|PT|B630.|RCD|Myeloma|9732/3
C0026764|T191|SY|B630.|RCD|Myelomatosis|9732/3
C0026764|T191|IS|BBn0.|RCD|Plasma cell myeloma|9732/3
C0026764|T191|SY|B630.|RCD|Plasmacytic myeloma|9732/3
C0026764|T191|SY|109989006|SNOMEDCT_US|Kahler's disease|9732/3
C0026764|T191|OF|94705007|SNOMEDCT_US|Multiple myeloma|9732/3
C0026764|T191|PT|109989006|SNOMEDCT_US|Multiple myeloma|9732/3
C0026764|T191|PT|55921005|SNOMEDCT_US|Multiple myeloma|9732/3
C0026764|T191|OAP|94705007|SNOMEDCT_US|Multiple myeloma|9732/3
C0026764|T191|SY|55921005|SNOMEDCT_US|Multiple myeloma, no ICD-O subtype|9732/3
C0026764|T191|SY|55921005|SNOMEDCT_US|Multiple myeloma, no International Classification of Diseases for Oncology subtype|9732/3
C0026764|T191|OF|154585004|SNOMEDCT_US|Myeloma|9732/3
C0026764|T191|SY|109989006|SNOMEDCT_US|Myeloma|9732/3
C0026764|T191|SY|55921005|SNOMEDCT_US|Myeloma|9732/3
C0026764|T191|OAP|154585004|SNOMEDCT_US|Myeloma|9732/3
C0026764|T191|IS|55921005|SNOMEDCT_US|Myeloma, NOS|9732/3
C0026764|T191|SY|55921005|SNOMEDCT_US|Myelomatosis|9732/3
C0026764|T191|SY|109989006|SNOMEDCT_US|Myelomatosis|9732/3
C0026764|T191|SY|55921005|SNOMEDCT_US|Plasma cell myeloma|9732/3
C1532559|T191|PT|415109007|SNOMEDCT_US|Plasma cell myeloma - category|9732/3
C0026764|T191|SY|109989006|SNOMEDCT_US|Plasmacytic myeloma|9732/3
C0026764|T191|IT|0583|WHO|MULTIPLE MYELOMA|9732/3
C0026764|T191|PT|0583|WHO|MYELOMATOSIS MULTIPLE|9732/3
C0023484|T191|PT|0044399|CCPSS|LEUKEMIA PLASMA CELL|9733/3
C0023484|T191|SY|0000007349|CHV|cells leukemia plasma|9733/3
C0023484|T191|SY|0000007349|CHV|plasma cell leukaemia|9733/3
C0023484|T191|PT|0000007349|CHV|plasma cell leukemia|9733/3
C0023484|T191|ET|2004-4789|CSP|plasma cell leukemia|9733/3
C0023484|T191|PT|2004-4789|CSP|plasmacytic leukemia|9733/3
C0023484|T191|GT|LEUKEMIA|CST|LEUKEMIA PLASMACYTIC|9733/3
C0023484|T191|DI|U001053|DXP|LEUKEMIA, PLASMA CELL|9733/3
C0023484|T191|SY|NOCODE|DXP|LEUKEMIA, PLASMACYTIC|9733/3
C0023484|T191|PT|C90.1|ICD10|Plasma cell leukaemia|9733/3
C0023484|T191|PT|C90.1|ICD10AE|Plasma cell leukemia|9733/3
C0023484|T191|AB|C90.1|ICD10CM|Plasma cell leukemia|9733/3
C0023484|T191|HT|C90.1|ICD10CM|Plasma cell leukemia|9733/3
C0023484|T191|ET|C90.10|ICD10CM|Plasma cell leukemia NOS|9733/3
C0023484|T191|ET|C90.1|ICD10CM|Plasmacytic leukemia|9733/3
C0023484|T191|HT|203.1|ICD9CM|Plasma cell leukemia|9733/3
C0023484|T191|PT|MTHU044794|ICPC2ICD10ENG|leukemia; plasma cell|9733/3
C0023484|T191|PT|MTHU059925|ICPC2ICD10ENG|plasma cell; leukemia|9733/3
C0023484|T191|PT|sh85103090|LCH_NW|Plasmacytic leukemia|9733/3
C0023484|T191|LLT|10024318|MDR|Leukaemia plasmacytic|9733/3
C0023484|T191|LLT|10024357|MDR|Leukemia plasmacytic|9733/3
C0023484|T191|LLT|10035222|MDR|Plasma cell leukaemia|9733/3
C0023484|T191|PT|10035222|MDR|Plasma cell leukaemia|9733/3
C0023484|T191|LLT|10035223|MDR|Plasma cell leukemia|9733/3
C0023484|T191|MTH_PT|10035222|MDR|Plasma cell leukemia|9733/3
C0023484|T191|SY|97730|MEDCIN|plasma cell leukaemia|9733/3
C0023484|T191|PT|97730|MEDCIN|plasma cell leukemia|9733/3
C0023484|T191|MH|D007952|MSH|Leukemia, Plasma Cell|9733/3
C0023484|T191|ET|D007952|MSH|Leukemia, Plasmacytic|9733/3
C0023484|T191|PM|D007952|MSH|Leukemias, Plasma Cell|9733/3
C0023484|T191|PM|D007952|MSH|Leukemias, Plasmacytic|9733/3
C0023484|T191|ET|D007952|MSH|Plasma Cell Leukemia|9733/3
C0023484|T191|PM|D007952|MSH|Plasma Cell Leukemias|9733/3
C0023484|T191|ET|D007952|MSH|Plasmacytic Leukemia|9733/3
C0023484|T191|PM|D007952|MSH|Plasmacytic Leukemias|9733/3
C0023484|T191|ET|203.1|MTHICD9|Plasmacytic leukemia|9733/3
C0023484|T191|SY|C3180|NCI|Leukemia Plasmacytic|9733/3
C0023484|T191|PT|C3180|NCI|Plasma Cell Leukemia|9733/3
C0023484|T191|SY|C3180|NCI|Plasmacytic Leukemia|9733/3
C0023484|T191|PT|C3180|NCI_CPTAC|Plasma Cell Leukemia|9733/3
C0023484|T191|DN|C3180|NCI_CTRP|Plasma Cell Leukemia|9733/3
C0023484|T191|PT|XaBB3|RCD|Plasma cell leukaemia|9733/3
C0023484|T191|PT|XaBB3|RCDAE|Plasma cell leukemia|9733/3
C0023484|T191|PT|BBr30|RCDSA|Plasma cell leukemia|9733/3
C0023484|T191|OP|BBr3z|RCDSA|Plasma cell leukemia NOS|9733/3
C0023484|T191|OP|BBr3.|RCDSA|Plasma cell leukemias|9733/3
C0023484|T191|PT|BBr30|RCDSY|Plasma cell leukaemia|9733/3
C0023484|T191|OP|BBr3z|RCDSY|Plasma cell leukaemia NOS|9733/3
C0023484|T191|OP|BBr3.|RCDSY|Plasma cell leukaemias|9733/3
C0023484|T191|OAP|188722001|SNOMEDCT_US|Plasma cell leukaemia|9733/3
C0023484|T191|OAP|39193004|SNOMEDCT_US|Plasma cell leukaemia|9733/3
C0023484|T191|PTGB|95210003|SNOMEDCT_US|Plasma cell leukaemia|9733/3
C0023484|T191|OAS|154586003|SNOMEDCT_US|Plasma cell leukaemia|9733/3
C0023484|T191|PTGB|128922003|SNOMEDCT_US|Plasma cell leukaemia|9733/3
C0023484|T191|OAS|269630009|SNOMEDCT_US|Plasma cell leukaemia|9733/3
C0023484|T191|OF|188722001|SNOMEDCT_US|Plasma cell leukaemia|9733/3
C0023484|T191|IS|39193004|SNOMEDCT_US|Plasma cell leukaemia -RETIRED-|9733/3
C0023484|T191|SYGB|95210003|SNOMEDCT_US|Plasma cell leukaemia, disease|9733/3
C0023484|T191|SYGB|128922003|SNOMEDCT_US|Plasma cell leukaemia, morphology|9733/3
C0023484|T191|PT|95210003|SNOMEDCT_US|Plasma cell leukemia|9733/3
C0023484|T191|OAP|39193004|SNOMEDCT_US|Plasma cell leukemia|9733/3
C0023484|T191|PT|128922003|SNOMEDCT_US|Plasma cell leukemia|9733/3
C0023484|T191|OAP|188722001|SNOMEDCT_US|Plasma cell leukemia|9733/3
C0023484|T191|OAS|269630009|SNOMEDCT_US|Plasma cell leukemia|9733/3
C0023484|T191|OAS|154586003|SNOMEDCT_US|Plasma cell leukemia|9733/3
C0023484|T191|IS|39193004|SNOMEDCT_US|Plasma cell leukemia -RETIRED-|9733/3
C0023484|T191|OF|39193004|SNOMEDCT_US|Plasma cell leukemia -RETIRED-|9733/3
C0023484|T191|SY|95210003|SNOMEDCT_US|Plasma cell leukemia, disease|9733/3
C0023484|T191|SY|128922003|SNOMEDCT_US|Plasma cell leukemia, morphology|9733/3
C0023484|T191|SYGB|128922003|SNOMEDCT_US|Plasmacytic leukaemia|9733/3
C0023484|T191|IS|39193004|SNOMEDCT_US|Plasmacytic leukemia|9733/3
C0023484|T191|SY|128922003|SNOMEDCT_US|Plasmacytic leukemia|9733/3
C0278619|T191|PT|0000027203|CHV|extramedullary plasmacytoma|9734/3
C0278619|T191|PT|C90.2|ICD10|Plasmacytoma, extramedullary|9734/3
C0278619|T191|AB|C90.2|ICD10CM|Extramedullary plasmacytoma|9734/3
C0278619|T191|HT|C90.2|ICD10CM|Extramedullary plasmacytoma|9734/3
C0278619|T191|ET|C90.20|ICD10CM|Extramedullary plasmacytoma NOS|9734/3
C0278619|T191|LLT|10066883|MDR|Extramedullary plasmacytoma|9734/3
C0278619|T191|PT|271576|MEDCIN|extramedullary plasmacytoma|9734/3
C1275323|T191|PT|357443|MEDCIN|Primary cutaneous plasmacytoma|9734/3
C1275323|T191|SY|357443|MEDCIN|skin malignant lymphoma non-hodgkin's primary cutaneous plasmacytoma|9734/3
C0278619|T191|PN|NOCODE|MTH|Extramedullary Plasmacytoma|9734/3
C0278619|T191|SY|C4002|NCI|Extramedullary Plasmacytoma|9734/3
C0278619|T191|PT|C4002|NCI|Extraosseous Plasmacytoma|9734/3
C0278619|T191|SY|TCGA|NCI|Extraosseous Plasmacytoma|9734/3
C0278619|T191|DN|C4002|NCI_CTRP|Extraosseous Plasmacytoma|9734/3
C0278619|T191|PT|CDR0000041865|PDQ|extramedullary plasmacytoma|9734/3
C0278619|T191|SY|CDR0000041865|PDQ|Extraosseous Plasmacytoma|9734/3
C0278619|T191|SY|CDR0000041865|PDQ|plasmacytoma, extramedullary|9734/3
C0278619|T191|AB|B6300|RCD|M plsma cel neo,extram p'cytom|9734/3
C0278619|T191|PT|B6300|RCD|Malignant plasma cell neoplasm, extramedullary plasmacytoma|9734/3
C0278619|T191|PT|188718006|SNOMEDCT_US|Extramedullary plasmacytoma|9734/3
C0278619|T191|IS|10639003|SNOMEDCT_US|Extramedullary plasmacytoma|9734/3
C0278619|T191|SY|128921005|SNOMEDCT_US|Extramedullary plasmacytoma|9734/3
C0278619|T191|SY|188718006|SNOMEDCT_US|Malignant plasma cell neoplasm, extramedullary plasmacytoma|9734/3
C1275323|T191|SY|404142007|SNOMEDCT_US|Primary cutaneous plasmacytic B-cell lymphoma|9734/3
C1275323|T191|PT|418789003|SNOMEDCT_US|Primary cutaneous plasmacytoma|9734/3
C1275323|T191|PT|404142007|SNOMEDCT_US|Primary cutaneous plasmacytoma|9734/3
C3472614|T191|ET|C83.3|ICD10CM|Plasmablastic diffuse large B-cell lymphoma|9735/3
C3472614|T191|PT|10065039|MDR|Plasmablastic lymphoma|9735/3
C3472614|T191|LLT|10065039|MDR|Plasmablastic lymphoma|9735/3
C3472614|T191|PT|391490|MEDCIN|Plasmablastic lymphoma|9735/3
C3472614|T191|PM|D000069293|MSH|Lymphoma, Plasmablastic|9735/3
C3472614|T191|PM|D000069293|MSH|Lymphomas, Plasmablastic|9735/3
C3472614|T191|PM|D000069293|MSH|Plasmablastic Diffuse Large B cell Lymphoma|9735/3
C3472614|T191|ET|D000069293|MSH|Plasmablastic Diffuse Large B-cell Lymphoma|9735/3
C3472614|T191|MH|D000069293|MSH|Plasmablastic Lymphoma|9735/3
C3472614|T191|PM|D000069293|MSH|Plasmablastic Lymphomas|9735/3
C3472614|T191|PM|D000069293|MSH|Plasmablasts Diffuse Large B cell Lymphoma|9735/3
C3472614|T191|ET|D000069293|MSH|Plasmablasts Diffuse Large B-cell Lymphoma|9735/3
C3472614|T191|PN|NOCODE|MTH|Plasmablastic lymphoma|9735/3
C3472614|T191|AB|C7224|NCI|PBL|9735/3
C3472614|T191|PT|C7224|NCI|Plasmablastic Lymphoma|9735/3
C3472614|T191|PT|724648008|SNOMEDCT_US|Plasmablastic lymphoma|9735/3
C3472614|T191|PT|450909005|SNOMEDCT_US|Plasmablastic lymphoma|9735/3
C1333294|T191|PT|366458|MEDCIN|Anaplastic lymphoma kinase positive large B-cell lymphoma|9737/3
C1333294|T191|AB|C7225|NCI|ALK-DLBCL|9737/3
C1333294|T191|PT|C7225|NCI|ALK-Positive Large B-Cell Lymphoma|9737/3
C1333294|T191|SY|C7225|NCI|Diffuse Large B-Cell Lymphoma with Expression of Full-Length ALK|9737/3
C1333294|T191|SY|C7225|NCI|Diffuse Large B-Cell Lymphoma with Expression of Full-Length Anaplastic Lymphoma Kinase|9737/3
C1333294|T191|PT|450910000|SNOMEDCT_US|ALK positive large B-cell lymphoma|9737/3
C1333294|T191|PT|715950008|SNOMEDCT_US|ALK-positive large B-cell lymphoma|9737/3
C1333294|T191|SY|715950008|SNOMEDCT_US|Anaplastic lymphoma kinase positive large B-cell lymphoma|9737/3
C1333294|T191|SY|450910000|SNOMEDCT_US|Anaplastic lymphoma kinase positive large B-cell lymphoma|9737/3
C3472615|T191|PT|C27856|NCI|Diffuse Large B-Cell Lymphoma Arising in HHV8-Positive Multicentric Castleman Disease|9738/3
C3472615|T191|SY|C27856|NCI|Kaposi Sarcoma-Associated Human Herpes Virus 8 Positive Extracavity Lymphoma|9738/3
C3472615|T191|SY|C27856|NCI|Kaposi's Sarcoma-Associated Human Herpes Virus 8 Positive Extracavity Lymphoma|9738/3
C3472615|T191|SY|C27856|NCI|Kaposi's Sarcoma-Associated Human Herpes Virus 8+ Extracavity Lymphoma|9738/3
C3472615|T191|AB|C27856|NCI|KSHV-8 Positive Extracavity Lymphoma|9738/3
C3472615|T191|AB|C27856|NCI|KSHV-8+ Extracavity Lymphoma|9738/3
C3472615|T191|SY|C27856|NCI|KSHV-Associated Non-Hodgkin Lymphoma|9738/3
C3472615|T191|SY|C27856|NCI|Large B-Cell Lymphoma Arising in HHV 8-Associated Multicentric Castleman Disease|9738/3
C3472615|T191|SY|C27856|NCI|Large B-Cell Lymphoma Arising in HHV8-Associated Multicentric Castleman Disease|9738/3
C3472615|T191|SY|C27856|NCI|Large B-Cell Lymphoma Arising in Human Herpes Virus 8-Associated Multicentric Castleman Disease|9738/3
C3472615|T191|DN|C27856|NCI_CTRP|Diffuse Large B-Cell Lymphoma Arising in HHV8-Positive Multicentric Castleman Disease|9738/3
C3472615|T191|PT|450911001|SNOMEDCT_US|Large B-cell lymphoma arising in HHV8 associated multicentric Castleman disease|9738/3
C3472615|T191|SY|450911001|SNOMEDCT_US|Large B-cell lymphoma arising in human herpesvirus type 8 associated multicentric Castleman disease|9738/3
C0042111|T191|PT|0035296|CCPSS|URTICARIA PIGMENTOSA|9740/1
C0042111|T191|SY|0000012811|CHV|pigmentosa urticaria|9740/1
C0042111|T191|SY|0000012811|CHV|urticaria pigmentosa|9740/1
C0024897|T191|SY|2004-8021|CSP|mastocytoma|9740/1
C0042111|T191|PT|2716-7072|CSP|urticaria pigmentosa|9740/1
C0042111|T191|DI|U001972|DXP|URTICARIA PIGMENTOSA|9740/1
C1136033|T191|PT|HP:0200151|HPO|Cutaneous mastocytosis|9740/1
C1136033|T191|AB|D47.01|ICD10CM|Cutaneous mastocytosis|9740/1
C1136033|T191|PT|D47.01|ICD10CM|Cutaneous mastocytosis|9740/1
C0024901|T191|ET|D47.01|ICD10CM|Diffuse cutaneous mastocytosis|9740/1
C0272202|T191|ET|D47.09|ICD10CM|Extracutaneous mastocytoma|9740/1
C0042111|T191|ET|D47.01|ICD10CM|Maculopapular cutaneous mastocytosis|9740/1
C0024897|T191|ET|D47.09|ICD10CM|Mastocytoma NOS|9740/1
C0343115|T191|ET|D47.01|ICD10CM|Solitary mastocytoma|9740/1
C0042111|T191|ET|D47.01|ICD10CM|Urticaria pigmentosa|9740/1
C0024897|T191|PT|MTHU047644|ICPC2ICD10ENG|mastocytoma|9740/1
C0042111|T191|PT|MTHU059456|ICPC2ICD10ENG|pigmentation; congenital, urticaria pigmentosa|9740/1
C0042111|T191|PT|MTHU059476|ICPC2ICD10ENG|pigmentosa; urticaria|9740/1
C0042111|T191|PT|MTHU078316|ICPC2ICD10ENG|urticaria; pigmentosa|9740/1
C0024901|T191|LLT|10012812|MDR|Diffuse cutaneous mastocytosis|9740/1
C0024901|T191|PT|10012812|MDR|Diffuse cutaneous mastocytosis|9740/1
C0024897|T191|PT|10026890|MDR|Mastocytoma|9740/1
C0024897|T191|LLT|10026890|MDR|Mastocytoma|9740/1
C0042111|T191|PT|10046752|MDR|Urticaria pigmentosa|9740/1
C0042111|T191|LLT|10046752|MDR|Urticaria pigmentosa|9740/1
C1136033|T191|PT|365415|MEDCIN|cutaneous mastocytosis|9740/1
C0024901|T191|PT|365416|MEDCIN|Diffuse cutaneous mastocytosis|9740/1
C0272202|T191|PT|353717|MEDCIN|Localized extracutaneous mastocytosis|9740/1
C0042111|T191|PT|365417|MEDCIN|maculopapular cutaneous mastocytosis|9740/1
C0343115|T191|PT|356411|MEDCIN|Mast cell nevus|9740/1
C0024897|T191|PT|213227|MEDCIN|mastocytoma|9740/1
C0272202|T191|SY|353717|MEDCIN|mastocytosis - localized extracutaneous|9740/1
C0343115|T191|SY|356411|MEDCIN|neoplasm of mast cell nevus|9740/1
C0024901|T191|SY|365416|MEDCIN|neoplasm uncert behav of histio & mast cells diffuse cutaneous mastocytosis|9740/1
C0042111|T191|SY|365417|MEDCIN|neoplasm uncert behav of histio & mast cells maculopap cutaneous mastocytosis|9740/1
C1136033|T191|SY|365415|MEDCIN|neoplasm uncert behavior of histiocytic & mast cells cutaneous mastocytosis|9740/1
C0343115|T191|PT|356412|MEDCIN|Solitary cutaneous mastocytoma|9740/1
C0042111|T191|PT|33124|MEDCIN|urticaria pigmentosa|9740/1
C1136033|T191|PM|D034701|MSH|Cutaneous Mastocytoses|9740/1
C0024901|T191|PM|D034701|MSH|Cutaneous Mastocytoses, Diffuse|9740/1
C0042111|T191|PM|D014582|MSH|Cutaneous Mastocytoses, Maculopapular|9740/1
C1136033|T191|ET|D034701|MSH|Cutaneous Mastocytosis|9740/1
C0024901|T191|PM|D034701|MSH|Cutaneous Mastocytosis, Diffuse|9740/1
C0042111|T191|PM|D014582|MSH|Cutaneous Mastocytosis, Maculopapular|9740/1
C0272202|T191|PEP|D034801|MSH|Extracutaneous Mastocytoma|9740/1
C0272202|T191|PM|D034801|MSH|Extracutaneous Mastocytomas|9740/1
C0042111|T191|PM|D014582|MSH|Maculopapular Cutaneous Mastocytoses|9740/1
C0042111|T191|ET|D014582|MSH|Maculopapular Cutaneous Mastocytosis|9740/1
C0272202|T191|ET|D034801|MSH|Mastocytoma, Extracutaneous|9740/1
C0343115|T191|MH|D054705|MSH|Mastocytoma, Skin|9740/1
C0272202|T191|PM|D034801|MSH|Mastocytomas, Extracutaneous|9740/1
C1136033|T191|PM|D034701|MSH|Mastocytoses, Cutaneous|9740/1
C1136033|T191|PM|D034701|MSH|Mastocytoses, Skin|9740/1
C1136033|T191|MH|D034701|MSH|Mastocytosis, Cutaneous|9740/1
C0024901|T191|PEP|D034701|MSH|Mastocytosis, Diffuse Cutaneous|9740/1
C1136033|T191|PM|D034701|MSH|Mastocytosis, Skin|9740/1
C0343115|T191|ET|D054705|MSH|Skin Mastocytoma|9740/1
C1136033|T191|PM|D034701|MSH|Skin Mastocytoses|9740/1
C1136033|T191|ET|D034701|MSH|Skin Mastocytosis|9740/1
C0343115|T191|ET|D054705|MSH|Solitary Mastocytoma of Skin|9740/1
C0042111|T191|MH|D014582|MSH|Urticaria Pigmentosa|9740/1
C1136033|T191|PN|NOCODE|MTH|Cutaneous Mastocytosis|9740/1
C0024897|T191|PN|NOCODE|MTH|Mastocytoma|9740/1
C0343115|T191|PN|NOCODE|MTH|Skin Mastocytoma|9740/1
C0042111|T191|PN|NOCODE|MTH|Urticaria Pigmentosa|9740/1
C0024897|T191|ET|238.5|MTHICD9|Mastocytoma NOS|9740/1
C0042111|T191|ET|757.33|MTHICD9|Urticaria pigmentosa|9740/1
C1136033|T191|AB|C7137|NCI|CM|9740/1
C1136033|T191|PT|C7137|NCI|Cutaneous Mastocytosis|9740/1
C0343115|T191|SY|C7138|NCI|Cutaneous Solitary Mastocytoma|9740/1
C0024901|T191|PT|C3218|NCI|Diffuse Cutaneous Mastocytosis|9740/1
C0272202|T191|PT|C7136|NCI|Extracutaneous Mastocytoma|9740/1
C0024897|T191|PT|C9303|NCI|Mastocytoma|9740/1
C0343115|T191|SY|C7138|NCI|Skin Solitary Mastocytoma|9740/1
C0343115|T191|SY|C7138|NCI|Solitary Mastocytoma of Skin|9740/1
C0343115|T191|PT|C7138|NCI|Solitary Mastocytoma of the Skin|9740/1
C0042111|T191|AB|C3433|NCI|UP/MPCM|9740/1
C0042111|T191|SY|C3433|NCI|Urticaria Pigmentosa|9740/1
C0042111|T191|PT|C3433|NCI|Urticaria Pigmentosa/Maculopapular Cutaneous Mastocytosis|9740/1
C0272202|T191|DN|C7136|NCI_CTRP|Extracutaneous Mastocytoma|9740/1
C0042111|T191|DN|C3433|NCI_CTRP|Urticaria Pigmentosa/Maculopapular Cutaneous Mastocytosis|9740/1
C0024897|T191|PT|CDR0000044607|NCI_NCI-GLOSS|mastocytoma|9740/1
C1136033|T191|AB|CDR0000553272|PDQ|CM|9740/1
C1136033|T191|PT|CDR0000553272|PDQ|cutaneous mastocytosis|9740/1
C0272202|T191|PT|CDR0000701775|PDQ|extracutaneous mastocytoma|9740/1
C0042111|T191|AB|CDR0000553281|PDQ|UP/MPCM|9740/1
C0042111|T191|SY|CDR0000553281|PDQ|Urticaria Pigmentosa|9740/1
C0042111|T191|PT|CDR0000553281|PDQ|urticaria pigmentosa/maculopapular cutaneous mastocytosis|9740/1
C0343115|T191|PT|X50KK|RCD|Mast cell naevus|9740/1
C0024897|T191|PT|Xa9AC|RCD|Mastocytoma|9740/1
C0343115|T191|SY|X50KK|RCD|Mastocytoma of skin|9740/1
C0042111|T191|PT|PH321|RCD|Urticaria pigmentosa|9740/1
C0343115|T191|PT|X50KK|RCDAE|Mast cell nevus|9740/1
C0024897|T191|OP|BBp0.|RCDSY|Mastocytoma NOS|9740/1
C0343115|T191|SY|397013007|SNOMEDCT_US|Cutaneous mastocytoma|9740/1
C1136033|T191|PT|703827008|SNOMEDCT_US|Cutaneous mastocytosis|9740/1
C1136033|T191|PT|397012002|SNOMEDCT_US|Cutaneous mastocytosis|9740/1
C0024901|T191|PT|703826004|SNOMEDCT_US|Diffuse cutaneous mastocytosis|9740/1
C0272202|T191|SY|63175003|SNOMEDCT_US|Extracutaneous mastocytoma|9740/1
C0042111|T191|SYGB|78745000|SNOMEDCT_US|Localised cutaneous mastocytosis|9740/1
C0272202|T191|PTGB|63175003|SNOMEDCT_US|Localised extracutaneous mastocytosis|9740/1
C0042111|T191|SY|78745000|SNOMEDCT_US|Localized cutaneous mastocytosis|9740/1
C0042111|T191|IS|78745000|SNOMEDCT_US|Localized cutaneous mastocytosis, NOS|9740/1
C0272202|T191|PT|63175003|SNOMEDCT_US|Localized extracutaneous mastocytosis|9740/1
C0343115|T191|IS|404171008|SNOMEDCT_US|Mast cell naevus|9740/1
C0343115|T191|PTGB|239147000|SNOMEDCT_US|Mast cell naevus|9740/1
C0343115|T191|PT|239147000|SNOMEDCT_US|Mast cell nevus|9740/1
C0343115|T191|IS|404171008|SNOMEDCT_US|Mast cell nevus|9740/1
C0024897|T191|PT|404171008|SNOMEDCT_US|Mastocytoma|9740/1
C0024897|T191|PT|89796001|SNOMEDCT_US|Mastocytoma|9740/1
C0024897|T191|OAP|134333006|SNOMEDCT_US|Mastocytoma|9740/1
C0024897|T191|OF|134333006|SNOMEDCT_US|Mastocytoma|9740/1
C0024897|T191|OAS|189506005|SNOMEDCT_US|Mastocytoma NOS|9740/1
C0343115|T191|SY|239147000|SNOMEDCT_US|Mastocytoma of skin|9740/1
C0024897|T191|IS|89796001|SNOMEDCT_US|Mastocytoma, NOS|9740/1
C0343115|T191|PT|397013007|SNOMEDCT_US|Solitary cutaneous mastocytoma|9740/1
C0343115|T191|SY|397013007|SNOMEDCT_US|Solitary mastocytoma|9740/1
C0343115|T191|PT|703836007|SNOMEDCT_US|Solitary mastocytoma of skin|9740/1
C0042111|T191|OAP|205566001|SNOMEDCT_US|Urticaria pigmentosa|9740/1
C0042111|T191|PT|703828003|SNOMEDCT_US|Urticaria pigmentosa|9740/1
C0042111|T191|PT|78745000|SNOMEDCT_US|Urticaria pigmentosa|9740/1
C0042111|T191|IS|78745000|SNOMEDCT_US|Urticaria pigmentosa, NOS|9740/1
C0036221|T191|PT|C96.2|ICD10|Malignant mast cell tumour|9740/3
C0036221|T191|PT|C96.2|ICD10AE|Malignant mast cell tumor|9740/3
C0036221|T191|AB|C96.2|ICD10CM|Malignant mast cell neoplasm|9740/3
C0036221|T191|HT|C96.2|ICD10CM|Malignant mast cell neoplasm|9740/3
C0036221|T191|AB|C96.22|ICD10CM|Mast cell sarcoma|9740/3
C0036221|T191|PT|C96.22|ICD10CM|Mast cell sarcoma|9740/3
C0036221|T191|HT|202.6|ICD9CM|Malignant mast cell tumors|9740/3
C0036221|T191|PT|MTHU047299|ICPC2ICD10ENG|malignant; mastocytoma|9740/3
C0036221|T191|PT|MTHU048976|ICPC2ICD10ENG|mast cell; sarcoma|9740/3
C0036221|T191|PT|MTHU048978|ICPC2ICD10ENG|mast cell; tumor, malignant|9740/3
C0036221|T191|PT|MTHU047645|ICPC2ICD10ENG|mastocytoma; malignant|9740/3
C0036221|T191|PT|MTHU065922|ICPC2ICD10ENG|sarcoma; mast cell|9740/3
C0036221|T191|PT|MTHU077100|ICPC2ICD10ENG|tumor; mast cell, malignant|9740/3
C0036221|T191|LLT|10025638|MDR|Malignant mast cell neoplasm|9740/3
C0036221|T191|PT|10025638|MDR|Malignant mast cell neoplasm|9740/3
C0036221|T191|OL|10025639|MDR|Malignant mast cell tumors|9740/3
C0036221|T191|MTH_OL|10026708|MDR|Malignant-mast cell tumors|9740/3
C0036221|T191|OL|10026708|MDR|Malignant-mast cell tumours|9740/3
C0036221|T191|PT|338575|MEDCIN|malignant mast cell tumor|9740/3
C0036221|T191|PT|213228|MEDCIN|malignant mastocytoma|9740/3
C0036221|T191|SY|338575|MEDCIN|malignant neoplasm lymphatic/hematopoietic neoplasm mast cell tumor|9740/3
C0036221|T191|PT|272059|MEDCIN|mast cell sarcoma|9740/3
C0036221|T191|PM|D012515|MSH|Malignant Mastocytoma|9740/3
C0036221|T191|PM|D012515|MSH|Malignant Mastocytomas|9740/3
C0036221|T191|PM|D012515|MSH|Mast Cell Sarcoma|9740/3
C0036221|T191|MH|D012515|MSH|Mast-Cell Sarcoma|9740/3
C0036221|T191|PM|D012515|MSH|Mast-Cell Sarcomas|9740/3
C0036221|T191|ET|D012515|MSH|Mastocytoma, Malignant|9740/3
C0036221|T191|PM|D012515|MSH|Mastocytomas, Malignant|9740/3
C0036221|T191|PM|D012515|MSH|Sarcoma, Mast Cell|9740/3
C0036221|T191|ET|D012515|MSH|Sarcoma, Mast-Cell|9740/3
C0036221|T191|PM|D012515|MSH|Sarcomas, Mast-Cell|9740/3
C0036221|T191|PN|NOCODE|MTH|Mast-Cell Sarcoma|9740/3
C0036221|T191|ET|202.6|MTHICD9|Malignant mastocytoma|9740/3
C0036221|T191|ET|202.6|MTHICD9|Mast cell sarcoma|9740/3
C0036221|T191|PT|C9348|NCI|Mast Cell Sarcoma|9740/3
C0036221|T191|SY|TCGA|NCI|Mast Cell Sarcoma|9740/3
C0036221|T191|AB|C9348|NCI|MCS|9740/3
C0036221|T191|DN|C9348|NCI_CTRP|Mast Cell Sarcoma|9740/3
C0036221|T191|PT|CDR0000701774|PDQ|mast cell sarcoma|9740/3
C0036221|T191|AB|CDR0000701774|PDQ|MCS|9740/3
C0036221|T191|SY|XaBAk|RCD|Malignant mast cell tumour|9740/3
C0036221|T191|OP|B626z|RCD|Malignant mast cell tumour NOS|9740/3
C0036221|T191|OP|B626.|RCD|Malignant mast cell tumours|9740/3
C0036221|T191|OA|B6260|RCD|Mast cell malignancy ? site|9740/3
C0036221|T191|OP|B6260|RCD|Mast cell malignancy of unspecified site|9740/3
C0036221|T191|PT|BBp1.|RCD|Mast cell sarcoma|9740/3
C0036221|T191|SY|XaBAk|RCDAE|Malignant mast cell tumor|9740/3
C0036221|T191|OP|B626z|RCDAE|Malignant mast cell tumor NOS|9740/3
C0036221|T191|OP|B626.|RCDAE|Malignant mast cell tumors|9740/3
C0036221|T191|PT|397010005|SNOMEDCT_US|Malignant mast cell neoplasm|9740/3
C0036221|T191|OAS|307591004|SNOMEDCT_US|Malignant mast cell tumor|9740/3
C0036221|T191|SY|13583002|SNOMEDCT_US|Malignant mast cell tumor|9740/3
C0036221|T191|SY|118615008|SNOMEDCT_US|Malignant mast cell tumor|9740/3
C0036221|T191|OAP|188670002|SNOMEDCT_US|Malignant mast cell tumor NOS|9740/3
C0036221|T191|PT|188660004|SNOMEDCT_US|Malignant mast cell tumors|9740/3
C0036221|T191|OAS|307591004|SNOMEDCT_US|Malignant mast cell tumour|9740/3
C0036221|T191|SYGB|13583002|SNOMEDCT_US|Malignant mast cell tumour|9740/3
C0036221|T191|SYGB|118615008|SNOMEDCT_US|Malignant mast cell tumour|9740/3
C0036221|T191|OAP|188670002|SNOMEDCT_US|Malignant mast cell tumour NOS|9740/3
C0036221|T191|PTGB|188660004|SNOMEDCT_US|Malignant mast cell tumours|9740/3
C0036221|T191|SY|13583002|SNOMEDCT_US|Malignant mastocytoma|9740/3
C0036221|T191|OAP|188661000|SNOMEDCT_US|Mast cell malignancy of unspecified site|9740/3
C0036221|T191|SY|118615008|SNOMEDCT_US|Mast cell sarcoma|9740/3
C0036221|T191|PT|13583002|SNOMEDCT_US|Mast cell sarcoma|9740/3
C0272203|T191|ET|D47.02|ICD10CM|Indolent systemic mastocytosis|9741/1
C0272203|T191|LLT|10056452|MDR|Indolent systemic mastocytosis|9741/1
C0272203|T191|SY|352954|MEDCIN|anomalies of skin mastocytosis indolent systemic|9741/1
C0272203|T191|PT|352954|MEDCIN|Indolent systemic mastocytosis|9741/1
C0272203|T191|PM|D034721|MSH|Indolent Systemic Mastocytoses|9741/1
C0272203|T191|PEP|D034721|MSH|Indolent Systemic Mastocytosis|9741/1
C0272203|T191|PM|D034721|MSH|Mastocytoses, Indolent Systemic|9741/1
C0272203|T191|PM|D034721|MSH|Mastocytosis, Indolent Systemic|9741/1
C0272203|T191|PM|D034721|MSH|Systemic Mastocytoses, Indolent|9741/1
C0272203|T191|PM|D034721|MSH|Systemic Mastocytosis, Indolent|9741/1
C0272203|T191|PN|NOCODE|MTH|Indolent Systemic Mastocytosis|9741/1
C0272203|T191|SY|TCGA|NCI|Indolent Systemic Mastocytosis|9741/1
C0272203|T191|PT|C9286|NCI|Indolent Systemic Mastocytosis|9741/1
C0272203|T191|AB|C9286|NCI|ISM|9741/1
C0272203|T191|DN|C9286|NCI_CTRP|Indolent Systemic Mastocytosis|9741/1
C0272203|T191|PT|CDR0000613597|PDQ|indolent systemic mastocytosis|9741/1
C0272203|T191|AB|CDR0000613597|PDQ|ISM|9741/1
C0272203|T191|PT|70910003|SNOMEDCT_US|Indolent systemic mastocytosis|9741/1
C0272203|T191|PT|397356009|SNOMEDCT_US|Indolent systemic mastocytosis|9741/1
C1112486|T191|AB|C96.21|ICD10CM|Aggressive systemic mastocytosis|9741/3
C1112486|T191|PT|C96.21|ICD10CM|Aggressive systemic mastocytosis|9741/3
C1541840|T191|PT|MTHU047300|ICPC2ICD10ENG|malignant; mastocytosis|9741/3
C1541840|T191|PT|MTHU047647|ICPC2ICD10ENG|mastocytosis; malignant|9741/3
C1112486|T191|LLT|10056453|MDR|Aggressive systemic mastocytosis|9741/3
C1112486|T191|PT|365413|MEDCIN|Aggressive systemic mastocytosis|9741/3
C1112486|T191|PT|356718|MEDCIN|agressive lymphadenopathic mastocytosis with eosinophilia|9741/3
C1112486|T191|SY|365413|MEDCIN|malignant mast cell tumor aggressive systemic mastocytosis|9741/3
C1541840|T191|PT|31762|MEDCIN|malignant mastocytosis|9741/3
C1541840|T191|PT|272064|MEDCIN|malignant mastocytosis of reticuloendothelial system|9741/3
C1301365|T191|SY|356719|MEDCIN|systemic mastocytosis w/ assoc clonal hematologic non-mast cell lineage disease|9741/3
C1301365|T191|PT|356719|MEDCIN|systemic mastocytosis with associated clonal hematologic non-mast cell lineage disease|9741/3
C1112486|T191|PM|D034721|MSH|Aggressive Systemic Mastocytoses|9741/3
C1112486|T191|PEP|D034721|MSH|Aggressive Systemic Mastocytosis|9741/3
C1112486|T191|PM|D034721|MSH|Mastocytoses, Aggressive Systemic|9741/3
C1112486|T191|PM|D034721|MSH|Mastocytosis, Aggressive Systemic|9741/3
C1112486|T191|PM|D034721|MSH|Systemic Mastocytoses, Aggressive|9741/3
C1112486|T191|PM|D034721|MSH|Systemic Mastocytosis, Aggressive|9741/3
C1112486|T191|PN|NOCODE|MTH|Aggressive Systemic Mastocytosis|9741/3
C1541840|T191|PN|NOCODE|MTH|Malignant mastocytosis|9741/3
C1541840|T191|ET|202.6|MTHICD9|Malignant mastocytosis|9741/3
C1112486|T191|SY|TCGA|NCI|Aggressive Systemic Mastocytosis|9741/3
C1112486|T191|PT|C9285|NCI|Aggressive Systemic Mastocytosis|9741/3
C1112486|T191|AB|C9285|NCI|ASM|9741/3
C1541840|T191|PT|C8991|NCI|Malignant Mastocytosis|9741/3
C1301365|T191|AB|C9284|NCI|SM-AHN|9741/3
C1301365|T191|AB|C9284|NCI|SM-AHNMD|9741/3
C1301365|T191|PT|C9284|NCI|Systemic Mastocytosis with an Associated Hematological Neoplasm|9741/3
C1301365|T191|SY|C9284|NCI|Systemic Mastocytosis with Associated Clonal Hematological non-Mast-Cell Lineage Disease|9741/3
C1541840|T191|PT|C8991|NCI_CDISC|MAST CELL TUMOR, MALIGNANT|9741/3
C1541840|T191|PT|C8991|NCI_CPTAC|Malignant Mastocytosis|9741/3
C1112486|T191|DN|C9285|NCI_CTRP|Aggressive Systemic Mastocytosis|9741/3
C1112486|T191|PT|CDR0000613596|PDQ|aggressive systemic mastocytosis|9741/3
C1112486|T191|AB|CDR0000613596|PDQ|ASM|9741/3
C1301365|T191|AB|CDR0000778560|PDQ|SM-AHN|9741/3
C1301365|T191|AB|CDR0000778560|PDQ|SM-AHNMD|9741/3
C1301365|T191|PT|CDR0000778560|PDQ|systemic mastocytosis with an associated hematological neoplasm|9741/3
C1301365|T191|SY|CDR0000778560|PDQ|systemic mastocytosis with associated clonal hematological non-mast-cell lineage disease|9741/3
C1541840|T191|PT|XaBAk|RCD|Malignant mastocytosis|9741/3
C1541840|T191|PT|BBp2.|RCDSY|Malignant mastocytosis|9741/3
C1112486|T191|PT|397008008|SNOMEDCT_US|Aggressive lymphadenopathic mastocytosis with eosinophilia|9741/3
C1112486|T191|PT|716655008|SNOMEDCT_US|Aggressive systemic mastocytosis|9741/3
C1112486|T191|IS|397008008|SNOMEDCT_US|Aggressive systemic mastocytosis|9741/3
C1112486|T191|PT|397358005|SNOMEDCT_US|Aggressive systemic mastocytosis|9741/3
C1112486|T191|SY|397008008|SNOMEDCT_US|Lymphadenopathic mastocytosis with eosinophilia|9741/3
C1541840|T191|PT|50150000|SNOMEDCT_US|Malignant mastocytosis|9741/3
C1541840|T191|OAP|307591004|SNOMEDCT_US|Malignant mastocytosis|9741/3
C1541840|T191|OAP|123311009|SNOMEDCT_US|Malignant mastocytosis|9741/3
C1541840|T191|IS|123311009|SNOMEDCT_US|Malignant mastocytosis -RETIRED-|9741/3
C1541840|T191|OF|123311009|SNOMEDCT_US|Malignant mastocytosis -RETIRED-|9741/3
C1301365|T191|SY|397357000|SNOMEDCT_US|Systemic mastocytosis with AHNMD|9741/3
C1301365|T191|PTGB|397015000|SNOMEDCT_US|Systemic mastocytosis with associated clonal haematological non-mast cell lineage disease|9741/3
C1301365|T191|PT|397015000|SNOMEDCT_US|Systemic mastocytosis with associated clonal hematological non-mast cell lineage disease|9741/3
C1301365|T191|PTGB|397357000|SNOMEDCT_US|Systemic mastocytosis with associated clonal, haematologic non-mast-cell lineage disease|9741/3
C1301365|T191|PT|397357000|SNOMEDCT_US|Systemic mastocytosis with associated clonal, hematologic non-mast-cell lineage disease|9741/3
C1301365|T191|SYGB|397357000|SNOMEDCT_US|Systemic mastocytosis with associated haematological clonal non-mast cell disorder|9741/3
C1301365|T191|SY|397357000|SNOMEDCT_US|Systemic mastocytosis with associated hematological clonal non-mast cell disorder|9741/3
C0023461|T191|SY|0000007340|CHV|mast cell leukaemia|9742/3
C0023461|T191|PT|0000007340|CHV|mast cell leukemia|9742/3
C0023461|T191|PT|C94.3|ICD10|Mast cell leukaemia|9742/3
C0023461|T191|PT|C94.3|ICD10AE|Mast cell leukemia|9742/3
C0023461|T191|AB|C94.3|ICD10CM|Mast cell leukemia|9742/3
C0023461|T191|HT|C94.3|ICD10CM|Mast cell leukemia|9742/3
C0023461|T191|ET|C94.30|ICD10CM|Mast cell leukemia NOS|9742/3
C0023461|T191|PT|MTHU044771|ICPC2ICD10ENG|leukemia; mast cell|9742/3
C0023461|T191|PT|MTHU048975|ICPC2ICD10ENG|mast cell; leukemia|9742/3
C0023461|T191|PT|10056450|MDR|Mastocytic leukaemia|9742/3
C0023461|T191|LLT|10056450|MDR|Mastocytic leukaemia|9742/3
C0023461|T191|LLT|10056451|MDR|Mastocytic leukemia|9742/3
C0023461|T191|MTH_PT|10056450|MDR|Mastocytic leukemia|9742/3
C0023461|T191|PT|31471|MEDCIN|mast cell leukemia|9742/3
C0023461|T191|PM|D007946|MSH|Leukemia, Mast Cell|9742/3
C0023461|T191|MH|D007946|MSH|Leukemia, Mast-Cell|9742/3
C0023461|T191|PM|D007946|MSH|Leukemias, Mast-Cell|9742/3
C0023461|T191|PM|D007946|MSH|Mast Cell Leukemia|9742/3
C0023461|T191|ET|D007946|MSH|Mast-Cell Leukemia|9742/3
C0023461|T191|PM|D007946|MSH|Mast-Cell Leukemias|9742/3
C0023461|T191|PN|NOCODE|MTH|Leukemia, Mast-Cell|9742/3
C0023461|T191|PT|C3169|NCI|Mast Cell Leukemia|9742/3
C0023461|T191|SY|TCGA|NCI|Mast Cell Leukemia|9742/3
C0023461|T191|PT|C3169|NCI_CPTAC|Mast Cell Leukemia|9742/3
C0023461|T191|DN|C3169|NCI_CTRP|Mast Cell Leukemia|9742/3
C0023461|T191|PT|CDR0000466588|PDQ|mast cell leukemia|9742/3
C0023461|T191|AB|CDR0000466588|PDQ|MCL|9742/3
C0023461|T191|OP|B673.|RCD|Mast cell leukaemia|9742/3
C0023461|T191|OP|B673.|RCDAE|Mast cell leukemia|9742/3
C0023461|T191|PT|BBrA0|RCDSA|Mast cell leukemia|9742/3
C0023461|T191|PT|BBrA0|RCDSY|Mast cell leukaemia|9742/3
C0023461|T191|OAP|188755006|SNOMEDCT_US|Mast cell leukaemia|9742/3
C0023461|T191|PTGB|128924002|SNOMEDCT_US|Mast cell leukaemia|9742/3
C0023461|T191|SYGB|110002002|SNOMEDCT_US|Mast cell leukaemia|9742/3
C0023461|T191|OAP|70798001|SNOMEDCT_US|Mast cell leukaemia|9742/3
C0023461|T191|IS|70798001|SNOMEDCT_US|Mast cell leukaemia -RETIRED-|9742/3
C0023461|T191|SY|110002002|SNOMEDCT_US|Mast cell leukemia|9742/3
C0023461|T191|OAP|188755006|SNOMEDCT_US|Mast cell leukemia|9742/3
C0023461|T191|PT|128924002|SNOMEDCT_US|Mast cell leukemia|9742/3
C0023461|T191|OAP|70798001|SNOMEDCT_US|Mast cell leukemia|9742/3
C0023461|T191|IS|70798001|SNOMEDCT_US|Mast cell leukemia -RETIRED-|9742/3
C0023461|T191|OF|70798001|SNOMEDCT_US|Mast cell leukemia -RETIRED-|9742/3
C0023461|T191|IS|70798001|SNOMEDCT_US|Noncutaneous systemic mastocytosis|9742/3
C0878675|T047|SY|0000051996|CHV|chester disease erdheim|9750/1
C0878675|T047|PT|0000051996|CHV|erdheim chester disease|9750/1
C0878675|T047|SY|0000051996|CHV|erdheim-chester disease|9750/1
C0878675|T047|PT|29792|DDB|Erdheim-Chester disease|9750/1
C0878675|T047|PT|10060801|MDR|Erdheim-Chester disease|9750/1
C0878675|T047|LLT|10060801|MDR|Erdheim-Chester disease|9750/1
C0878675|T047|SY|313968|MEDCIN|Erdheim-Chester syndrome|9750/1
C0878675|T047|PT|313968|MEDCIN|polyostotic sclerosing histiocytosis|9750/1
C0878675|T047|PM|D031249|MSH|Erdheim Chester Disease|9750/1
C0878675|T047|MH|D031249|MSH|Erdheim-Chester Disease|9750/1
C0878675|T047|ET|D031249|MSH|Granulomatosis, Lipid|9750/1
C0878675|T047|PM|D031249|MSH|Lipid Granulomatosis|9750/1
C0878675|T047|PN|NOCODE|MTH|Erdheim-Chester Disease|9750/1
C0878675|T047|PT|C53972|NCI|Erdheim-Chester Disease|9750/1
C0878675|T047|SY|C53972|NCI|Lipogranulomatosis|9750/1
C0878675|T047|SY|C53972|NCI|Polyostotic Sclerosing Histiocytosis|9750/1
C0878675|T047|PT|CDR0000710367|PDQ|Erdheim-Chester disease|9750/1
C0878675|T047|SY|CDR0000710367|PDQ|lipogranulomatosis|9750/1
C0878675|T047|SY|CDR0000710367|PDQ|polyostotic sclerosing histiocytosis|9750/1
C0878675|T047|SY|699537002|SNOMEDCT_US|Erdheim-Chester disease|9750/1
C0878675|T047|OAP|703711007|SNOMEDCT_US|Erdheim-Chester disease|9750/1
C0878675|T047|SY|699537002|SNOMEDCT_US|Erdheim-Chester syndrome|9750/1
C0878675|T047|PT|699537002|SNOMEDCT_US|Polyostotic sclerosing histiocytosis|9750/1
C0019623|T191|SY|0000006166|CHV|angiocentric lymphoma|9750/3
C0019623|T191|SY|0000006166|CHV|angiocentric t-cell lymphoma|9750/3
C0019623|T191|SY|0000006166|CHV|histiocytic medullary reticulosis|9750/3
C0019623|T191|SY|0000006166|CHV|histiocytosis malignant|9750/3
C0019623|T191|SY|0000006166|CHV|lymphoma nasal t-cell|9750/3
C0019623|T191|PT|0000006166|CHV|malignant histiocytosis|9750/3
C0019623|T191|SY|0000006166|CHV|nasal t-cell lymphoma|9750/3
C0019623|T191|SY|0000006166|CHV|polymorphic reticulosis|9750/3
C0019623|T191|SY|0000006166|CHV|stewart's granuloma|9750/3
C0019623|T191|DI|U000848|DXP|HISTIOCYTOSIS, MALIGNANT|9750/3
C0019623|T191|SY|NOCODE|DXP|RETICULOSIS, ALEUKEMIC|9750/3
C0019623|T191|SY|NOCODE|DXP|RETICULOSIS, MALIGNANT|9750/3
C0019623|T191|SY|NOCODE|DXP|RETICULOSIS, MALIGNANT MIDLINE|9750/3
C0019623|T191|SY|NOCODE|DXP|RETICULOSIS, POLYMORPHORIC|9750/3
C0019623|T191|PT|C96.1|ICD10|Malignant histiocytosis|9750/3
C0019623|T191|ET|C96.A|ICD10CM|Malignant histiocytosis|9750/3
C0019623|T191|HT|202.3|ICD9CM|Malignant histiocytosis|9750/3
C0019623|T191|PT|MTHU035175|ICPC2ICD10ENG|histiocytosis; malignant|9750/3
C0019623|T191|PT|MTHU047290|ICPC2ICD10ENG|malignant; histiocytosis|9750/3
C0019623|T191|PT|MTHU047309|ICPC2ICD10ENG|malignant; reticuloendotheliosis|9750/3
C0019623|T191|PT|MTHU047310|ICPC2ICD10ENG|malignant; reticulosis|9750/3
C0019623|T191|PT|MTHU060950|ICPC2ICD10ENG|polymorphic; reticulosis|9750/3
C0019623|T191|PT|MTHU064352|ICPC2ICD10ENG|reticuloendotheliosis; malignant|9750/3
C0019623|T191|PT|MTHU064369|ICPC2ICD10ENG|reticulosis; malignant|9750/3
C0019623|T191|PT|MTHU064371|ICPC2ICD10ENG|reticulosis; polymorphic|9750/3
C0019623|T191|LLT|10025581|MDR|Malignant histiocytosis|9750/3
C0019623|T191|PT|10025581|MDR|Malignant histiocytosis|9750/3
C0019623|T191|LLT|10027591|MDR|Midline malignant reticulosis|9750/3
C0019623|T191|LLT|10028772|MDR|Nasal T-cell lymphoma|9750/3
C0019623|T191|LLT|10036088|MDR|Polymorphic reticulosis|9750/3
C0019623|T191|PT|272065|MEDCIN|malignant histiocytosis|9750/3
C0019623|T191|PM|D054747|MSH|Histiocytoses, Malignant|9750/3
C0019623|T191|PEP|D054747|MSH|Histiocytosis, Malignant|9750/3
C0019623|T191|PM|D054747|MSH|Malignant Histiocytoses|9750/3
C0019623|T191|ET|D054747|MSH|Malignant Histiocytosis|9750/3
C0019623|T191|PN|NOCODE|MTH|Malignant histiocytosis|9750/3
C0019623|T191|ET|202.3|MTHICD9|Malignant reticuloendotheliosis|9750/3
C0019623|T191|ET|202.3|MTHICD9|Malignant reticulosis|9750/3
C0019623|T191|OP|C7202|NCI|Histiocytic Medullary Reticulosis|9750/3
C0019623|T191|OP|C7202|NCI|Malignant Histiocytosis|9750/3
C0019623|T191|PT|C7202|NCI|Malignant Histiocytosis|9750/3
C0019623|T191|PT|B623.|RCD|Malignant histiocytosis|9750/3
C0019623|T191|OP|B623z|RCD|Malignant histiocytosis NOS|9750/3
C0019623|T191|SY|G753.|RCD|Malignant midline reticulosis|9750/3
C0019623|T191|AB|Xa0To|RCD|Malignant reticuloendothelios|9750/3
C0019623|T191|SY|Xa0To|RCD|Malignant reticuloendotheliosis|9750/3
C0019623|T191|SY|B623.|RCD|Malignant reticulosis|9750/3
C0019623|T191|SY|Xa0To|RCD|Malignant reticulosis|9750/3
C0019623|T191|SY|Xa0To|RCD|Polymorphic reticulosis|9750/3
C0019623|T191|SY|Xa0To|RCD|Stewart's granuloma|9750/3
C0019623|T191|OP|BBm1.|RCDSY|Malignant histiocytosis|9750/3
C0019623|T191|IS|BBm1.|RCDSY|Malignant reticulosis|9750/3
C0019623|T191|SY|118612006|SNOMEDCT_US|Malignant histiocytosis|9750/3
C0019623|T191|OAP|8139000|SNOMEDCT_US|Malignant histiocytosis|9750/3
C0019623|T191|OAP|188690006|SNOMEDCT_US|Malignant histiocytosis|9750/3
C0019623|T191|PT|128920006|SNOMEDCT_US|Malignant histiocytosis|9750/3
C0019623|T191|OF|188690006|SNOMEDCT_US|Malignant histiocytosis|9750/3
C0019623|T191|IS|8139000|SNOMEDCT_US|Malignant histiocytosis -RETIRED-|9750/3
C0019623|T191|OF|8139000|SNOMEDCT_US|Malignant histiocytosis -RETIRED-|9750/3
C0019623|T191|OAP|188643009|SNOMEDCT_US|Malignant histiocytosis NOS|9750/3
C0019623|T191|IS|66855003|SNOMEDCT_US|Malignant midline reticulosis|9750/3
C0019623|T191|OAS|277648007|SNOMEDCT_US|Malignant reticuloendotheliosis|9750/3
C0019623|T191|SY|118612006|SNOMEDCT_US|Malignant reticulosis|9750/3
C0019623|T191|OAS|277648007|SNOMEDCT_US|Malignant reticulosis|9750/3
C0019623|T191|IS|66855003|SNOMEDCT_US|Malignant reticulosis, NOS|9750/3
C0019623|T191|IS|66855003|SNOMEDCT_US|Polymorphic reticulosis|9750/3
C0019623|T191|OAS|277648007|SNOMEDCT_US|Polymorphic reticulosis|9750/3
C0019623|T191|OAS|277648007|SNOMEDCT_US|Stewart's granuloma|9750/3
C0019621|T191|SY|0000006165|CHV|cell granulomatosis langerhans|9751/1
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhan|9751/1
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhans|9751/1
C0019621|T191|SY|0000006165|CHV|cells histiocytosis langerhans|9751/1
C0019621|T191|SY|0000026274|CHV|christian disease hand schuller|9751/1
C0019621|T191|SY|0000026274|CHV|christian diseases hand schuller|9751/1
C0019621|T191|SY|0000026274|CHV|disease hand schuller christian|9751/1
C0019621|T191|SY|0000007324|CHV|generalized histiocytosis|9751/1
C0019621|T191|SY|0000026274|CHV|hand christian schuller disease|9751/1
C0019621|T191|SY|0000026274|CHV|hand schuller christian disease|9751/1
C0019621|T191|SY|0000026274|CHV|hand-schueller-christian disease|9751/1
C0019621|T191|PT|0000026274|CHV|hand-schuller-christian disease|9751/1
C0019621|T191|PT|0000006165|CHV|histiocytosis x|9751/1
C0019621|T191|SY|0000006165|CHV|histiocytosis-x|9751/1
C0019621|T191|SY|0000006165|CHV|langerhan's cell histiocytosis|9751/1
C0019621|T191|SY|0000006165|CHV|langerhans cell disease|9751/1
C0019621|T191|SY|0000006165|CHV|langerhans cell granulomatosis|9751/1
C0019621|T191|SY|0000006165|CHV|langerhans cell histiocytosis|9751/1
C0019621|T191|SY|0000026274|CHV|schuller christian syndrome|9751/1
C0019621|T191|ET|0427-5330|CSP|Hand Schuller Christian disease|9751/1
C0019621|T191|PT|0427-5330|CSP|histiocytosis X|9751/1
C0019621|T191|ET|0427-5330|CSP|Langerhans cell granulomatosis|9751/1
C0019621|T191|SY|NOCODE|DXP|EOSINOPHILIC GRANULOMA, MULTIFOCAL|9751/1
C0019621|T191|DI|U000766|DXP|HAND-SCHUELLER-CHRISTIAN SYNDROME|9751/1
C0019621|T191|SY|NOCODE|DXP|HISTIOCYTOSIS X II|9751/1
C0019621|T191|SY|NOCODE|DXP|SCHUELLER-CHRISTIAN DISEASE|9751/1
C0019621|T191|ET|C96.5|ICD10CM|Hand-Schüller-Christian disease|9751/1
C0019621|T191|ET|C96.6|ICD10CM|Langerhans-cell histiocytosis NOS|9751/1
C0019621|T191|PT|MTHU033317|ICPC2ICD10ENG|Hand-Schüller-Christian|9751/1
C0019621|T191|PT|MTHU035172|ICPC2ICD10ENG|histiocytosis; Langerhans' cell|9751/1
C0019621|T191|PT|MTHU035180|ICPC2ICD10ENG|histiocytosis; X|9751/1
C0019621|T191|PT|MTHU035182|ICPC2ICD10ENG|histiocytosis; X, chronic|9751/1
C0019621|T191|PT|MTHU042862|ICPC2ICD10ENG|Langerhans' cell; histiocytosis|9751/1
C0019621|T191|PT|MTHU066496|ICPC2ICD10ENG|Schüller-Christian|9751/1
C0019621|T191|PT|MTHU082788|ICPC2ICD10ENG|X; histiocytosis|9751/1
C0019621|T191|PT|MTHU082790|ICPC2ICD10ENG|X; histiocytosis, chronic|9751/1
C0019621|T191|PT|U002076|LCH|Hand-Schueller-Christian syndrome|9751/1
C0019621|T191|PT|sh85058638|LCH_NW|Hand-Schueller-Christian syndrome|9751/1
C0019621|T191|LLT|10053133|MDR|Chronic idiopathic xanthomatosis|9751/1
C0019621|T191|LLT|10053135|MDR|Hand-Schueller-Christian disease|9751/1
C0019621|T191|LLT|10023688|MDR|Langerhans' cell granulomatosis|9751/1
C0019621|T191|LLT|10069698|MDR|Langerhans' cell histiocytosis|9751/1
C0019621|T191|PT|10069698|MDR|Langerhans' cell histiocytosis|9751/1
C0019621|T191|SY|31815|MEDCIN|Hand-Schuller-Christian disease|9751/1
C0019621|T191|PT|315032|MEDCIN|Langerhans cell histiocytosis|9751/1
C0019621|T191|PT|31815|MEDCIN|multifocal eosinophilic granuloma|9751/1
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendothelioses, Systemic|9751/1
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendotheliosis, Systemic|9751/1
C0019621|T191|PM|D006646|MSH|Cell Granulomatoses, Langerhans|9751/1
C0019621|T191|PM|D006646|MSH|Cell Granulomatosis, Langerhans|9751/1
C0019621|T191|PM|D006646|MSH|Cell Histiocytoses, Langerhans|9751/1
C0019621|T191|PM|D006646|MSH|Cell Histiocytosis, Langerhans|9751/1
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schueller-Christian|9751/1
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schüller-Christian|9751/1
C0019621|T191|PM|D006646|MSH|Disease, Letterer-Siwe|9751/1
C0019621|T191|PM|D006646|MSH|Disease, Schueller-Christian|9751/1
C0019621|T191|PM|D006646|MSH|Generalized Histiocytoses|9751/1
C0019621|T191|PM|D006646|MSH|Generalized Histiocytosis|9751/1
C0019621|T191|PM|D006646|MSH|Granulomatoses, Langerhans Cell|9751/1
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans Cell|9751/1
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans-Cell|9751/1
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Disease|9751/1
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Syndrome|9751/1
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Disease|9751/1
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Syndrome|9751/1
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Disease|9751/1
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Syndrome|9751/1
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Disease|9751/1
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Syndrome|9751/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Generalized|9751/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Langerhans Cell|9751/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Type 2|9751/1
C0019621|T191|ET|D006646|MSH|Histiocytosis X|9751/1
C0019621|T191|ET|D006646|MSH|Histiocytosis-X|9751/1
C0019621|T191|ET|D006646|MSH|Histiocytosis, Generalized|9751/1
C0019621|T191|PM|D006646|MSH|Histiocytosis, Langerhans Cell|9751/1
C0019621|T191|MH|D006646|MSH|Histiocytosis, Langerhans-Cell|9751/1
C0019621|T191|PM|D006646|MSH|Histiocytosis, Type 2|9751/1
C0019621|T191|PM|D006646|MSH|Langerhans Cell Granulomatoses|9751/1
C0019621|T191|ET|D006646|MSH|Langerhans Cell Granulomatosis|9751/1
C0019621|T191|PM|D006646|MSH|Langerhans Cell Histiocytoses|9751/1
C0019621|T191|ET|D006646|MSH|Langerhans Cell Histiocytosis|9751/1
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Granulomatosis|9751/1
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Histiocytosis|9751/1
C0019621|T191|DEV|D006646|MSH|LETTERER SIWE DIS|9751/1
C0019621|T191|PM|D006646|MSH|Letterer Siwe Disease|9751/1
C0019621|T191|ET|D006646|MSH|Letterer-Siwe Disease|9751/1
C0019621|T191|PM|D006646|MSH|Non Lipid Reticuloendotheliosis|9751/1
C0019621|T191|PM|D006646|MSH|Non-Lipid Reticuloendothelioses|9751/1
C0019621|T191|ET|D006646|MSH|Non-Lipid Reticuloendotheliosis|9751/1
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Non-Lipid|9751/1
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Systemic Aleukemic|9751/1
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Non-Lipid|9751/1
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Systemic Aleukemic|9751/1
C0019621|T191|DEV|D006646|MSH|SCHUELLER CHRISTIAN DIS|9751/1
C0019621|T191|PM|D006646|MSH|Schueller Christian Disease|9751/1
C0019621|T191|ET|D006646|MSH|Schueller-Christian Disease|9751/1
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schueller-Christian|9751/1
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schüller-Christian|9751/1
C0019621|T191|PM|D006646|MSH|Systemic Aleukemic Reticuloendothelioses|9751/1
C0019621|T191|ET|D006646|MSH|Systemic Aleukemic Reticuloendotheliosis|9751/1
C0019621|T191|PM|D006646|MSH|Type 2 Histiocytoses|9751/1
C0019621|T191|ET|D006646|MSH|Type 2 Histiocytosis|9751/1
C0019621|T191|PN|NOCODE|MTH|Histiocytosis, Langerhans-Cell|9751/1
C0019621|T191|ET|277.89|MTHICD9|Chronic Histiocytosis X|9751/1
C0019621|T191|ET|277.89|MTHICD9|Hand-Schuller-Christian disease|9751/1
C0019621|T191|ET|277.89|MTHICD9|Histiocytosis X|9751/1
C0019621|T191|PT|C6920|NCI|Hand-Schuller-Christian Disease|9751/1
C0019621|T191|OP|C3107|NCI|Histiocytosis X|9751/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Granulomatosis|9751/1
C0019621|T191|PT|C3107|NCI|Langerhans Cell Histiocytosis|9751/1
C0019621|T191|SY|TCGA|NCI|Langerhans Cell Histiocytosis|9751/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, NOS|9751/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, Not Otherwise Specified|9751/1
C0019621|T191|AB|C3107|NCI|LCH|9751/1
C0019621|T191|PT|C6920|NCI_CPTAC|Hand-Schuller-Christian Disease|9751/1
C0019621|T191|PT|10025581|NCI_CTEP-SDC|Langerhans cell histiocytosis|9751/1
C0019621|T191|DN|C3107|NCI_CTRP|Langerhans Cell Histiocytosis|9751/1
C0019621|T191|PT|CDR0000471787|NCI_NCI-GLOSS|Langerhans cell histiocytosis|9751/1
C0019621|T191|PT|CDR0000513054|NCI_NCI-GLOSS|LCH|9751/1
C0019621|T191|SY|C6920|NCI_NICHD|Classic Multifocal Langerhans Cell Histiocytosis|9751/1
C0019621|T191|SY|C6920|NCI_NICHD|Hand-Schüller-Christian Disease|9751/1
C0019621|T191|OP|C3107|NCI_NICHD|Histiocytosis X|9751/1
C0019621|T191|PT|C3107|NCI_NICHD|Langerhans Cell Histiocytosis|9751/1
C0019621|T191|PT|C6920|NCI_NICHD|Multifocal Unisystem Langerhans Cell Histiocytosis|9751/1
C0019621|T191|SY|CDR0000039054|PDQ|histiocytosis X|9751/1
C0019621|T191|PT|CDR0000641624|PDQ|Langerhans cell histiocytosis|9751/1
C0019621|T191|AB|X20E9|RCD|Different progress histiocyto|9751/1
C0019621|T191|SY|X20E9|RCD|Differentiated progressive histiocytosis|9751/1
C0019621|T191|AB|C37y0|RCD|Hand-Schuller-Christian diseas|9751/1
C0019621|T191|SY|C37y0|RCD|Hand-Schuller-Christian disease|9751/1
C0019621|T191|OP|C37y6|RCD|Histiocytosis X , unspecified|9751/1
C0019621|T191|PT|C37y5|RCD|Histiocytosis X syndrome|9751/1
C0019621|T191|PT|X20E9|RCD|Langerhan's cell histiocytosis|9751/1
C0019621|T191|AB|X20E9|RCD|Langerhans histiocyt syndrome|9751/1
C0019621|T191|SY|X20E9|RCD|Langerhans histiocytic syndrome|9751/1
C0019621|T191|SY|X20E9|RCD|LCH - Langerhan's cell histiocytosis|9751/1
C0019621|T191|AB|X20E9|RCD|LCH-Langerh cell histiocytosis|9751/1
C0019621|T191|PT|C37y0|RCD|Schuller-Christian syndrome|9751/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic differentiated progressive histiocytosis|9751/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic disseminated histiocytosis X|9751/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic histiocytosis X|9751/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic idiopathic xanthomatosis|9751/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Differentiated progressive histiocytosis|9751/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Differentiated progressive histiocytosis|9751/1
C0019621|T191|SYGB|39795003|SNOMEDCT_US|Generalised histiocytosis of bones|9751/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Generalized histiocytosis of bones|9751/1
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand - Schuller - Christian disease|9751/1
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand - Schuller - Christian disease|9751/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Hand-Schuller-Christian disease|9751/1
C0019621|T191|PT|39795003|SNOMEDCT_US|Hand-Schüller-Christian disease|9751/1
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9751/1
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9751/1
C0019621|T191|OAS|154583006|SNOMEDCT_US|Histiocytosis X|9751/1
C0019621|T191|OAS|269628007|SNOMEDCT_US|Histiocytosis X|9751/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Histiocytosis X|9751/1
C0019621|T191|IS|190960001|SNOMEDCT_US|Histiocytosis X , chronic|9751/1
C0019621|T191|IS|190956004|SNOMEDCT_US|Histiocytosis X , unspecified|9751/1
C0019621|T191|PT|190955000|SNOMEDCT_US|Histiocytosis X syndrome|9751/1
C0019621|T191|IS|65399007|SNOMEDCT_US|Histiocytosis X, NOS|9751/1
C0019621|T191|OAP|190956004|SNOMEDCT_US|Histiocytosis X, unspecified|9751/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhan's cell histiocytosis|9751/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhan's cell histiocytosis|9751/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans cell disease|9751/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhans cell disease|9751/1
C0019621|T191|IS|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9751/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9751/1
C0019621|T191|OAP|234439008|SNOMEDCT_US|Langerhans cell histiocytosis|9751/1
C0019621|T191|PT|65399007|SNOMEDCT_US|Langerhans cell histiocytosis|9751/1
C0019621|T191|PT|128809007|SNOMEDCT_US|Langerhans cell histiocytosis|9751/1
C0019621|T191|PT|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, multifocal|9751/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no ICD-O subtype|9751/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no International Classification of Diseases for Oncology subtype|9751/1
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, poly-ostotic|9751/1
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, polyostotic|9751/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans histiocytic syndrome|9751/1
C0019621|T191|OAP|110450007|SNOMEDCT_US|Langerhans' cell histiocytosis|9751/1
C0019621|T191|SY|65399007|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9751/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9751/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Multifocal and unisystemic Langerhans cell histiocytosis|9751/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Schuller-Christian syndrome|9751/1
C0019621|T191|SY|0000006165|CHV|cell granulomatosis langerhans|9751/3
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhan|9751/3
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhans|9751/3
C0019621|T191|SY|0000006165|CHV|cells histiocytosis langerhans|9751/3
C0019621|T191|SY|0000026274|CHV|christian disease hand schuller|9751/3
C0019621|T191|SY|0000026274|CHV|christian diseases hand schuller|9751/3
C0019621|T191|SY|0000026274|CHV|disease hand schuller christian|9751/3
C0019621|T191|SY|0000007324|CHV|generalized histiocytosis|9751/3
C0019621|T191|SY|0000026274|CHV|hand christian schuller disease|9751/3
C0019621|T191|SY|0000026274|CHV|hand schuller christian disease|9751/3
C0019621|T191|SY|0000026274|CHV|hand-schueller-christian disease|9751/3
C0019621|T191|PT|0000026274|CHV|hand-schuller-christian disease|9751/3
C0019621|T191|PT|0000006165|CHV|histiocytosis x|9751/3
C0019621|T191|SY|0000006165|CHV|histiocytosis-x|9751/3
C0019621|T191|SY|0000006165|CHV|langerhan's cell histiocytosis|9751/3
C0019621|T191|SY|0000006165|CHV|langerhans cell disease|9751/3
C0019621|T191|SY|0000006165|CHV|langerhans cell granulomatosis|9751/3
C0019621|T191|SY|0000006165|CHV|langerhans cell histiocytosis|9751/3
C0019621|T191|SY|0000026274|CHV|schuller christian syndrome|9751/3
C0019621|T191|ET|0427-5330|CSP|Hand Schuller Christian disease|9751/3
C0019621|T191|PT|0427-5330|CSP|histiocytosis X|9751/3
C0019621|T191|ET|0427-5330|CSP|Langerhans cell granulomatosis|9751/3
C0019621|T191|SY|NOCODE|DXP|EOSINOPHILIC GRANULOMA, MULTIFOCAL|9751/3
C0019621|T191|DI|U000766|DXP|HAND-SCHUELLER-CHRISTIAN SYNDROME|9751/3
C0019621|T191|SY|NOCODE|DXP|HISTIOCYTOSIS X II|9751/3
C0019621|T191|SY|NOCODE|DXP|SCHUELLER-CHRISTIAN DISEASE|9751/3
C0019621|T191|ET|C96.5|ICD10CM|Hand-Schüller-Christian disease|9751/3
C0019621|T191|ET|C96.6|ICD10CM|Langerhans-cell histiocytosis NOS|9751/3
C0019621|T191|PT|MTHU033317|ICPC2ICD10ENG|Hand-Schüller-Christian|9751/3
C0019621|T191|PT|MTHU035172|ICPC2ICD10ENG|histiocytosis; Langerhans' cell|9751/3
C0019621|T191|PT|MTHU035180|ICPC2ICD10ENG|histiocytosis; X|9751/3
C0019621|T191|PT|MTHU035182|ICPC2ICD10ENG|histiocytosis; X, chronic|9751/3
C0019621|T191|PT|MTHU042862|ICPC2ICD10ENG|Langerhans' cell; histiocytosis|9751/3
C0019621|T191|PT|MTHU066496|ICPC2ICD10ENG|Schüller-Christian|9751/3
C0019621|T191|PT|MTHU082788|ICPC2ICD10ENG|X; histiocytosis|9751/3
C0019621|T191|PT|MTHU082790|ICPC2ICD10ENG|X; histiocytosis, chronic|9751/3
C0019621|T191|PT|U002076|LCH|Hand-Schueller-Christian syndrome|9751/3
C0019621|T191|PT|sh85058638|LCH_NW|Hand-Schueller-Christian syndrome|9751/3
C0019621|T191|LLT|10053133|MDR|Chronic idiopathic xanthomatosis|9751/3
C0019621|T191|LLT|10053135|MDR|Hand-Schueller-Christian disease|9751/3
C0019621|T191|LLT|10023688|MDR|Langerhans' cell granulomatosis|9751/3
C0019621|T191|LLT|10069698|MDR|Langerhans' cell histiocytosis|9751/3
C0019621|T191|PT|10069698|MDR|Langerhans' cell histiocytosis|9751/3
C0019621|T191|SY|31815|MEDCIN|Hand-Schuller-Christian disease|9751/3
C0019621|T191|PT|315032|MEDCIN|Langerhans cell histiocytosis|9751/3
C0019621|T191|PT|31815|MEDCIN|multifocal eosinophilic granuloma|9751/3
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendothelioses, Systemic|9751/3
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendotheliosis, Systemic|9751/3
C0019621|T191|PM|D006646|MSH|Cell Granulomatoses, Langerhans|9751/3
C0019621|T191|PM|D006646|MSH|Cell Granulomatosis, Langerhans|9751/3
C0019621|T191|PM|D006646|MSH|Cell Histiocytoses, Langerhans|9751/3
C0019621|T191|PM|D006646|MSH|Cell Histiocytosis, Langerhans|9751/3
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schueller-Christian|9751/3
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schüller-Christian|9751/3
C0019621|T191|PM|D006646|MSH|Disease, Letterer-Siwe|9751/3
C0019621|T191|PM|D006646|MSH|Disease, Schueller-Christian|9751/3
C0019621|T191|PM|D006646|MSH|Generalized Histiocytoses|9751/3
C0019621|T191|PM|D006646|MSH|Generalized Histiocytosis|9751/3
C0019621|T191|PM|D006646|MSH|Granulomatoses, Langerhans Cell|9751/3
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans Cell|9751/3
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans-Cell|9751/3
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Disease|9751/3
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Syndrome|9751/3
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Disease|9751/3
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Syndrome|9751/3
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Disease|9751/3
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Syndrome|9751/3
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Disease|9751/3
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Syndrome|9751/3
C0019621|T191|PM|D006646|MSH|Histiocytoses, Generalized|9751/3
C0019621|T191|PM|D006646|MSH|Histiocytoses, Langerhans Cell|9751/3
C0019621|T191|PM|D006646|MSH|Histiocytoses, Type 2|9751/3
C0019621|T191|ET|D006646|MSH|Histiocytosis X|9751/3
C0019621|T191|ET|D006646|MSH|Histiocytosis-X|9751/3
C0019621|T191|ET|D006646|MSH|Histiocytosis, Generalized|9751/3
C0019621|T191|PM|D006646|MSH|Histiocytosis, Langerhans Cell|9751/3
C0019621|T191|MH|D006646|MSH|Histiocytosis, Langerhans-Cell|9751/3
C0019621|T191|PM|D006646|MSH|Histiocytosis, Type 2|9751/3
C0019621|T191|PM|D006646|MSH|Langerhans Cell Granulomatoses|9751/3
C0019621|T191|ET|D006646|MSH|Langerhans Cell Granulomatosis|9751/3
C0019621|T191|PM|D006646|MSH|Langerhans Cell Histiocytoses|9751/3
C0019621|T191|ET|D006646|MSH|Langerhans Cell Histiocytosis|9751/3
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Granulomatosis|9751/3
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Histiocytosis|9751/3
C0019621|T191|DEV|D006646|MSH|LETTERER SIWE DIS|9751/3
C0019621|T191|PM|D006646|MSH|Letterer Siwe Disease|9751/3
C0019621|T191|ET|D006646|MSH|Letterer-Siwe Disease|9751/3
C0019621|T191|PM|D006646|MSH|Non Lipid Reticuloendotheliosis|9751/3
C0019621|T191|PM|D006646|MSH|Non-Lipid Reticuloendothelioses|9751/3
C0019621|T191|ET|D006646|MSH|Non-Lipid Reticuloendotheliosis|9751/3
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Non-Lipid|9751/3
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Systemic Aleukemic|9751/3
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Non-Lipid|9751/3
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Systemic Aleukemic|9751/3
C0019621|T191|DEV|D006646|MSH|SCHUELLER CHRISTIAN DIS|9751/3
C0019621|T191|PM|D006646|MSH|Schueller Christian Disease|9751/3
C0019621|T191|ET|D006646|MSH|Schueller-Christian Disease|9751/3
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schueller-Christian|9751/3
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schüller-Christian|9751/3
C0019621|T191|PM|D006646|MSH|Systemic Aleukemic Reticuloendothelioses|9751/3
C0019621|T191|ET|D006646|MSH|Systemic Aleukemic Reticuloendotheliosis|9751/3
C0019621|T191|PM|D006646|MSH|Type 2 Histiocytoses|9751/3
C0019621|T191|ET|D006646|MSH|Type 2 Histiocytosis|9751/3
C0019621|T191|PN|NOCODE|MTH|Histiocytosis, Langerhans-Cell|9751/3
C0019621|T191|ET|277.89|MTHICD9|Chronic Histiocytosis X|9751/3
C0019621|T191|ET|277.89|MTHICD9|Hand-Schuller-Christian disease|9751/3
C0019621|T191|ET|277.89|MTHICD9|Histiocytosis X|9751/3
C0019621|T191|PT|C6920|NCI|Hand-Schuller-Christian Disease|9751/3
C0019621|T191|OP|C3107|NCI|Histiocytosis X|9751/3
C0019621|T191|SY|C3107|NCI|Langerhans Cell Granulomatosis|9751/3
C0019621|T191|PT|C3107|NCI|Langerhans Cell Histiocytosis|9751/3
C0019621|T191|SY|TCGA|NCI|Langerhans Cell Histiocytosis|9751/3
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, NOS|9751/3
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, Not Otherwise Specified|9751/3
C0019621|T191|AB|C3107|NCI|LCH|9751/3
C0019621|T191|PT|C6920|NCI_CPTAC|Hand-Schuller-Christian Disease|9751/3
C0019621|T191|PT|10025581|NCI_CTEP-SDC|Langerhans cell histiocytosis|9751/3
C0019621|T191|DN|C3107|NCI_CTRP|Langerhans Cell Histiocytosis|9751/3
C0019621|T191|PT|CDR0000471787|NCI_NCI-GLOSS|Langerhans cell histiocytosis|9751/3
C0019621|T191|PT|CDR0000513054|NCI_NCI-GLOSS|LCH|9751/3
C0019621|T191|SY|C6920|NCI_NICHD|Classic Multifocal Langerhans Cell Histiocytosis|9751/3
C0019621|T191|SY|C6920|NCI_NICHD|Hand-Schüller-Christian Disease|9751/3
C0019621|T191|OP|C3107|NCI_NICHD|Histiocytosis X|9751/3
C0019621|T191|PT|C3107|NCI_NICHD|Langerhans Cell Histiocytosis|9751/3
C0019621|T191|PT|C6920|NCI_NICHD|Multifocal Unisystem Langerhans Cell Histiocytosis|9751/3
C0019621|T191|SY|CDR0000039054|PDQ|histiocytosis X|9751/3
C0019621|T191|PT|CDR0000641624|PDQ|Langerhans cell histiocytosis|9751/3
C0019621|T191|AB|X20E9|RCD|Different progress histiocyto|9751/3
C0019621|T191|SY|X20E9|RCD|Differentiated progressive histiocytosis|9751/3
C0019621|T191|AB|C37y0|RCD|Hand-Schuller-Christian diseas|9751/3
C0019621|T191|SY|C37y0|RCD|Hand-Schuller-Christian disease|9751/3
C0019621|T191|OP|C37y6|RCD|Histiocytosis X , unspecified|9751/3
C0019621|T191|PT|C37y5|RCD|Histiocytosis X syndrome|9751/3
C0019621|T191|PT|X20E9|RCD|Langerhan's cell histiocytosis|9751/3
C0019621|T191|AB|X20E9|RCD|Langerhans histiocyt syndrome|9751/3
C0019621|T191|SY|X20E9|RCD|Langerhans histiocytic syndrome|9751/3
C0019621|T191|SY|X20E9|RCD|LCH - Langerhan's cell histiocytosis|9751/3
C0019621|T191|AB|X20E9|RCD|LCH-Langerh cell histiocytosis|9751/3
C0019621|T191|PT|C37y0|RCD|Schuller-Christian syndrome|9751/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic differentiated progressive histiocytosis|9751/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic disseminated histiocytosis X|9751/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic histiocytosis X|9751/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic idiopathic xanthomatosis|9751/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|Differentiated progressive histiocytosis|9751/3
C0019621|T191|SY|65399007|SNOMEDCT_US|Differentiated progressive histiocytosis|9751/3
C0019621|T191|SYGB|39795003|SNOMEDCT_US|Generalised histiocytosis of bones|9751/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Generalized histiocytosis of bones|9751/3
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand - Schuller - Christian disease|9751/3
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand - Schuller - Christian disease|9751/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Hand-Schuller-Christian disease|9751/3
C0019621|T191|PT|39795003|SNOMEDCT_US|Hand-Schüller-Christian disease|9751/3
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9751/3
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9751/3
C0019621|T191|SY|65399007|SNOMEDCT_US|Histiocytosis X|9751/3
C0019621|T191|OAS|154583006|SNOMEDCT_US|Histiocytosis X|9751/3
C0019621|T191|OAS|269628007|SNOMEDCT_US|Histiocytosis X|9751/3
C0019621|T191|IS|190960001|SNOMEDCT_US|Histiocytosis X , chronic|9751/3
C0019621|T191|IS|190956004|SNOMEDCT_US|Histiocytosis X , unspecified|9751/3
C0019621|T191|PT|190955000|SNOMEDCT_US|Histiocytosis X syndrome|9751/3
C0019621|T191|IS|65399007|SNOMEDCT_US|Histiocytosis X, NOS|9751/3
C0019621|T191|OAP|190956004|SNOMEDCT_US|Histiocytosis X, unspecified|9751/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhan's cell histiocytosis|9751/3
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhan's cell histiocytosis|9751/3
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhans cell disease|9751/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans cell disease|9751/3
C0019621|T191|IS|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9751/3
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9751/3
C0019621|T191|PT|65399007|SNOMEDCT_US|Langerhans cell histiocytosis|9751/3
C0019621|T191|PT|128809007|SNOMEDCT_US|Langerhans cell histiocytosis|9751/3
C0019621|T191|OAP|234439008|SNOMEDCT_US|Langerhans cell histiocytosis|9751/3
C0019621|T191|PT|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, multifocal|9751/3
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no ICD-O subtype|9751/3
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no International Classification of Diseases for Oncology subtype|9751/3
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, poly-ostotic|9751/3
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, polyostotic|9751/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans histiocytic syndrome|9751/3
C0019621|T191|OAP|110450007|SNOMEDCT_US|Langerhans' cell histiocytosis|9751/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9751/3
C0019621|T191|SY|65399007|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9751/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Multifocal and unisystemic Langerhans cell histiocytosis|9751/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Schuller-Christian syndrome|9751/3
C0019621|T191|SY|0000006165|CHV|cell granulomatosis langerhans|9752/1
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhan|9752/1
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhans|9752/1
C0019621|T191|SY|0000006165|CHV|cells histiocytosis langerhans|9752/1
C0019621|T191|SY|0000026274|CHV|christian disease hand schuller|9752/1
C0019621|T191|SY|0000026274|CHV|christian diseases hand schuller|9752/1
C0019621|T191|SY|0000026274|CHV|disease hand schuller christian|9752/1
C0014461|T046|PT|0000004531|CHV|eosinophilic granuloma|9752/1
C0019621|T191|SY|0000007324|CHV|generalized histiocytosis|9752/1
C0014461|T046|SY|0000004531|CHV|granuloma eosinophilic|9752/1
C0019621|T191|SY|0000026274|CHV|hand christian schuller disease|9752/1
C0019621|T191|SY|0000026274|CHV|hand schuller christian disease|9752/1
C0019621|T191|SY|0000026274|CHV|hand-schueller-christian disease|9752/1
C0019621|T191|PT|0000026274|CHV|hand-schuller-christian disease|9752/1
C0019621|T191|PT|0000006165|CHV|histiocytosis x|9752/1
C0019621|T191|SY|0000006165|CHV|histiocytosis-x|9752/1
C0019621|T191|SY|0000006165|CHV|langerhan's cell histiocytosis|9752/1
C0019621|T191|SY|0000006165|CHV|langerhans cell disease|9752/1
C0019621|T191|SY|0000006165|CHV|langerhans cell granulomatosis|9752/1
C0019621|T191|SY|0000006165|CHV|langerhans cell histiocytosis|9752/1
C0019621|T191|SY|0000026274|CHV|schuller christian syndrome|9752/1
C0014461|T046|PT|NOCODE|COSTAR|Eosinophilic Granuloma|9752/1
C0014461|T046|PT|0427-5503|CSP|eosinophilic granuloma|9752/1
C0019621|T191|ET|0427-5330|CSP|Hand Schuller Christian disease|9752/1
C0019621|T191|PT|0427-5330|CSP|histiocytosis X|9752/1
C0019621|T191|ET|0427-5330|CSP|Langerhans cell granulomatosis|9752/1
C0014461|T046|GT|GRANULOMA|CST|EOSINOPHILIC GRANULOMA|9752/1
C0014461|T046|DI|U000571|DXP|EOSINOPHILIC GRANULOMA|9752/1
C0019621|T191|SY|NOCODE|DXP|EOSINOPHILIC GRANULOMA, MULTIFOCAL|9752/1
C0019621|T191|DI|U000766|DXP|HAND-SCHUELLER-CHRISTIAN SYNDROME|9752/1
C0019621|T191|SY|NOCODE|DXP|HISTIOCYTOSIS X II|9752/1
C0019621|T191|SY|NOCODE|DXP|SCHUELLER-CHRISTIAN DISEASE|9752/1
C0014461|T046|PT|HP:0032253|HPO|Eosinophilic granuloma|9752/1
C0014461|T046|ET|K13.4|ICD10CM|Eosinophilic granuloma|9752/1
C0014461|T046|ET|C96.6|ICD10CM|Eosinophilic granuloma|9752/1
C0019621|T191|ET|C96.5|ICD10CM|Hand-Schüller-Christian disease|9752/1
C0019621|T191|ET|C96.6|ICD10CM|Langerhans-cell histiocytosis NOS|9752/1
C1306599|T191|PT|C96.6|ICD10CM|Unifocal Langerhans-cell histiocytosis|9752/1
C1306599|T191|AB|C96.6|ICD10CM|Unifocal Langerhans-cell histiocytosis|9752/1
C0014461|T046|PT|MTHU026437|ICPC2ICD10ENG|eosinophilic; granuloma|9752/1
C0014461|T046|PT|MTHU032745|ICPC2ICD10ENG|granuloma; eosinophilic|9752/1
C0019621|T191|PT|MTHU033317|ICPC2ICD10ENG|Hand-Schüller-Christian|9752/1
C0019621|T191|PT|MTHU035172|ICPC2ICD10ENG|histiocytosis; Langerhans' cell|9752/1
C0019621|T191|PT|MTHU035180|ICPC2ICD10ENG|histiocytosis; X|9752/1
C0019621|T191|PT|MTHU035182|ICPC2ICD10ENG|histiocytosis; X, chronic|9752/1
C0019621|T191|PT|MTHU042862|ICPC2ICD10ENG|Langerhans' cell; histiocytosis|9752/1
C0019621|T191|PT|MTHU066496|ICPC2ICD10ENG|Schüller-Christian|9752/1
C0019621|T191|PT|MTHU082788|ICPC2ICD10ENG|X; histiocytosis|9752/1
C0019621|T191|PT|MTHU082790|ICPC2ICD10ENG|X; histiocytosis, chronic|9752/1
C0014461|T046|PT|U001621|LCH|Eosinophilic granuloma|9752/1
C0019621|T191|PT|U002076|LCH|Hand-Schueller-Christian syndrome|9752/1
C0014461|T046|PT|sh85044244|LCH_NW|Eosinophilic granuloma|9752/1
C0019621|T191|PT|sh85058638|LCH_NW|Hand-Schueller-Christian syndrome|9752/1
C0019621|T191|LLT|10053133|MDR|Chronic idiopathic xanthomatosis|9752/1
C0014461|T046|LLT|10014956|MDR|Eosinophilic granuloma|9752/1
C0019621|T191|LLT|10053135|MDR|Hand-Schueller-Christian disease|9752/1
C0019621|T191|LLT|10023688|MDR|Langerhans' cell granulomatosis|9752/1
C0019621|T191|PT|10069698|MDR|Langerhans' cell histiocytosis|9752/1
C0019621|T191|LLT|10069698|MDR|Langerhans' cell histiocytosis|9752/1
C0014461|T046|PT|97091|MEDCIN|eosinophilic granuloma|9752/1
C0019621|T191|SY|31815|MEDCIN|Hand-Schuller-Christian disease|9752/1
C0014461|T046|PT|31814|MEDCIN|histiocytoses - unifocal eosinophilic granuloma|9752/1
C0019621|T191|PT|315032|MEDCIN|Langerhans cell histiocytosis|9752/1
C0019621|T191|PT|31815|MEDCIN|multifocal eosinophilic granuloma|9752/1
C0014461|T046|SY|31814|MEDCIN|unifocal eosinophilic granuloma|9752/1
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendothelioses, Systemic|9752/1
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendotheliosis, Systemic|9752/1
C0019621|T191|PM|D006646|MSH|Cell Granulomatoses, Langerhans|9752/1
C0019621|T191|PM|D006646|MSH|Cell Granulomatosis, Langerhans|9752/1
C0019621|T191|PM|D006646|MSH|Cell Histiocytoses, Langerhans|9752/1
C0019621|T191|PM|D006646|MSH|Cell Histiocytosis, Langerhans|9752/1
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schueller-Christian|9752/1
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schüller-Christian|9752/1
C0019621|T191|PM|D006646|MSH|Disease, Letterer-Siwe|9752/1
C0019621|T191|PM|D006646|MSH|Disease, Schueller-Christian|9752/1
C0014461|T046|MH|D004803|MSH|Eosinophilic Granuloma|9752/1
C0014461|T046|PM|D004803|MSH|Eosinophilic Granulomas|9752/1
C0019621|T191|PM|D006646|MSH|Generalized Histiocytoses|9752/1
C0019621|T191|PM|D006646|MSH|Generalized Histiocytosis|9752/1
C0014461|T046|ET|D004803|MSH|Granuloma, Eosinophilic|9752/1
C0014461|T046|PM|D004803|MSH|Granulomas, Eosinophilic|9752/1
C0019621|T191|PM|D006646|MSH|Granulomatoses, Langerhans Cell|9752/1
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans Cell|9752/1
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans-Cell|9752/1
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Disease|9752/1
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Syndrome|9752/1
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Disease|9752/1
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Syndrome|9752/1
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Disease|9752/1
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Syndrome|9752/1
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Disease|9752/1
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Syndrome|9752/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Generalized|9752/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Langerhans Cell|9752/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Type 2|9752/1
C0019621|T191|ET|D006646|MSH|Histiocytosis X|9752/1
C0019621|T191|ET|D006646|MSH|Histiocytosis-X|9752/1
C0019621|T191|ET|D006646|MSH|Histiocytosis, Generalized|9752/1
C0019621|T191|PM|D006646|MSH|Histiocytosis, Langerhans Cell|9752/1
C0019621|T191|MH|D006646|MSH|Histiocytosis, Langerhans-Cell|9752/1
C0019621|T191|PM|D006646|MSH|Histiocytosis, Type 2|9752/1
C0019621|T191|PM|D006646|MSH|Langerhans Cell Granulomatoses|9752/1
C0019621|T191|ET|D006646|MSH|Langerhans Cell Granulomatosis|9752/1
C0019621|T191|PM|D006646|MSH|Langerhans Cell Histiocytoses|9752/1
C0019621|T191|ET|D006646|MSH|Langerhans Cell Histiocytosis|9752/1
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Granulomatosis|9752/1
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Histiocytosis|9752/1
C0019621|T191|DEV|D006646|MSH|LETTERER SIWE DIS|9752/1
C0019621|T191|PM|D006646|MSH|Letterer Siwe Disease|9752/1
C0019621|T191|ET|D006646|MSH|Letterer-Siwe Disease|9752/1
C0019621|T191|PM|D006646|MSH|Non Lipid Reticuloendotheliosis|9752/1
C0019621|T191|PM|D006646|MSH|Non-Lipid Reticuloendothelioses|9752/1
C0019621|T191|ET|D006646|MSH|Non-Lipid Reticuloendotheliosis|9752/1
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Non-Lipid|9752/1
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Systemic Aleukemic|9752/1
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Non-Lipid|9752/1
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Systemic Aleukemic|9752/1
C0019621|T191|DEV|D006646|MSH|SCHUELLER CHRISTIAN DIS|9752/1
C0019621|T191|PM|D006646|MSH|Schueller Christian Disease|9752/1
C0019621|T191|ET|D006646|MSH|Schueller-Christian Disease|9752/1
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schueller-Christian|9752/1
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schüller-Christian|9752/1
C0019621|T191|PM|D006646|MSH|Systemic Aleukemic Reticuloendothelioses|9752/1
C0019621|T191|ET|D006646|MSH|Systemic Aleukemic Reticuloendotheliosis|9752/1
C0019621|T191|PM|D006646|MSH|Type 2 Histiocytoses|9752/1
C0019621|T191|ET|D006646|MSH|Type 2 Histiocytosis|9752/1
C0019621|T191|PN|NOCODE|MTH|Histiocytosis, Langerhans-Cell|9752/1
C0019621|T191|ET|277.89|MTHICD9|Chronic Histiocytosis X|9752/1
C0019621|T191|ET|277.89|MTHICD9|Hand-Schuller-Christian disease|9752/1
C0019621|T191|ET|277.89|MTHICD9|Histiocytosis X|9752/1
C0014461|T046|PT|C3016|NCI|Eosinophilic Granuloma|9752/1
C0014461|T046|SY|C3016|NCI|Eosinophilic Xanthomatous Granuloma|9752/1
C0019621|T191|PT|C6920|NCI|Hand-Schuller-Christian Disease|9752/1
C0019621|T191|OP|C3107|NCI|Histiocytosis X|9752/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Granulomatosis|9752/1
C0019621|T191|PT|C3107|NCI|Langerhans Cell Histiocytosis|9752/1
C0019621|T191|SY|TCGA|NCI|Langerhans Cell Histiocytosis|9752/1
C1306599|T191|PT|C150701|NCI|Langerhans Cell Histiocytosis, Monostotic|9752/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, NOS|9752/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, Not Otherwise Specified|9752/1
C0019621|T191|AB|C3107|NCI|LCH|9752/1
C0019621|T191|PT|C6920|NCI_CPTAC|Hand-Schuller-Christian Disease|9752/1
C0019621|T191|PT|10025581|NCI_CTEP-SDC|Langerhans cell histiocytosis|9752/1
C0019621|T191|DN|C3107|NCI_CTRP|Langerhans Cell Histiocytosis|9752/1
C0019621|T191|PT|CDR0000471787|NCI_NCI-GLOSS|Langerhans cell histiocytosis|9752/1
C0019621|T191|PT|CDR0000513054|NCI_NCI-GLOSS|LCH|9752/1
C0014461|T046|SY|C3016|NCI_NICHD|Chronic Unifocal Langerhans Cell Histiocytosis|9752/1
C0019621|T191|SY|C6920|NCI_NICHD|Classic Multifocal Langerhans Cell Histiocytosis|9752/1
C0014461|T046|SY|C3016|NCI_NICHD|Eosinophilic Granuloma|9752/1
C0014461|T046|SY|C3016|NCI_NICHD|Eosinophilic Xanthomatous Granuloma|9752/1
C0019621|T191|SY|C6920|NCI_NICHD|Hand-Schüller-Christian Disease|9752/1
C0019621|T191|OP|C3107|NCI_NICHD|Histiocytosis X|9752/1
C0019621|T191|PT|C3107|NCI_NICHD|Langerhans Cell Histiocytosis|9752/1
C0014461|T046|SY|C3016|NCI_NICHD|Monostotic Langerhans Cell Histiocytosis|9752/1
C0019621|T191|PT|C6920|NCI_NICHD|Multifocal Unisystem Langerhans Cell Histiocytosis|9752/1
C0014461|T046|PT|C3016|NCI_NICHD|Unifocal Langerhans Cell Histiocytosis|9752/1
C0019621|T191|SY|CDR0000039054|PDQ|histiocytosis X|9752/1
C0019621|T191|PT|CDR0000641624|PDQ|Langerhans cell histiocytosis|9752/1
C0019621|T191|AB|X20E9|RCD|Different progress histiocyto|9752/1
C0019621|T191|SY|X20E9|RCD|Differentiated progressive histiocytosis|9752/1
C0014461|T046|PT|C37y1|RCD|Eosinophilic granuloma|9752/1
C0014461|T046|AB|C37y1|RCD|Eosinophilic xanthom granuloma|9752/1
C0014461|T046|SY|C37y1|RCD|Eosinophilic xanthomatous granuloma|9752/1
C0019621|T191|AB|C37y0|RCD|Hand-Schuller-Christian diseas|9752/1
C0019621|T191|SY|C37y0|RCD|Hand-Schuller-Christian disease|9752/1
C0019621|T191|OP|C37y6|RCD|Histiocytosis X , unspecified|9752/1
C0019621|T191|PT|C37y5|RCD|Histiocytosis X syndrome|9752/1
C0019621|T191|PT|X20E9|RCD|Langerhan's cell histiocytosis|9752/1
C0019621|T191|AB|X20E9|RCD|Langerhans histiocyt syndrome|9752/1
C0019621|T191|SY|X20E9|RCD|Langerhans histiocytic syndrome|9752/1
C0019621|T191|SY|X20E9|RCD|LCH - Langerhan's cell histiocytosis|9752/1
C0019621|T191|AB|X20E9|RCD|LCH-Langerh cell histiocytosis|9752/1
C0019621|T191|PT|C37y0|RCD|Schuller-Christian syndrome|9752/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic differentiated progressive histiocytosis|9752/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic disseminated histiocytosis X|9752/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic histiocytosis X|9752/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic idiopathic xanthomatosis|9752/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Differentiated progressive histiocytosis|9752/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Differentiated progressive histiocytosis|9752/1
C0014461|T046|SY|129000002|SNOMEDCT_US|Eosinophilic granuloma|9752/1
C0014461|T046|SY|128810002|SNOMEDCT_US|Eosinophilic granuloma|9752/1
C0014461|T046|OAP|77239009|SNOMEDCT_US|Eosinophilic granuloma|9752/1
C0014461|T046|IS|77239009|SNOMEDCT_US|Eosinophilic granuloma -RETIRED-|9752/1
C0014461|T046|OF|77239009|SNOMEDCT_US|Eosinophilic granuloma -RETIRED-|9752/1
C0014461|T046|IS|77239009|SNOMEDCT_US|Eosinophilic xanthomatous granuloma|9752/1
C0014461|T046|SY|129000002|SNOMEDCT_US|Eosinophilic xanthomatous granuloma|9752/1
C0019621|T191|SYGB|39795003|SNOMEDCT_US|Generalised histiocytosis of bones|9752/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Generalized histiocytosis of bones|9752/1
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand - Schuller - Christian disease|9752/1
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand - Schuller - Christian disease|9752/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Hand-Schuller-Christian disease|9752/1
C0019621|T191|PT|39795003|SNOMEDCT_US|Hand-Schüller-Christian disease|9752/1
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9752/1
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9752/1
C0019621|T191|OAS|269628007|SNOMEDCT_US|Histiocytosis X|9752/1
C0019621|T191|OAS|154583006|SNOMEDCT_US|Histiocytosis X|9752/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Histiocytosis X|9752/1
C0019621|T191|IS|190960001|SNOMEDCT_US|Histiocytosis X , chronic|9752/1
C0019621|T191|IS|190956004|SNOMEDCT_US|Histiocytosis X , unspecified|9752/1
C0019621|T191|PT|190955000|SNOMEDCT_US|Histiocytosis X syndrome|9752/1
C0019621|T191|IS|65399007|SNOMEDCT_US|Histiocytosis X, NOS|9752/1
C0019621|T191|OAP|190956004|SNOMEDCT_US|Histiocytosis X, unspecified|9752/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhan's cell histiocytosis|9752/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhan's cell histiocytosis|9752/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans cell disease|9752/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhans cell disease|9752/1
C0019621|T191|IS|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9752/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9752/1
C1306599|T191|SY|128810002|SNOMEDCT_US|Langerhans cell granulomatosis, unifocal|9752/1
C0019621|T191|OAP|234439008|SNOMEDCT_US|Langerhans cell histiocytosis|9752/1
C0019621|T191|PT|65399007|SNOMEDCT_US|Langerhans cell histiocytosis|9752/1
C0019621|T191|PT|128809007|SNOMEDCT_US|Langerhans cell histiocytosis|9752/1
C1306599|T191|SY|128810002|SNOMEDCT_US|Langerhans cell histiocytosis, mono-ostotic|9752/1
C1306599|T191|SY|128810002|SNOMEDCT_US|Langerhans cell histiocytosis, monostotic|9752/1
C0019621|T191|PT|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, multifocal|9752/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no ICD-O subtype|9752/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no International Classification of Diseases for Oncology subtype|9752/1
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, poly-ostotic|9752/1
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, polyostotic|9752/1
C1306599|T191|PT|128810002|SNOMEDCT_US|Langerhans cell histiocytosis, unifocal|9752/1
C1306599|T191|SY|129000002|SNOMEDCT_US|Langerhans cell histiocytosis, unifocal|9752/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans histiocytic syndrome|9752/1
C0019621|T191|OAP|110450007|SNOMEDCT_US|Langerhans' cell histiocytosis|9752/1
C0019621|T191|SY|65399007|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9752/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9752/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Multifocal and unisystemic Langerhans cell histiocytosis|9752/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Schuller-Christian syndrome|9752/1
C0014461|T046|PT|0815|WHO|EOSINOPHILIC GRANULOMA|9752/1
C0019621|T191|SY|0000006165|CHV|cell granulomatosis langerhans|9753/1
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhan|9753/1
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhans|9753/1
C0019621|T191|SY|0000006165|CHV|cells histiocytosis langerhans|9753/1
C0019621|T191|SY|0000026274|CHV|christian disease hand schuller|9753/1
C0019621|T191|SY|0000026274|CHV|christian diseases hand schuller|9753/1
C0019621|T191|SY|0000026274|CHV|disease hand schuller christian|9753/1
C0019621|T191|SY|0000007324|CHV|generalized histiocytosis|9753/1
C0019621|T191|SY|0000026274|CHV|hand christian schuller disease|9753/1
C0019621|T191|SY|0000026274|CHV|hand schuller christian disease|9753/1
C0019621|T191|SY|0000026274|CHV|hand-schueller-christian disease|9753/1
C0019621|T191|PT|0000026274|CHV|hand-schuller-christian disease|9753/1
C0019621|T191|PT|0000006165|CHV|histiocytosis x|9753/1
C0019621|T191|SY|0000006165|CHV|histiocytosis-x|9753/1
C0019621|T191|SY|0000006165|CHV|langerhan's cell histiocytosis|9753/1
C0019621|T191|SY|0000006165|CHV|langerhans cell disease|9753/1
C0019621|T191|SY|0000006165|CHV|langerhans cell granulomatosis|9753/1
C0019621|T191|SY|0000006165|CHV|langerhans cell histiocytosis|9753/1
C0019621|T191|SY|0000026274|CHV|schuller christian syndrome|9753/1
C0019621|T191|ET|0427-5330|CSP|Hand Schuller Christian disease|9753/1
C0019621|T191|PT|0427-5330|CSP|histiocytosis X|9753/1
C0019621|T191|ET|0427-5330|CSP|Langerhans cell granulomatosis|9753/1
C0019621|T191|SY|NOCODE|DXP|EOSINOPHILIC GRANULOMA, MULTIFOCAL|9753/1
C0019621|T191|DI|U000766|DXP|HAND-SCHUELLER-CHRISTIAN SYNDROME|9753/1
C0019621|T191|SY|NOCODE|DXP|HISTIOCYTOSIS X II|9753/1
C0019621|T191|SY|NOCODE|DXP|SCHUELLER-CHRISTIAN DISEASE|9753/1
C0019621|T191|ET|C96.5|ICD10CM|Hand-Schüller-Christian disease|9753/1
C0019621|T191|ET|C96.6|ICD10CM|Langerhans-cell histiocytosis NOS|9753/1
C0019621|T191|PT|MTHU033317|ICPC2ICD10ENG|Hand-Schüller-Christian|9753/1
C0019621|T191|PT|MTHU035172|ICPC2ICD10ENG|histiocytosis; Langerhans' cell|9753/1
C0019621|T191|PT|MTHU035180|ICPC2ICD10ENG|histiocytosis; X|9753/1
C0019621|T191|PT|MTHU035182|ICPC2ICD10ENG|histiocytosis; X, chronic|9753/1
C0019621|T191|PT|MTHU042862|ICPC2ICD10ENG|Langerhans' cell; histiocytosis|9753/1
C0019621|T191|PT|MTHU066496|ICPC2ICD10ENG|Schüller-Christian|9753/1
C0019621|T191|PT|MTHU082788|ICPC2ICD10ENG|X; histiocytosis|9753/1
C0019621|T191|PT|MTHU082790|ICPC2ICD10ENG|X; histiocytosis, chronic|9753/1
C0019621|T191|PT|U002076|LCH|Hand-Schueller-Christian syndrome|9753/1
C0019621|T191|PT|sh85058638|LCH_NW|Hand-Schueller-Christian syndrome|9753/1
C0019621|T191|LLT|10053133|MDR|Chronic idiopathic xanthomatosis|9753/1
C0019621|T191|LLT|10053135|MDR|Hand-Schueller-Christian disease|9753/1
C0019621|T191|LLT|10023688|MDR|Langerhans' cell granulomatosis|9753/1
C0019621|T191|LLT|10069698|MDR|Langerhans' cell histiocytosis|9753/1
C0019621|T191|PT|10069698|MDR|Langerhans' cell histiocytosis|9753/1
C0019621|T191|SY|31815|MEDCIN|Hand-Schuller-Christian disease|9753/1
C0019621|T191|PT|315032|MEDCIN|Langerhans cell histiocytosis|9753/1
C0019621|T191|PT|31815|MEDCIN|multifocal eosinophilic granuloma|9753/1
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendothelioses, Systemic|9753/1
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendotheliosis, Systemic|9753/1
C0019621|T191|PM|D006646|MSH|Cell Granulomatoses, Langerhans|9753/1
C0019621|T191|PM|D006646|MSH|Cell Granulomatosis, Langerhans|9753/1
C0019621|T191|PM|D006646|MSH|Cell Histiocytoses, Langerhans|9753/1
C0019621|T191|PM|D006646|MSH|Cell Histiocytosis, Langerhans|9753/1
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schueller-Christian|9753/1
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schüller-Christian|9753/1
C0019621|T191|PM|D006646|MSH|Disease, Letterer-Siwe|9753/1
C0019621|T191|PM|D006646|MSH|Disease, Schueller-Christian|9753/1
C0019621|T191|PM|D006646|MSH|Generalized Histiocytoses|9753/1
C0019621|T191|PM|D006646|MSH|Generalized Histiocytosis|9753/1
C0019621|T191|PM|D006646|MSH|Granulomatoses, Langerhans Cell|9753/1
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans Cell|9753/1
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans-Cell|9753/1
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Disease|9753/1
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Syndrome|9753/1
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Disease|9753/1
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Syndrome|9753/1
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Disease|9753/1
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Syndrome|9753/1
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Disease|9753/1
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Syndrome|9753/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Generalized|9753/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Langerhans Cell|9753/1
C0019621|T191|PM|D006646|MSH|Histiocytoses, Type 2|9753/1
C0019621|T191|ET|D006646|MSH|Histiocytosis X|9753/1
C0019621|T191|ET|D006646|MSH|Histiocytosis-X|9753/1
C0019621|T191|ET|D006646|MSH|Histiocytosis, Generalized|9753/1
C0019621|T191|PM|D006646|MSH|Histiocytosis, Langerhans Cell|9753/1
C0019621|T191|MH|D006646|MSH|Histiocytosis, Langerhans-Cell|9753/1
C0019621|T191|PM|D006646|MSH|Histiocytosis, Type 2|9753/1
C0019621|T191|PM|D006646|MSH|Langerhans Cell Granulomatoses|9753/1
C0019621|T191|ET|D006646|MSH|Langerhans Cell Granulomatosis|9753/1
C0019621|T191|PM|D006646|MSH|Langerhans Cell Histiocytoses|9753/1
C0019621|T191|ET|D006646|MSH|Langerhans Cell Histiocytosis|9753/1
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Granulomatosis|9753/1
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Histiocytosis|9753/1
C0019621|T191|DEV|D006646|MSH|LETTERER SIWE DIS|9753/1
C0019621|T191|PM|D006646|MSH|Letterer Siwe Disease|9753/1
C0019621|T191|ET|D006646|MSH|Letterer-Siwe Disease|9753/1
C0019621|T191|PM|D006646|MSH|Non Lipid Reticuloendotheliosis|9753/1
C0019621|T191|PM|D006646|MSH|Non-Lipid Reticuloendothelioses|9753/1
C0019621|T191|ET|D006646|MSH|Non-Lipid Reticuloendotheliosis|9753/1
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Non-Lipid|9753/1
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Systemic Aleukemic|9753/1
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Non-Lipid|9753/1
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Systemic Aleukemic|9753/1
C0019621|T191|DEV|D006646|MSH|SCHUELLER CHRISTIAN DIS|9753/1
C0019621|T191|PM|D006646|MSH|Schueller Christian Disease|9753/1
C0019621|T191|ET|D006646|MSH|Schueller-Christian Disease|9753/1
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schueller-Christian|9753/1
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schüller-Christian|9753/1
C0019621|T191|PM|D006646|MSH|Systemic Aleukemic Reticuloendothelioses|9753/1
C0019621|T191|ET|D006646|MSH|Systemic Aleukemic Reticuloendotheliosis|9753/1
C0019621|T191|PM|D006646|MSH|Type 2 Histiocytoses|9753/1
C0019621|T191|ET|D006646|MSH|Type 2 Histiocytosis|9753/1
C0019621|T191|PN|NOCODE|MTH|Histiocytosis, Langerhans-Cell|9753/1
C0019621|T191|ET|277.89|MTHICD9|Chronic Histiocytosis X|9753/1
C0019621|T191|ET|277.89|MTHICD9|Hand-Schuller-Christian disease|9753/1
C0019621|T191|ET|277.89|MTHICD9|Histiocytosis X|9753/1
C0019621|T191|PT|C6920|NCI|Hand-Schuller-Christian Disease|9753/1
C0019621|T191|OP|C3107|NCI|Histiocytosis X|9753/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Granulomatosis|9753/1
C0019621|T191|PT|C3107|NCI|Langerhans Cell Histiocytosis|9753/1
C0019621|T191|SY|TCGA|NCI|Langerhans Cell Histiocytosis|9753/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, NOS|9753/1
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, Not Otherwise Specified|9753/1
C0019621|T191|AB|C3107|NCI|LCH|9753/1
C0019621|T191|PT|C6920|NCI_CPTAC|Hand-Schuller-Christian Disease|9753/1
C0019621|T191|PT|10025581|NCI_CTEP-SDC|Langerhans cell histiocytosis|9753/1
C0019621|T191|DN|C3107|NCI_CTRP|Langerhans Cell Histiocytosis|9753/1
C0019621|T191|PT|CDR0000471787|NCI_NCI-GLOSS|Langerhans cell histiocytosis|9753/1
C0019621|T191|PT|CDR0000513054|NCI_NCI-GLOSS|LCH|9753/1
C0019621|T191|SY|C6920|NCI_NICHD|Classic Multifocal Langerhans Cell Histiocytosis|9753/1
C0019621|T191|SY|C6920|NCI_NICHD|Hand-Schüller-Christian Disease|9753/1
C0019621|T191|OP|C3107|NCI_NICHD|Histiocytosis X|9753/1
C0019621|T191|PT|C3107|NCI_NICHD|Langerhans Cell Histiocytosis|9753/1
C0019621|T191|PT|C6920|NCI_NICHD|Multifocal Unisystem Langerhans Cell Histiocytosis|9753/1
C0019621|T191|SY|CDR0000039054|PDQ|histiocytosis X|9753/1
C0019621|T191|PT|CDR0000641624|PDQ|Langerhans cell histiocytosis|9753/1
C0019621|T191|AB|X20E9|RCD|Different progress histiocyto|9753/1
C0019621|T191|SY|X20E9|RCD|Differentiated progressive histiocytosis|9753/1
C0019621|T191|AB|C37y0|RCD|Hand-Schuller-Christian diseas|9753/1
C0019621|T191|SY|C37y0|RCD|Hand-Schuller-Christian disease|9753/1
C0019621|T191|OP|C37y6|RCD|Histiocytosis X , unspecified|9753/1
C0019621|T191|PT|C37y5|RCD|Histiocytosis X syndrome|9753/1
C0019621|T191|PT|X20E9|RCD|Langerhan's cell histiocytosis|9753/1
C0019621|T191|AB|X20E9|RCD|Langerhans histiocyt syndrome|9753/1
C0019621|T191|SY|X20E9|RCD|Langerhans histiocytic syndrome|9753/1
C0019621|T191|SY|X20E9|RCD|LCH - Langerhan's cell histiocytosis|9753/1
C0019621|T191|AB|X20E9|RCD|LCH-Langerh cell histiocytosis|9753/1
C0019621|T191|PT|C37y0|RCD|Schuller-Christian syndrome|9753/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic differentiated progressive histiocytosis|9753/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic disseminated histiocytosis X|9753/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic histiocytosis X|9753/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic idiopathic xanthomatosis|9753/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Differentiated progressive histiocytosis|9753/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Differentiated progressive histiocytosis|9753/1
C0019621|T191|SYGB|39795003|SNOMEDCT_US|Generalised histiocytosis of bones|9753/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Generalized histiocytosis of bones|9753/1
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand - Schuller - Christian disease|9753/1
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand - Schuller - Christian disease|9753/1
C0019621|T191|PT|39795003|SNOMEDCT_US|Hand-Schüller-Christian disease|9753/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Hand-Schuller-Christian disease|9753/1
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9753/1
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9753/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Histiocytosis X|9753/1
C0019621|T191|OAS|154583006|SNOMEDCT_US|Histiocytosis X|9753/1
C0019621|T191|OAS|269628007|SNOMEDCT_US|Histiocytosis X|9753/1
C0019621|T191|IS|190960001|SNOMEDCT_US|Histiocytosis X , chronic|9753/1
C0019621|T191|IS|190956004|SNOMEDCT_US|Histiocytosis X , unspecified|9753/1
C0019621|T191|PT|190955000|SNOMEDCT_US|Histiocytosis X syndrome|9753/1
C0019621|T191|IS|65399007|SNOMEDCT_US|Histiocytosis X, NOS|9753/1
C0019621|T191|OAP|190956004|SNOMEDCT_US|Histiocytosis X, unspecified|9753/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhan's cell histiocytosis|9753/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhan's cell histiocytosis|9753/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans cell disease|9753/1
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhans cell disease|9753/1
C0019621|T191|IS|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9753/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9753/1
C0019621|T191|PT|65399007|SNOMEDCT_US|Langerhans cell histiocytosis|9753/1
C0019621|T191|PT|128809007|SNOMEDCT_US|Langerhans cell histiocytosis|9753/1
C0019621|T191|OAP|234439008|SNOMEDCT_US|Langerhans cell histiocytosis|9753/1
C0019621|T191|PT|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, multifocal|9753/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no ICD-O subtype|9753/1
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no International Classification of Diseases for Oncology subtype|9753/1
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, poly-ostotic|9753/1
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, polyostotic|9753/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans histiocytic syndrome|9753/1
C0019621|T191|OAP|110450007|SNOMEDCT_US|Langerhans' cell histiocytosis|9753/1
C0019621|T191|OAS|234439008|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9753/1
C0019621|T191|SY|65399007|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9753/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Multifocal and unisystemic Langerhans cell histiocytosis|9753/1
C0019621|T191|SY|39795003|SNOMEDCT_US|Schuller-Christian syndrome|9753/1
C0019621|T191|SY|0000006165|CHV|cell granulomatosis langerhans|9754/3
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhan|9754/3
C0019621|T191|SY|0000006165|CHV|cell histiocytosis langerhans|9754/3
C0019621|T191|SY|0000006165|CHV|cells histiocytosis langerhans|9754/3
C0019621|T191|SY|0000026274|CHV|christian disease hand schuller|9754/3
C0019621|T191|SY|0000026274|CHV|christian diseases hand schuller|9754/3
C0019621|T191|SY|0000026274|CHV|disease hand schuller christian|9754/3
C0019621|T191|SY|0000007324|CHV|generalized histiocytosis|9754/3
C0019621|T191|SY|0000026274|CHV|hand christian schuller disease|9754/3
C0019621|T191|SY|0000026274|CHV|hand schuller christian disease|9754/3
C0019621|T191|SY|0000026274|CHV|hand-schueller-christian disease|9754/3
C0019621|T191|PT|0000026274|CHV|hand-schuller-christian disease|9754/3
C0019621|T191|PT|0000006165|CHV|histiocytosis x|9754/3
C0023381|T047|PT|0000007324|CHV|histiocytosis x|9754/3
C0019621|T191|SY|0000006165|CHV|histiocytosis-x|9754/3
C0019621|T191|SY|0000006165|CHV|langerhan's cell histiocytosis|9754/3
C0019621|T191|SY|0000006165|CHV|langerhans cell disease|9754/3
C0019621|T191|SY|0000006165|CHV|langerhans cell granulomatosis|9754/3
C0019621|T191|SY|0000006165|CHV|langerhans cell histiocytosis|9754/3
C0023381|T047|SY|0000007324|CHV|letterer - siwe disease|9754/3
C0023381|T047|SY|0000007324|CHV|letterer siwe disease|9754/3
C0023381|T047|SY|0000007324|CHV|letterer-siwe disease|9754/3
C0019621|T191|SY|0000026274|CHV|schuller christian syndrome|9754/3
C0019621|T191|ET|0427-5330|CSP|Hand Schuller Christian disease|9754/3
C0019621|T191|PT|0427-5330|CSP|histiocytosis X|9754/3
C0019621|T191|ET|0427-5330|CSP|Langerhans cell granulomatosis|9754/3
C0023381|T047|ET|0427-5330|CSP|Letterer Siwe disease|9754/3
C0023381|T047|SY|NOCODE|DXP|ABT-LETTERER-SIWE DISEASE|9754/3
C0019621|T191|SY|NOCODE|DXP|EOSINOPHILIC GRANULOMA, MULTIFOCAL|9754/3
C0019621|T191|DI|U000766|DXP|HAND-SCHUELLER-CHRISTIAN SYNDROME|9754/3
C0023381|T047|SY|NOCODE|DXP|HISTIOCYTOSIS X I|9754/3
C0019621|T191|SY|NOCODE|DXP|HISTIOCYTOSIS X II|9754/3
C0023381|T047|DI|U001043|DXP|LETTERER-SIWE DISEASE|9754/3
C0023381|T047|SY|NOCODE|DXP|RETICULOENDOTHELIOSIS, SYSTEMIC ALEUKEMIC|9754/3
C0019621|T191|SY|NOCODE|DXP|SCHUELLER-CHRISTIAN DISEASE|9754/3
C0023381|T047|PT|C96.0|ICD10|Letterer-Siwe disease|9754/3
C0019621|T191|ET|C96.5|ICD10CM|Hand-Schüller-Christian disease|9754/3
C0023381|T047|ET|C96.6|ICD10CM|Histiocytosis X NOS|9754/3
C0019621|T191|ET|C96.6|ICD10CM|Langerhans-cell histiocytosis NOS|9754/3
C0023381|T047|ET|C96.0|ICD10CM|Letterer-Siwe disease|9754/3
C0023381|T047|HT|202.5|ICD9CM|Letterer-Siwe disease|9754/3
C0023381|T047|PT|MTHU003129|ICPC2ICD10ENG|acute; differentiated progressive, histiocytosis|9754/3
C0023381|T047|PT|MTHU003204|ICPC2ICD10ENG|acute; reticuloendotheliosis, acute infantile|9754/3
C0019621|T191|PT|MTHU033317|ICPC2ICD10ENG|Hand-Schüller-Christian|9754/3
C0023381|T047|PT|MTHU035171|ICPC2ICD10ENG|histiocytosis; acute differentiated progressive|9754/3
C0019621|T191|PT|MTHU035172|ICPC2ICD10ENG|histiocytosis; Langerhans' cell|9754/3
C0019621|T191|PT|MTHU035180|ICPC2ICD10ENG|histiocytosis; X|9754/3
C0019621|T191|PT|MTHU035182|ICPC2ICD10ENG|histiocytosis; X, chronic|9754/3
C0019621|T191|PT|MTHU042862|ICPC2ICD10ENG|Langerhans' cell; histiocytosis|9754/3
C0023381|T047|PT|MTHU044732|ICPC2ICD10ENG|Letterer-Siwe|9754/3
C0023381|T047|PT|MTHU053302|ICPC2ICD10ENG|nonlipid; reticuloendotheliosis|9754/3
C0023381|T047|PT|MTHU064350|ICPC2ICD10ENG|reticuloendotheliosis; acute infantile|9754/3
C0023381|T047|PT|MTHU064353|ICPC2ICD10ENG|reticuloendotheliosis; nonlipid|9754/3
C0019621|T191|PT|MTHU066496|ICPC2ICD10ENG|Schüller-Christian|9754/3
C0019621|T191|PT|MTHU082788|ICPC2ICD10ENG|X; histiocytosis|9754/3
C0019621|T191|PT|MTHU082790|ICPC2ICD10ENG|X; histiocytosis, chronic|9754/3
C0019621|T191|PT|U002076|LCH|Hand-Schueller-Christian syndrome|9754/3
C0023381|T047|PT|U002660|LCH|Letterer-Siwe disease|9754/3
C0019621|T191|PT|sh85058638|LCH_NW|Hand-Schueller-Christian syndrome|9754/3
C0023381|T047|PT|sh85076237|LCH_NW|Letterer-Siwe disease|9754/3
C0019621|T191|LLT|10053133|MDR|Chronic idiopathic xanthomatosis|9754/3
C0019621|T191|LLT|10053135|MDR|Hand-Schueller-Christian disease|9754/3
C0019621|T191|LLT|10023688|MDR|Langerhans' cell granulomatosis|9754/3
C0019621|T191|LLT|10069698|MDR|Langerhans' cell histiocytosis|9754/3
C0019621|T191|PT|10069698|MDR|Langerhans' cell histiocytosis|9754/3
C0023381|T047|LLT|10024265|MDR|Letterer-Siwe disease|9754/3
C0019621|T191|SY|31815|MEDCIN|Hand-Schuller-Christian disease|9754/3
C0019621|T191|PT|315032|MEDCIN|Langerhans cell histiocytosis|9754/3
C0023381|T047|PT|31816|MEDCIN|Letterer-Siwe disease|9754/3
C0019621|T191|PT|31815|MEDCIN|multifocal eosinophilic granuloma|9754/3
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendothelioses, Systemic|9754/3
C0019621|T191|PM|D006646|MSH|Aleukemic Reticuloendotheliosis, Systemic|9754/3
C0019621|T191|PM|D006646|MSH|Cell Granulomatoses, Langerhans|9754/3
C0019621|T191|PM|D006646|MSH|Cell Granulomatosis, Langerhans|9754/3
C0019621|T191|PM|D006646|MSH|Cell Histiocytoses, Langerhans|9754/3
C0019621|T191|PM|D006646|MSH|Cell Histiocytosis, Langerhans|9754/3
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schueller-Christian|9754/3
C0019621|T191|PM|D006646|MSH|Disease, Hand-Schüller-Christian|9754/3
C0019621|T191|PM|D006646|MSH|Disease, Letterer-Siwe|9754/3
C0019621|T191|PM|D006646|MSH|Disease, Schueller-Christian|9754/3
C0023381|T047|NM|C538636|MSH|Familial Letterer-Siwe disease|9754/3
C0019621|T191|PM|D006646|MSH|Generalized Histiocytoses|9754/3
C0019621|T191|PM|D006646|MSH|Generalized Histiocytosis|9754/3
C0019621|T191|PM|D006646|MSH|Granulomatoses, Langerhans Cell|9754/3
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans Cell|9754/3
C0019621|T191|PM|D006646|MSH|Granulomatosis, Langerhans-Cell|9754/3
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Disease|9754/3
C0019621|T191|PM|D006646|MSH|Hand Schueller Christian Syndrome|9754/3
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Disease|9754/3
C0019621|T191|PM|D006646|MSH|Hand Schüller Christian Syndrome|9754/3
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Disease|9754/3
C0019621|T191|ET|D006646|MSH|Hand-Schueller-Christian Syndrome|9754/3
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Disease|9754/3
C0019621|T191|ET|D006646|MSH|Hand-Schüller-Christian Syndrome|9754/3
C0019621|T191|PM|D006646|MSH|Histiocytoses, Generalized|9754/3
C0019621|T191|PM|D006646|MSH|Histiocytoses, Langerhans Cell|9754/3
C0019621|T191|PM|D006646|MSH|Histiocytoses, Type 2|9754/3
C0019621|T191|ET|D006646|MSH|Histiocytosis X|9754/3
C0023381|T047|CE|C538636|MSH|Histiocytosis X, acute disseminated|9754/3
C0019621|T191|ET|D006646|MSH|Histiocytosis-X|9754/3
C0019621|T191|ET|D006646|MSH|Histiocytosis, Generalized|9754/3
C0019621|T191|PM|D006646|MSH|Histiocytosis, Langerhans Cell|9754/3
C0019621|T191|MH|D006646|MSH|Histiocytosis, Langerhans-Cell|9754/3
C0019621|T191|PM|D006646|MSH|Histiocytosis, Type 2|9754/3
C0019621|T191|PM|D006646|MSH|Langerhans Cell Granulomatoses|9754/3
C0019621|T191|ET|D006646|MSH|Langerhans Cell Granulomatosis|9754/3
C0019621|T191|PM|D006646|MSH|Langerhans Cell Histiocytoses|9754/3
C0019621|T191|ET|D006646|MSH|Langerhans Cell Histiocytosis|9754/3
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Granulomatosis|9754/3
C0019621|T191|ET|D006646|MSH|Langerhans-Cell Histiocytosis|9754/3
C0019621|T191|DEV|D006646|MSH|LETTERER SIWE DIS|9754/3
C0019621|T191|PM|D006646|MSH|Letterer Siwe Disease|9754/3
C0019621|T191|ET|D006646|MSH|Letterer-Siwe Disease|9754/3
C0019621|T191|PM|D006646|MSH|Non Lipid Reticuloendotheliosis|9754/3
C0019621|T191|PM|D006646|MSH|Non-Lipid Reticuloendothelioses|9754/3
C0019621|T191|ET|D006646|MSH|Non-Lipid Reticuloendotheliosis|9754/3
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Non-Lipid|9754/3
C0019621|T191|PM|D006646|MSH|Reticuloendothelioses, Systemic Aleukemic|9754/3
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Non-Lipid|9754/3
C0019621|T191|PM|D006646|MSH|Reticuloendotheliosis, Systemic Aleukemic|9754/3
C0019621|T191|DEV|D006646|MSH|SCHUELLER CHRISTIAN DIS|9754/3
C0019621|T191|PM|D006646|MSH|Schueller Christian Disease|9754/3
C0019621|T191|ET|D006646|MSH|Schueller-Christian Disease|9754/3
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schueller-Christian|9754/3
C0019621|T191|PM|D006646|MSH|Syndrome, Hand-Schüller-Christian|9754/3
C0019621|T191|PM|D006646|MSH|Systemic Aleukemic Reticuloendothelioses|9754/3
C0019621|T191|ET|D006646|MSH|Systemic Aleukemic Reticuloendotheliosis|9754/3
C0019621|T191|PM|D006646|MSH|Type 2 Histiocytoses|9754/3
C0019621|T191|ET|D006646|MSH|Type 2 Histiocytosis|9754/3
C0019621|T191|PN|NOCODE|MTH|Histiocytosis, Langerhans-Cell|9754/3
C0023381|T047|PN|NOCODE|MTH|Letterer-Siwe Disease|9754/3
C0023381|T047|ET|202.5|MTHICD9|Acute differentiated progressive histiocytosis|9754/3
C0023381|T047|ET|202.5|MTHICD9|Acute histiocytosis X|9754/3
C0023381|T047|ET|202.5|MTHICD9|Acute infantile reticuloendotheliosis|9754/3
C0023381|T047|ET|202.5|MTHICD9|Acute progressive histiocytosis X|9754/3
C0023381|T047|ET|202.5|MTHICD9|Acute reticulosis of infancy|9754/3
C0019621|T191|ET|277.89|MTHICD9|Chronic Histiocytosis X|9754/3
C0019621|T191|ET|277.89|MTHICD9|Hand-Schuller-Christian disease|9754/3
C0019621|T191|ET|277.89|MTHICD9|Histiocytosis X|9754/3
C0019621|T191|PT|C6920|NCI|Hand-Schuller-Christian Disease|9754/3
C0019621|T191|OP|C3107|NCI|Histiocytosis X|9754/3
C0019621|T191|SY|C3107|NCI|Langerhans Cell Granulomatosis|9754/3
C0019621|T191|SY|TCGA|NCI|Langerhans Cell Histiocytosis|9754/3
C0019621|T191|PT|C3107|NCI|Langerhans Cell Histiocytosis|9754/3
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, NOS|9754/3
C0019621|T191|SY|C3107|NCI|Langerhans Cell Histiocytosis, Not Otherwise Specified|9754/3
C0019621|T191|AB|C3107|NCI|LCH|9754/3
C0023381|T047|PT|C3160|NCI|Letterer-Siwe Disease|9754/3
C0019621|T191|PT|C6920|NCI_CPTAC|Hand-Schuller-Christian Disease|9754/3
C0023381|T047|PT|C3160|NCI_CPTAC|Letterer-Siwe Disease|9754/3
C0019621|T191|PT|10025581|NCI_CTEP-SDC|Langerhans cell histiocytosis|9754/3
C0019621|T191|DN|C3107|NCI_CTRP|Langerhans Cell Histiocytosis|9754/3
C0019621|T191|PT|CDR0000471787|NCI_NCI-GLOSS|Langerhans cell histiocytosis|9754/3
C0019621|T191|PT|CDR0000513054|NCI_NCI-GLOSS|LCH|9754/3
C0023381|T047|SY|C3160|NCI_NICHD|Acute Disseminated Langerhans Cell Histiocytosis|9754/3
C0019621|T191|SY|C6920|NCI_NICHD|Classic Multifocal Langerhans Cell Histiocytosis|9754/3
C0019621|T191|SY|C6920|NCI_NICHD|Hand-Schüller-Christian Disease|9754/3
C0019621|T191|OP|C3107|NCI_NICHD|Histiocytosis X|9754/3
C0019621|T191|PT|C3107|NCI_NICHD|Langerhans Cell Histiocytosis|9754/3
C0023381|T047|SY|C3160|NCI_NICHD|Letterer-Siwe Disease|9754/3
C0023381|T047|PT|C3160|NCI_NICHD|Multifocal Multisystem Langerhans Cell Histiocytosis|9754/3
C0019621|T191|PT|C6920|NCI_NICHD|Multifocal Unisystem Langerhans Cell Histiocytosis|9754/3
C0019621|T191|SY|CDR0000039054|PDQ|histiocytosis X|9754/3
C0019621|T191|PT|CDR0000641624|PDQ|Langerhans cell histiocytosis|9754/3
C0023381|T047|SY|B625.|RCD|Acute infancy reticulosis|9754/3
C0023381|T047|AB|B625.|RCD|Acute prog histiocytosis X|9754/3
C0023381|T047|SY|B625.|RCD|Acute progressive histiocytosis X|9754/3
C0019621|T191|AB|X20E9|RCD|Different progress histiocyto|9754/3
C0019621|T191|SY|X20E9|RCD|Differentiated progressive histiocytosis|9754/3
C0019621|T191|AB|C37y0|RCD|Hand-Schuller-Christian diseas|9754/3
C0019621|T191|SY|C37y0|RCD|Hand-Schuller-Christian disease|9754/3
C0023381|T047|SY|B625.|RCD|Histiocytosis X|9754/3
C0019621|T191|OP|C37y6|RCD|Histiocytosis X , unspecified|9754/3
C0019621|T191|PT|C37y5|RCD|Histiocytosis X syndrome|9754/3
C0019621|T191|PT|X20E9|RCD|Langerhan's cell histiocytosis|9754/3
C0019621|T191|AB|X20E9|RCD|Langerhans histiocyt syndrome|9754/3
C0019621|T191|SY|X20E9|RCD|Langerhans histiocytic syndrome|9754/3
C0019621|T191|SY|X20E9|RCD|LCH - Langerhan's cell histiocytosis|9754/3
C0019621|T191|AB|X20E9|RCD|LCH-Langerh cell histiocytosis|9754/3
C0023381|T047|OA|B6250|RCD|Letterer-Siwe dis.-unspec.site|9754/3
C0023381|T047|PT|B625.|RCD|Letterer-Siwe disease|9754/3
C0023381|T047|OP|B625z|RCD|Letterer-Siwe disease NOS|9754/3
C0023381|T047|OP|B6250|RCD|Letterer-Siwe disease of unspecified sites|9754/3
C0023381|T047|SY|B625.|RCD|LSD - Letterer-Siwe disease|9754/3
C0019621|T191|PT|C37y0|RCD|Schuller-Christian syndrome|9754/3
C0023381|T047|IS|BBm3.|RCDSY|Acute infancy reticulosis|9754/3
C0023381|T047|OA|BBm3.|RCDSY|Acute progress histiocyt X|9754/3
C0023381|T047|IS|BBm3.|RCDSY|Acute progressive histiocytosis X|9754/3
C0023381|T047|OP|BBm3.|RCDSY|Letterer - Siwe disease|9754/3
C0023381|T047|IS|67574008|SNOMEDCT_US|Acute differentiated progressive histiocytosis|9754/3
C0023381|T047|SY|118614007|SNOMEDCT_US|Acute infancy reticulosis|9754/3
C0023381|T047|OAS|366059005|SNOMEDCT_US|Acute infancy reticulosis|9754/3
C0023381|T047|SY|128812005|SNOMEDCT_US|Acute infancy reticulosis|9754/3
C0023381|T047|OAS|366059005|SNOMEDCT_US|Acute progressive histiocytosis X|9754/3
C0023381|T047|SY|118614007|SNOMEDCT_US|Acute progressive histiocytosis X|9754/3
C0023381|T047|IS|128812005|SNOMEDCT_US|Acute progressive histiocytosis X|9754/3
C0023381|T047|IS|67574008|SNOMEDCT_US|Acute progressive histiocytosis X|9754/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic differentiated progressive histiocytosis|9754/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic disseminated histiocytosis X|9754/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic histiocytosis X|9754/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Chronic idiopathic xanthomatosis|9754/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|Differentiated progressive histiocytosis|9754/3
C0019621|T191|SY|65399007|SNOMEDCT_US|Differentiated progressive histiocytosis|9754/3
C0019621|T191|SYGB|39795003|SNOMEDCT_US|Generalised histiocytosis of bones|9754/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Generalized histiocytosis of bones|9754/3
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand - Schuller - Christian disease|9754/3
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand - Schuller - Christian disease|9754/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Hand-Schuller-Christian disease|9754/3
C0019621|T191|PT|39795003|SNOMEDCT_US|Hand-Schüller-Christian disease|9754/3
C0019621|T191|OAS|267510005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9754/3
C0019621|T191|OAS|154773005|SNOMEDCT_US|Hand-Schuller-Christian syndr.|9754/3
C0019621|T191|SY|65399007|SNOMEDCT_US|Histiocytosis X|9754/3
C0019621|T191|OAS|154583006|SNOMEDCT_US|Histiocytosis X|9754/3
C0019621|T191|OAS|269628007|SNOMEDCT_US|Histiocytosis X|9754/3
C0019621|T191|IS|190960001|SNOMEDCT_US|Histiocytosis X , chronic|9754/3
C0019621|T191|IS|190956004|SNOMEDCT_US|Histiocytosis X , unspecified|9754/3
C0019621|T191|PT|190955000|SNOMEDCT_US|Histiocytosis X syndrome|9754/3
C0019621|T191|IS|65399007|SNOMEDCT_US|Histiocytosis X, NOS|9754/3
C0019621|T191|OAP|190956004|SNOMEDCT_US|Histiocytosis X, unspecified|9754/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhan's cell histiocytosis|9754/3
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhan's cell histiocytosis|9754/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans cell disease|9754/3
C0019621|T191|SY|65399007|SNOMEDCT_US|Langerhans cell disease|9754/3
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9754/3
C0019621|T191|IS|128809007|SNOMEDCT_US|Langerhans cell granulomatosis|9754/3
C0019621|T191|PT|65399007|SNOMEDCT_US|Langerhans cell histiocytosis|9754/3
C0019621|T191|PT|128809007|SNOMEDCT_US|Langerhans cell histiocytosis|9754/3
C0019621|T191|OAP|234439008|SNOMEDCT_US|Langerhans cell histiocytosis|9754/3
C0023381|T047|PT|128812005|SNOMEDCT_US|Langerhans cell histiocytosis, disseminated|9754/3
C0023381|T047|SY|118614007|SNOMEDCT_US|Langerhans cell histiocytosis, disseminated|9754/3
C0023381|T047|SYGB|128812005|SNOMEDCT_US|Langerhans cell histiocytosis, generalised|9754/3
C0023381|T047|SY|128812005|SNOMEDCT_US|Langerhans cell histiocytosis, generalized|9754/3
C0019621|T191|PT|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, multifocal|9754/3
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no ICD-O subtype|9754/3
C0019621|T191|SY|128809007|SNOMEDCT_US|Langerhans cell histiocytosis, no International Classification of Diseases for Oncology subtype|9754/3
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, poly-ostotic|9754/3
C0019621|T191|SY|128811003|SNOMEDCT_US|Langerhans cell histiocytosis, polyostotic|9754/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|Langerhans histiocytic syndrome|9754/3
C0019621|T191|OAP|110450007|SNOMEDCT_US|Langerhans' cell histiocytosis|9754/3
C0019621|T191|OAS|234439008|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9754/3
C0019621|T191|SY|65399007|SNOMEDCT_US|LCH - Langerhan's cell histiocytosis|9754/3
C0023381|T047|OAP|188654004|SNOMEDCT_US|Letterer-Siwe disease|9754/3
C0023381|T047|OAP|366059005|SNOMEDCT_US|Letterer-Siwe disease|9754/3
C0023381|T047|OAS|154583006|SNOMEDCT_US|Letterer-Siwe disease|9754/3
C0023381|T047|OAS|269628007|SNOMEDCT_US|Letterer-Siwe disease|9754/3
C0023381|T047|SY|128812005|SNOMEDCT_US|Letterer-Siwe disease|9754/3
C0023381|T047|OAP|188659009|SNOMEDCT_US|Letterer-Siwe disease NOS|9754/3
C0023381|T047|OAP|188655003|SNOMEDCT_US|Letterer-Siwe disease of unspecified sites|9754/3
C0023381|T047|OAP|67574008|SNOMEDCT_US|Letterer-Siwe's disease|9754/3
C0023381|T047|IS|67574008|SNOMEDCT_US|Letterer-Siwe's disease -RETIRED-|9754/3
C0023381|T047|OF|67574008|SNOMEDCT_US|Letterer-Siwe's disease -RETIRED-|9754/3
C0023381|T047|SY|118614007|SNOMEDCT_US|LSD - Letterer-Siwe disease|9754/3
C0023381|T047|OAS|366059005|SNOMEDCT_US|LSD - Letterer-Siwe disease|9754/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Multifocal and unisystemic Langerhans cell histiocytosis|9754/3
C0023381|T047|IS|67574008|SNOMEDCT_US|Nonlipid reticuloendotheliosis|9754/3
C0019621|T191|SY|39795003|SNOMEDCT_US|Schuller-Christian syndrome|9754/3
C0334663|T191|PT|0000030018|CHV|histiocytic sarcoma|9755/3
C0334663|T191|PT|C96.3|ICD10|True histiocytic lymphoma|9755/3
C0334663|T191|PT|C96.A|ICD10CM|Histiocytic sarcoma|9755/3
C0334663|T191|AB|C96.A|ICD10CM|Histiocytic sarcoma|9755/3
C0334663|T191|PT|MTHU035167|ICPC2ICD10ENG|histiocytic; lymphoma, true|9755/3
C0334663|T191|PT|MTHU046801|ICPC2ICD10ENG|lymphoma; histiocytic, true|9755/3
C0334663|T191|PT|MTHU046769|ICPC2ICD10ENG|lymphoma; true histiocytic|9755/3
C0334663|T191|PT|MTHU024682|ICPC2ICD10ENG|true histiocytic; lymphoma|9755/3
C0334663|T191|PT|10076876|MDR|Histiocytic sarcoma|9755/3
C0334663|T191|LLT|10076876|MDR|Histiocytic sarcoma|9755/3
C0334663|T191|PT|272060|MEDCIN|histiocytic sarcoma|9755/3
C0334663|T191|PM|D054747|MSH|Histiocytic Lymphoma, True|9755/3
C0334663|T191|PM|D054747|MSH|Histiocytic Lymphomas, True|9755/3
C0334663|T191|MH|D054747|MSH|Histiocytic Sarcoma|9755/3
C0334663|T191|PM|D054747|MSH|Histiocytic Sarcomas|9755/3
C0334663|T191|PM|D054747|MSH|Histiocytoses, True Malignant|9755/3
C0334663|T191|PM|D054747|MSH|Histiocytosis, True Malignant|9755/3
C0334663|T191|PM|D054747|MSH|Lymphoma, True Histiocytic|9755/3
C0334663|T191|PM|D054747|MSH|Lymphomas, True Histiocytic|9755/3
C0334663|T191|PM|D054747|MSH|Malignant Histiocytoses, True|9755/3
C0334663|T191|PM|D054747|MSH|Malignant Histiocytosis, True|9755/3
C0334663|T191|PM|D054747|MSH|Sarcoma, Histiocytic|9755/3
C0334663|T191|PM|D054747|MSH|Sarcomas, Histiocytic|9755/3
C0334663|T191|ET|D054747|MSH|True Histiocytic Lymphoma|9755/3
C0334663|T191|PM|D054747|MSH|True Histiocytic Lymphomas|9755/3
C0334663|T191|PM|D054747|MSH|True Malignant Histiocytoses|9755/3
C0334663|T191|ET|D054747|MSH|True Malignant Histiocytosis|9755/3
C0334663|T191|PN|NOCODE|MTH|Histiocytic sarcoma|9755/3
C0334663|T191|SY|TCGA|NCI|Histiocytic Sarcoma|9755/3
C0334663|T191|PT|C27349|NCI|Histiocytic Sarcoma|9755/3
C0334663|T191|OP|C35382|NCI|True Histiocytic Lymphoma|9755/3
C0334663|T191|PT|C35382|NCI|True Histiocytic Lymphoma|9755/3
C0334663|T191|PT|C27349|NCI_CDISC|SARCOMA, HISTIOCYTIC, MALIGNANT|9755/3
C0334663|T191|PT|C27349|NCI_CPTAC|Histiocytic Sarcoma|9755/3
C0334663|T191|PT|CDR0000373019|NCI_NCI-GLOSS|histiocytic lymphoma|9755/3
C0334663|T191|PT|CDR0000776971|PDQ|histiocytic sarcoma|9755/3
C0334663|T191|PT|Xa0Ty|RCD|True histiocytic lymphoma|9755/3
C0334663|T191|OP|BBm4.|RCDSY|True histiocytic lymphoma|9755/3
C0334663|T191|SY|109988003|SNOMEDCT_US|Histiocytic sarcoma|9755/3
C0334663|T191|PT|128813000|SNOMEDCT_US|Histiocytic sarcoma|9755/3
C0334663|T191|OAP|26640009|SNOMEDCT_US|True histiocytic lymphoma|9755/3
C0334663|T191|SY|128813000|SNOMEDCT_US|True histiocytic lymphoma|9755/3
C0334663|T191|OAP|188692003|SNOMEDCT_US|True histiocytic lymphoma|9755/3
C0334663|T191|SY|109988003|SNOMEDCT_US|True histiocytic lymphoma|9755/3
C0334663|T191|OF|188692003|SNOMEDCT_US|True histiocytic lymphoma|9755/3
C0334663|T191|OF|26640009|SNOMEDCT_US|True histiocytic lymphoma -RETIRED-|9755/3
C0334663|T191|IS|26640009|SNOMEDCT_US|True histiocytic lymphoma -RETIRED-|9755/3
C1260327|T191|ET|C96.4|ICD10CM|Langerhans cell sarcoma|9756/3
C1260327|T191|LLT|10078782|MDR|Langerhans cell sarcoma|9756/3
C1260327|T191|PT|10078782|MDR|Langerhans cell sarcoma|9756/3
C1260327|T191|PT|391486|MEDCIN|Langerhans cell sarcoma|9756/3
C1260327|T191|SY|391486|MEDCIN|sarcoma Langerhans cell|9756/3
C1260327|T191|MH|D054752|MSH|Langerhans Cell Sarcoma|9756/3
C1260327|T191|PM|D054752|MSH|Langerhans Cell Sarcomas|9756/3
C1260327|T191|PM|D054752|MSH|Sarcoma, Langerhans Cell|9756/3
C1260327|T191|PM|D054752|MSH|Sarcomas, Langerhans Cell|9756/3
C1260327|T191|ET|202.9|MTHICD9|Langerhans cell sarcoma|9756/3
C1260327|T191|SY|TCGA|NCI|Langerhans Cell Sarcoma|9756/3
C1260327|T191|PT|C6921|NCI|Langerhans Cell Sarcoma|9756/3
C1260327|T191|PT|C6921|NCI_CPTAC|Langerhans Cell Sarcoma|9756/3
C1260327|T191|PT|128814006|SNOMEDCT_US|Langerhans cell sarcoma|9756/3
C1260327|T191|PT|724649000|SNOMEDCT_US|Langerhans cell sarcoma|9756/3
C1260326|T191|PT|0000056321|CHV|dendritic cell sarcoma|9757/1
C1260326|T191|ET|C96.4|ICD10CM|Interdigitating dendritic cell sarcoma|9757/1
C1260326|T191|PT|272062|MEDCIN|interdigitating dendritic cell sarcoma|9757/1
C1260326|T191|MH|D054739|MSH|Dendritic Cell Sarcoma, Interdigitating|9757/1
C1260326|T191|ET|D054739|MSH|Interdigitating Cell Sarcoma|9757/1
C1260326|T191|PM|D054739|MSH|Interdigitating Cell Sarcomas|9757/1
C1260326|T191|ET|D054739|MSH|Interdigitating Dendritic Cell Sarcoma|9757/1
C1260326|T191|PM|D054739|MSH|Sarcoma, Interdigitating Cell|9757/1
C1260326|T191|PM|D054739|MSH|Sarcomas, Interdigitating Cell|9757/1
C1260326|T191|PN|NOCODE|MTH|Dendritic Cell Sarcoma, Interdigitating|9757/1
C1260326|T191|ET|202.9|MTHICD9|Interdigitating dendritic cell sarcoma|9757/1
C1260326|T191|SY|C9282|NCI|Interdigitating Cell Sarcoma/Tumor|9757/1
C1260326|T191|SY|TCGA|NCI|Interdigitating Dendritic Cell Sarcoma|9757/1
C1260326|T191|PT|C9282|NCI|Interdigitating Dendritic Cell Sarcoma|9757/1
C1260326|T191|SY|C9282|NCI|Interdigitating Dendritic Cell Sarcoma/Tumor|9757/1
C1260326|T191|PT|C9282|NCI_CPTAC|Interdigitating Dendritic Cell Sarcoma|9757/1
C1260326|T191|SY|128815007|SNOMEDCT_US|Interdigitating cell sarcoma|9757/1
C1260326|T191|PT|128815007|SNOMEDCT_US|Interdigitating dendritic cell sarcoma|9757/1
C1260326|T191|PT|0000056321|CHV|dendritic cell sarcoma|9757/3
C1260326|T191|ET|C96.4|ICD10CM|Interdigitating dendritic cell sarcoma|9757/3
C2825741|T191|SY|366682|MEDCIN|histiocytic dis interdigitating dendritic cell indeterminate neoplasm|9757/3
C2825741|T191|PT|366682|MEDCIN|Indeterminate dendritic cell neoplasm|9757/3
C1260326|T191|PT|272062|MEDCIN|interdigitating dendritic cell sarcoma|9757/3
C1301364|T191|PT|338577|MEDCIN|sarcoma of dendritic cell|9757/3
C1260326|T191|MH|D054739|MSH|Dendritic Cell Sarcoma, Interdigitating|9757/3
C1260326|T191|ET|D054739|MSH|Interdigitating Cell Sarcoma|9757/3
C1260326|T191|PM|D054739|MSH|Interdigitating Cell Sarcomas|9757/3
C1260326|T191|ET|D054739|MSH|Interdigitating Dendritic Cell Sarcoma|9757/3
C1260326|T191|PM|D054739|MSH|Sarcoma, Interdigitating Cell|9757/3
C1260326|T191|PM|D054739|MSH|Sarcomas, Interdigitating Cell|9757/3
C1260326|T191|PN|NOCODE|MTH|Dendritic Cell Sarcoma, Interdigitating|9757/3
C1301364|T191|PN|NOCODE|MTH|Dendritic cell sarcoma, not otherwise specified|9757/3
C1260326|T191|ET|202.9|MTHICD9|Interdigitating dendritic cell sarcoma|9757/3
C1301364|T191|OP|C27260|NCI|Dendritic Cell Sarcoma, NOS|9757/3
C1301364|T191|PT|C27260|NCI|Dendritic Cell Tumor, Not Otherwise Specified|9757/3
C1301364|T191|SY|TCGA|NCI|Dendritic Cell Tumor, Not Otherwise Specified|9757/3
C1301364|T191|OP|C27260|NCI|Dendritic Cell Tumor, Not Otherwise Specified|9757/3
C2825741|T191|SY|C81767|NCI|Indeterminate Cell Histiocytosis|9757/3
C2825741|T191|PT|C81767|NCI|Indeterminate Dendritic Cell Tumor|9757/3
C1260326|T191|SY|C9282|NCI|Interdigitating Cell Sarcoma/Tumor|9757/3
C1260326|T191|PT|C9282|NCI|Interdigitating Dendritic Cell Sarcoma|9757/3
C1260326|T191|SY|TCGA|NCI|Interdigitating Dendritic Cell Sarcoma|9757/3
C1260326|T191|SY|C9282|NCI|Interdigitating Dendritic Cell Sarcoma/Tumor|9757/3
C1260326|T191|PT|C9282|NCI_CPTAC|Interdigitating Dendritic Cell Sarcoma|9757/3
C1301364|T191|IS|128815007|SNOMEDCT_US|Dendritic cell sarcoma|9757/3
C1301364|T191|SY|397355008|SNOMEDCT_US|Dendritic cell sarcoma, no ICD-O subtype|9757/3
C1301364|T191|PT|397355008|SNOMEDCT_US|Dendritic cell sarcoma, no International Classification of Diseases for Oncology subtype|9757/3
C1301364|T191|OP|397355008|SNOMEDCT_US|Dendritic cell sarcoma, not otherwise specified|9757/3
C2825741|T191|PT|721313009|SNOMEDCT_US|Indeterminate dendritic cell neoplasm|9757/3
C2825741|T191|PT|703822002|SNOMEDCT_US|Indeterminate dendritic cell tumor|9757/3
C2825741|T191|SY|721313009|SNOMEDCT_US|Indeterminate dendritic cell tumor|9757/3
C2825741|T191|PTGB|703822002|SNOMEDCT_US|Indeterminate dendritic cell tumour|9757/3
C2825741|T191|SYGB|721313009|SNOMEDCT_US|Indeterminate dendritic cell tumour|9757/3
C1260326|T191|SY|128815007|SNOMEDCT_US|Interdigitating cell sarcoma|9757/3
C1260326|T191|PT|128815007|SNOMEDCT_US|Interdigitating dendritic cell sarcoma|9757/3
C1260325|T191|ET|C96.4|ICD10CM|Follicular dendritic cell sarcoma|9758/1
C1260325|T191|LLT|10075332|MDR|Follicular dendritic cell sarcoma|9758/1
C1260325|T191|PT|10075332|MDR|Follicular dendritic cell sarcoma|9758/1
C1260325|T191|PT|272063|MEDCIN|follicular dendritic cell sarcoma|9758/1
C1260325|T191|MH|D054740|MSH|Dendritic Cell Sarcoma, Follicular|9758/1
C1260325|T191|ET|D054740|MSH|Follicular Dendritic Cell Sarcoma|9758/1
C1260325|T191|ET|202.9|MTHICD9|Follicular dendritic cell sarcoma|9758/1
C1260325|T191|SY|TCGA|NCI|Follicular Dendritic Cell Sarcoma|9758/1
C1260325|T191|PT|C9281|NCI|Follicular Dendritic Cell Sarcoma|9758/1
C1260325|T191|SY|C9281|NCI|Follicular Dendritic Cell Sarcoma/Tumor|9758/1
C1260325|T191|PT|C9281|NCI_CPTAC|Follicular Dendritic Cell Sarcoma|9758/1
C1260325|T191|PT|128816008|SNOMEDCT_US|Follicular dendritic cell sarcoma|9758/1
C1260325|T191|SY|128816008|SNOMEDCT_US|Follicular dendritic cell tumor|9758/1
C1260325|T191|SYGB|128816008|SNOMEDCT_US|Follicular dendritic cell tumour|9758/1
C1260325|T191|ET|C96.4|ICD10CM|Follicular dendritic cell sarcoma|9758/3
C1260325|T191|LLT|10075332|MDR|Follicular dendritic cell sarcoma|9758/3
C1260325|T191|PT|10075332|MDR|Follicular dendritic cell sarcoma|9758/3
C1260325|T191|PT|272063|MEDCIN|follicular dendritic cell sarcoma|9758/3
C1260325|T191|MH|D054740|MSH|Dendritic Cell Sarcoma, Follicular|9758/3
C1260325|T191|ET|D054740|MSH|Follicular Dendritic Cell Sarcoma|9758/3
C1260325|T191|ET|202.9|MTHICD9|Follicular dendritic cell sarcoma|9758/3
C1260325|T191|SY|TCGA|NCI|Follicular Dendritic Cell Sarcoma|9758/3
C1260325|T191|PT|C9281|NCI|Follicular Dendritic Cell Sarcoma|9758/3
C1260325|T191|SY|C9281|NCI|Follicular Dendritic Cell Sarcoma/Tumor|9758/3
C1260325|T191|PT|C9281|NCI_CPTAC|Follicular Dendritic Cell Sarcoma|9758/3
C1260325|T191|PT|128816008|SNOMEDCT_US|Follicular dendritic cell sarcoma|9758/3
C1260325|T191|SY|128816008|SNOMEDCT_US|Follicular dendritic cell tumor|9758/3
C1260325|T191|SYGB|128816008|SNOMEDCT_US|Follicular dendritic cell tumour|9758/3
C2825739|T191|PT|366680|MEDCIN|Fibroblastic reticular cell neoplasm|9759/3
C2825739|T191|SY|366680|MEDCIN|malig neoplasm histiocytic disorder fibroblastic reticular cell neoplasm|9759/3
C2825739|T191|PT|C81758|NCI|Fibroblastic Reticular Cell Tumor|9759/3
C2825739|T191|PT|C81758|NCI_CPTAC|Fibroblastic Reticular Cell Tumor|9759/3
C2825739|T191|PT|721314003|SNOMEDCT_US|Fibroblastic reticular cell neoplasm|9759/3
C2825739|T191|PT|450912008|SNOMEDCT_US|Fibroblastic reticular cell tumor|9759/3
C2825739|T191|SY|721314003|SNOMEDCT_US|Fibroblastic reticular cell tumor|9759/3
C2825739|T191|PTGB|450912008|SNOMEDCT_US|Fibroblastic reticular cell tumour|9759/3
C2825739|T191|SYGB|721314003|SNOMEDCT_US|Fibroblastic reticular cell tumour|9759/3
C0021071|T191|SY|0000006611|CHV|alpha-chain disease|9760/3
C0021071|T191|SY|0000006611|CHV|chain alpha disease|9760/3
C0021070|T191|PT|0000006610|CHV|immunoproliferative disease|9760/3
C0021071|T191|PT|0000006611|CHV|ipsid|9760/3
C0021071|T191|SY|NOCODE|DXP|ALPHA CHAIN DISEASE|9760/3
C0021071|T191|SY|NOCODE|DXP|ALPHA HCD|9760/3
C0021071|T191|SY|NOCODE|DXP|ALPHA HEAVY CHAIN DISEASE|9760/3
C0021071|T191|SY|NOCODE|DXP|ALPHA-HEAVY CHAIN DISEASE|9760/3
C0021071|T191|SY|NOCODE|DXP|IGA HEAVY CHAIN DISEASE|9760/3
C0021071|T191|SY|NOCODE|DXP|IMMUNOPROLIFERATIVE SMALL INTESTINE DISEASE|9760/3
C0021071|T191|SY|NOCODE|DXP|IPSID|9760/3
C0021071|T191|ET|HP:0020194|HPO|Alpha heavy chain disease|9760/3
C0021071|T191|PT|C88.1|ICD10|Alpha heavy chain disease|9760/3
C0021071|T191|PT|C88.3|ICD10|Immunoproliferative small intestinal disease|9760/3
C0021071|T191|ET|C88.3|ICD10CM|Alpha heavy chain disease|9760/3
C0021070|T191|ET|C88.9|ICD10CM|Immunoproliferative disease NOS|9760/3
C0021071|T191|AB|C88.3|ICD10CM|Immunoproliferative small intestinal disease|9760/3
C0021071|T191|PT|C88.3|ICD10CM|Immunoproliferative small intestinal disease|9760/3
C0021071|T191|ET|C88.3|ICD10CM|Mediterranean lymphoma|9760/3
C0021071|T191|PT|MTHU005087|ICPC2ICD10ENG|alpha heavy chain; disease|9760/3
C0021071|T191|PT|MTHU004932|ICPC2ICD10ENG|alpha; alpha heavy chain disease|9760/3
C0021071|T191|PT|MTHU023293|ICPC2ICD10ENG|disease; alpha heavy chain|9760/3
C0021071|T191|PT|MTHU033693|ICPC2ICD10ENG|heavy chain alpha|9760/3
C0021070|T191|PT|MTHU090249|ICPC2ICD10ENG|immunoproliferative; disease|9760/3
C0021071|T191|PT|MTHU090250|ICPC2ICD10ENG|immunoproliferative; disease, small intestine|9760/3
C0021071|T191|PT|MTHU046826|ICPC2ICD10ENG|lymphoma; mediterranean|9760/3
C0021071|T191|PT|MTHU049176|ICPC2ICD10ENG|mediterranean; lymphoma|9760/3
C0021071|T191|PT|351185|MEDCIN|Alpha heavy chain disease|9760/3
C0021071|T191|PT|351186|MEDCIN|Alpha heavy chain disease, enteric form|9760/3
C0021071|T191|SY|351185|MEDCIN|heavy chain disease alpha|9760/3
C0021071|T191|SY|351186|MEDCIN|heavy chain disease alpha, enteric form|9760/3
C0021071|T191|SY|31572|MEDCIN|immunoproliferative intestinal disease|9760/3
C0021071|T191|PT|31572|MEDCIN|immunoproliferative small intestinal disease|9760/3
C0021071|T191|DEV|D007161|MSH|ALPHA CHAIN DIS|9760/3
C0021071|T191|PM|D007161|MSH|alpha Chain Disease|9760/3
C0021071|T191|ET|D007161|MSH|alpha-Chain Disease|9760/3
C0021071|T191|PM|D007161|MSH|alpha-Chain Diseases|9760/3
C0021071|T191|PM|D007161|MSH|Disease, alpha-Chain|9760/3
C0021071|T191|PM|D007161|MSH|Diseases, alpha-Chain|9760/3
C0021070|T191|PM|D007160|MSH|Disorder, Immunoproliferative|9760/3
C0021070|T191|PM|D007160|MSH|Disorders, Immunoproliferative|9760/3
C0021071|T191|DEV|D007161|MSH|HEAVY CHAIN DIS IGA TYPE|9760/3
C0021071|T191|ET|D007161|MSH|Heavy Chain Disease, IgA Type|9760/3
C0021070|T191|DEV|D007160|MSH|IMMUNOPROLIFERATIVE DIS|9760/3
C0021070|T191|PM|D007160|MSH|Immunoproliferative Disorder|9760/3
C0021070|T191|MH|D007160|MSH|Immunoproliferative Disorders|9760/3
C0021071|T191|DEV|D007161|MSH|IMMUNOPROLIFERATIVE SMALL INTESTINAL DIS|9760/3
C0021071|T191|MH|D007161|MSH|Immunoproliferative Small Intestinal Disease|9760/3
C0021071|T191|ET|D007161|MSH|IPSID|9760/3
C0021071|T191|ET|D007161|MSH|Lymphoma, Mediterranean|9760/3
C0021071|T191|PM|D007161|MSH|Mediterranean Lymphoma|9760/3
C0021071|T191|PT|C3132|NCI|Alpha Heavy Chain Disease|9760/3
C0021071|T191|SY|C3132|NCI|Immunoproliferative Small Intestinal Disease|9760/3
C0021071|T191|AB|C3132|NCI|IPSID|9760/3
C0021071|T191|SY|C3132|NCI|Mediterranean Abdominal Lymphoma|9760/3
C0021071|T191|SY|C3132|NCI|Mediterranean Lymphoma|9760/3
C0021071|T191|OP|C3331|RCD|Alpha heavy chain disease|9760/3
C0021071|T191|OP|BBm6.|RCDSY|Alpha heavy chain disease|9760/3
C0021071|T191|OP|BBmG.|RCDSY|Immunoproliferative small intestinal disease|9760/3
C0021071|T191|OA|BBmG.|RCDSY|Imunoprolif smal intest dis|9760/3
C0021071|T191|SY|109982002|SNOMEDCT_US|Alpha heavy chain disease|9760/3
C0021071|T191|OAP|190819007|SNOMEDCT_US|Alpha heavy chain disease|9760/3
C0021071|T191|SY|6381009|SNOMEDCT_US|Alpha heavy chain disease|9760/3
C0021071|T191|OAP|123312002|SNOMEDCT_US|Alpha heavy chain disease|9760/3
C0021071|T191|IS|123312002|SNOMEDCT_US|Alpha heavy chain disease -RETIRED-|9760/3
C0021071|T191|OF|123312002|SNOMEDCT_US|Alpha heavy chain disease -RETIRED-|9760/3
C0021071|T191|PT|123313007|SNOMEDCT_US|Alpha heavy chain disease, enteric form|9760/3
C0021071|T191|SY|27461004|SNOMEDCT_US|Alpha heavy chain disease, enteric form|9760/3
C0021071|T191|IS|123312002|SNOMEDCT_US|Alpha heavy chain disease, NOS|9760/3
C0021071|T191|SY|6381009|SNOMEDCT_US|IgA heavy chain disease|9760/3
C0021071|T191|IS|6381009|SNOMEDCT_US|IgA heavy chain disease, NOS|9760/3
C0021071|T191|IS|123312002|SNOMEDCT_US|IgA heavy chain disease, NOS|9760/3
C0021070|T191|PT|86295000|SNOMEDCT_US|Immunoproliferative disease|9760/3
C0021070|T191|OAP|134363002|SNOMEDCT_US|Immunoproliferative disease - morphology|9760/3
C0021070|T191|SY|86295000|SNOMEDCT_US|Immunoproliferative disease, no ICD-O subtype|9760/3
C0021070|T191|SY|86295000|SNOMEDCT_US|Immunoproliferative disease, no International Classification of Diseases for Oncology subtype|9760/3
C0021070|T191|IS|86295000|SNOMEDCT_US|Immunoproliferative disease, NOS|9760/3
C0021070|T191|PT|127071007|SNOMEDCT_US|Immunoproliferative disorder|9760/3
C0021071|T191|SY|109985000|SNOMEDCT_US|Immunoproliferative small intestinal disease|9760/3
C0021071|T191|IS|123313007|SNOMEDCT_US|Immunoproliferative small intestinal disease|9760/3
C0021071|T191|PT|27461004|SNOMEDCT_US|Immunoproliferative small intestinal disease|9760/3
C1532005|T191|PT|414646000|SNOMEDCT_US|Malignant immunoproliferative neoplasm|9760/3
C0021071|T191|IS|123313007|SNOMEDCT_US|Mediterranean lymphoma|9760/3
C0021071|T191|SY|27461004|SNOMEDCT_US|Mediterranean lymphoma|9760/3
C0024419|T191|ET|0000005754|AOD|macroglobulinemia|9761/3
C0334633|T191|PT|0000030014|CHV|immunocytoma|9761/3
C0024419|T191|SY|0000007643|CHV|lymphoplasmacytic lymphoma|9761/3
C0024419|T191|SY|0000007643|CHV|lymphoplasmacytoid lymphoma|9761/3
C0024419|T191|SY|0000007643|CHV|macroglobulinaemia|9761/3
C0024419|T191|PT|0000007643|CHV|macroglobulinemia|9761/3
C0024419|T191|SY|0000007643|CHV|macroglobulinemia waldenstrom|9761/3
C0024419|T191|SY|0000007643|CHV|macroglobulinemia waldenstrom's|9761/3
C0024419|T191|SY|0000007643|CHV|macroglobulinemia waldenstroms|9761/3
C0024419|T191|SY|0000007643|CHV|waldenstrom macroglobulinemia|9761/3
C0024419|T191|SY|0000007643|CHV|waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|SY|0000007643|CHV|waldenstrom's macroglobulinemia|9761/3
C0024419|T191|SY|0000007643|CHV|waldenstroms macroglobulinemia|9761/3
C0024419|T191|PT|NOCODE|COSTAR|Macroglobulinemia|9761/3
C0024419|T191|ET|0449-2705|CSP|macroglobulinemia|9761/3
C0024419|T191|ET|0449-8115|CSP|macroglobulinemia|9761/3
C0024419|T191|PT|0449-8115|CSP|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|DI|U001123|DXP|MACROGLOBULINEMIA, WALDENSTROM|9761/3
C0024419|T191|ET|HP:0005508|HPO|Waldenstrom macroglobulinemia|9761/3
C0024419|T191|PT|C88.0|ICD10|Waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|PT|C88.0|ICD10AE|Waldenstrom's macroglobulinemia|9761/3
C0334633|T191|ET|C83.0|ICD10CM|Lymphoplasmacytic lymphoma|9761/3
C0024419|T191|PT|C88.0|ICD10CM|Waldenström macroglobulinemia|9761/3
C0024419|T191|AB|C88.0|ICD10CM|Waldenstrom macroglobulinemia|9761/3
C0024419|T191|AB|273.3|ICD9CM|Macroglobulinemia|9761/3
C0024419|T191|PT|273.3|ICD9CM|Macroglobulinemia|9761/3
C0334633|T191|PT|MTHU037619|ICPC2ICD10ENG|immunocytoma|9761/3
C0334633|T191|PT|MTHU046823|ICPC2ICD10ENG|lymphoma; lymphoplasmacytoid|9761/3
C0334633|T191|PT|MTHU046851|ICPC2ICD10ENG|lymphoma; plasmacytic|9761/3
C0334633|T191|PT|MTHU046868|ICPC2ICD10ENG|lymphoplasmacytoid; lymphoma|9761/3
C0024419|T191|PT|MTHU047061|ICPC2ICD10ENG|macroglobulinemia|9761/3
C0024419|T191|PT|MTHU047062|ICPC2ICD10ENG|macroglobulinemia; Waldenström|9761/3
C0334633|T191|PT|MTHU059930|ICPC2ICD10ENG|plasmacytic; lymphoma|9761/3
C0024419|T191|PT|MTHU082024|ICPC2ICD10ENG|Waldenström; macroglobulinemia|9761/3
C0024419|T191|LLT|10062831|MDR|Macroglobulinaemia|9761/3
C0024419|T191|LLT|10025389|MDR|Macroglobulinaemia NOS|9761/3
C0024419|T191|LLT|10025390|MDR|Macroglobulinemia|9761/3
C0024419|T191|MTH_LLT|10025389|MDR|Macroglobulinemia NOS|9761/3
C0024419|T191|LLT|10081215|MDR|Primary macroglobulinaemia|9761/3
C0024419|T191|LLT|10081211|MDR|Primary macroglobulinemia|9761/3
C0024419|T191|LLT|10047714|MDR|Von Waldenstrom macroglobulinaemia|9761/3
C0024419|T191|LLT|10054693|MDR|Von Waldenstrom macroglobulinemia|9761/3
C0024419|T191|PT|10047801|MDR|Waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|LLT|10047801|MDR|Waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|LLT|10047803|MDR|Waldenstrom's macroglobulinaemia NOS|9761/3
C0024419|T191|HT|10047802|MDR|Waldenstrom's macroglobulinaemias|9761/3
C0024419|T191|LLT|10054695|MDR|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|MTH_PT|10047801|MDR|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|LLT|10054696|MDR|Waldenstrom's macroglobulinemia NOS|9761/3
C0334633|T191|PT|355928|MEDCIN|malignant lymphoplasmacytic lymphoma|9761/3
C0334633|T191|SY|355928|MEDCIN|malignant neoplasm lymphoma lymphoplasmacytic|9761/3
C0024419|T191|PT|31733|MEDCIN|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|ET|117|MEDLINEPLUS|Waldenstrom's Macroglobulinemia|9761/3
C0024419|T191|ET|D008258|MSH|Lymphoma, Lymphocytic, Plasmacytoid|9761/3
C0024419|T191|ET|D008258|MSH|Lymphoma, Lymphoplasmacytoid|9761/3
C0024419|T191|PM|D008258|MSH|Lymphomas, Lymphoplasmacytoid|9761/3
C0024419|T191|PM|D008258|MSH|Lymphoplasmacytoid Lymphoma|9761/3
C0024419|T191|PM|D008258|MSH|Lymphoplasmacytoid Lymphomas|9761/3
C0024419|T191|PM|D008258|MSH|Macroglobulinaemia, Waldenstrom's|9761/3
C0024419|T191|ET|D008258|MSH|Macroglobulinemia|9761/3
C0024419|T191|PM|D008258|MSH|Macroglobulinemia, Primary|9761/3
C0024419|T191|PM|D008258|MSH|Macroglobulinemia, Waldenstrom|9761/3
C0024419|T191|PM|D008258|MSH|Macroglobulinemia, Waldenstrom's|9761/3
C0024419|T191|ET|D008258|MSH|Primary Macroglobulinemia|9761/3
C0024419|T191|PM|D008258|MSH|Waldenstrom Macroglobulinaemia|9761/3
C0024419|T191|MH|D008258|MSH|Waldenstrom Macroglobulinemia|9761/3
C0024419|T191|ET|D008258|MSH|Waldenstrom's Macroglobulinaemia|9761/3
C0024419|T191|ET|D008258|MSH|Waldenstrom's Macroglobulinemia|9761/3
C0024419|T191|PM|D008258|MSH|Waldenstroms Macroglobulinaemia|9761/3
C0024419|T191|PM|D008258|MSH|Waldenstroms Macroglobulinemia|9761/3
C0334633|T191|PN|NOCODE|MTH|Malignant lymphoma - lymphoplasmacytic|9761/3
C0024419|T191|PN|NOCODE|MTH|Waldenstrom Macroglobulinemia|9761/3
C0334633|T191|ET|200.8|MTHICD9|Malignant lymphoplasmacytoid type lymphoma|9761/3
C0024419|T191|ET|273.3|MTHICD9|Primary macroglobulinemia|9761/3
C0024419|T191|ET|273.3|MTHICD9|Waldenstrom's macroglobulinemia|9761/3
C0334633|T191|OP|C3212|NCI|Immunocytoma, Lymphoplasmacytic Type|9761/3
C0334633|T191|SY|TCGA|NCI|Lymphoplasmacytic Lymphoma|9761/3
C0334633|T191|PT|C3212|NCI|Lymphoplasmacytic Lymphoma|9761/3
C0334633|T191|SY|C3212|NCI|Lymphoplasmacytoid Lymphoma|9761/3
C0024419|T191|SY|C80307|NCI|Waldenström Macroglobulinemia|9761/3
C0024419|T191|PT|C80307|NCI|Waldenstrom Macroglobulinemia|9761/3
C0024419|T191|SY|C80307|NCI|Waldenstrom's Macroglobulinemia|9761/3
C0334633|T191|SY|C3212|NCI_CDISC|Immunocytoma, Lymphoplasmacytic Type|9761/3
C0334633|T191|PT|C3212|NCI_CDISC|LYMPHOMA, LYMPHOPLASMACYTIC, MALIGNANT|9761/3
C0334633|T191|SY|C3212|NCI_CDISC|Lymphoma, Plasmacytic|9761/3
C0334633|T191|SY|C3212|NCI_CDISC|Lymphoplasmacytoid Lymphoma|9761/3
C0334633|T191|SY|10047803|NCI_CTEP-SDC|Lymphoplasmacytic lymphoma|9761/3
C0334633|T191|DN|C3212|NCI_CTRP|Lymphoplasmacytic Lymphoma|9761/3
C0024419|T191|DN|C80307|NCI_CTRP|Waldenstrom Macroglobulinemia|9761/3
C0334633|T191|PT|CDR0000409750|NCI_NCI-GLOSS|lymphoplasmacytic lymphoma|9761/3
C0024419|T191|PT|CDR0000044854|NCI_NCI-GLOSS|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|IS|CDR0000037790|PDQ|Immunocytoma, Lymphoplasmacytic Type|9761/3
C0024419|T191|SY|CDR0000037790|PDQ|lymphoplasmacytic lymphoma|9761/3
C0024419|T191|SY|CDR0000037790|PDQ|Lymphoplasmacytic Lymphoma/Waldenström Macroglobulinemia|9761/3
C0024419|T191|SY|CDR0000037790|PDQ|Lymphoplasmacytic Lymphoma/Waldenström's Macroglobulinemia|9761/3
C0024419|T191|SY|CDR0000037790|PDQ|lymphoplasmacytoid lymphoma|9761/3
C0024419|T191|SY|CDR0000037790|PDQ|macroglobulinemia|9761/3
C0024419|T191|SY|CDR0000037790|PDQ|macroglobulinemia, Waldenström's|9761/3
C0024419|T191|SY|CDR0000037790|PDQ|plasmacytoma, macroglobulinemia|9761/3
C0024419|T191|PT|CDR0000037790|PDQ|Waldenström macroglobulinemia|9761/3
C0024419|T191|SY|CDR0000037790|PDQ|Waldenström's macroglobulinemia|9761/3
C0024419|T191|PT|R0121913|QMR|WALDENSTROMS MACROGLOBULINEMIA|9761/3
C0334633|T191|SY|XaBBN|RCD|Immunocytoma|9761/3
C0024419|T191|PT|C333.|RCD|Macroglobulinaemia|9761/3
C0024419|T191|OP|C333z|RCD|Macroglobulinaemia NOS|9761/3
C0334633|T191|AB|XaBBN|RCD|Mal lymphoma, lymphoplasmacyt|9761/3
C0334633|T191|AB|XaBBN|RCD|Malignant lymph-lymphoplasmac|9761/3
C0334633|T191|PT|XaBBN|RCD|Malignant lymphoma - lymphoplasmacytic|9761/3
C0334633|T191|SY|XaBBN|RCD|Malignant lymphoma, lymphoplasmacytoid type|9761/3
C0334633|T191|SY|XaBBN|RCD|Plasmacytic lymphoma|9761/3
C0024419|T191|AB|C3330|RCD|Waldenstrom's macroglobulinaem|9761/3
C0024419|T191|PT|C3330|RCD|Waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|PT|C333.|RCDAE|Macroglobulinemia|9761/3
C0024419|T191|OP|C333z|RCDAE|Macroglobulinemia NOS|9761/3
C0024419|T191|PT|C3330|RCDAE|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|OP|XaBLz|RCDSA|Waldenstrom's macroglobulinemia|9761/3
C0334633|T191|AB|BBg7.|RCDSY|Malig.lymph,lymphoplasmacyt|9761/3
C0334633|T191|PT|BBg7.|RCDSY|Malignant lymphoma, lymphoplasmacytoid type|9761/3
C0024419|T191|OA|XaBLz|RCDSY|Waldenstrom's macroglobulin|9761/3
C0024419|T191|OP|XaBLz|RCDSY|Waldenstrom's macroglobulinaemia|9761/3
C0334633|T191|SY|307623001|SNOMEDCT_US|Immunocytoma|9761/3
C0334633|T191|SY|19340000|SNOMEDCT_US|Immunocytoma|9761/3
C0024419|T191|PTGB|190817009|SNOMEDCT_US|Macroglobulinaemia|9761/3
C0024419|T191|OAP|190821002|SNOMEDCT_US|Macroglobulinaemia NOS|9761/3
C0024419|T191|PT|190817009|SNOMEDCT_US|Macroglobulinemia|9761/3
C0024419|T191|OAP|190821002|SNOMEDCT_US|Macroglobulinemia NOS|9761/3
C0334633|T191|PT|307623001|SNOMEDCT_US|Malignant lymphoma - lymphoplasmacytic|9761/3
C0334633|T191|PT|19340000|SNOMEDCT_US|Malignant lymphoma, lymphoplasmacytic|9761/3
C0334633|T191|SY|19340000|SNOMEDCT_US|Malignant lymphoma, lymphoplasmacytoid|9761/3
C0334633|T191|SY|307623001|SNOMEDCT_US|Malignant lymphoma, lymphoplasmacytoid type|9761/3
C0334633|T191|SY|19340000|SNOMEDCT_US|Malignant lymphoma, plasmacytoid|9761/3
C0334633|T191|SY|307623001|SNOMEDCT_US|Plasmacytic lymphoma|9761/3
C0334633|T191|SY|19340000|SNOMEDCT_US|Plasmacytic lymphoma|9761/3
C0024419|T191|SYGB|35562000|SNOMEDCT_US|Primary macroglobulinaemia|9761/3
C0024419|T191|SY|35562000|SNOMEDCT_US|Primary macroglobulinemia|9761/3
C0024419|T191|PTGB|190818004|SNOMEDCT_US|Waldenström macroglobulinaemia|9761/3
C0024419|T191|SYGB|35562000|SNOMEDCT_US|Waldenstrom macroglobulinaemia|9761/3
C0024419|T191|SY|35562000|SNOMEDCT_US|Waldenstrom macroglobulinemia|9761/3
C0024419|T191|PT|190818004|SNOMEDCT_US|Waldenström macroglobulinemia|9761/3
C0024419|T191|OAS|154750002|SNOMEDCT_US|Waldenstrom's macroglob'naemia|9761/3
C0024419|T191|OAS|267503004|SNOMEDCT_US|Waldenstrom's macroglob'naemia|9761/3
C0024419|T191|PTGB|35562000|SNOMEDCT_US|Waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|OAS|267503004|SNOMEDCT_US|Waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|SYGB|190818004|SNOMEDCT_US|Waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|OAS|154750002|SNOMEDCT_US|Waldenstrom's macroglobulinaemia|9761/3
C0024419|T191|OAS|154750002|SNOMEDCT_US|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|PT|35562000|SNOMEDCT_US|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|OAS|267503004|SNOMEDCT_US|Waldenstrom's macroglobulinemia|9761/3
C0024419|T191|SY|190818004|SNOMEDCT_US|Waldenstrom's macroglobulinemia|9761/3
C0018852|T191|PT|0000005912|CHV|heavy chain disease|9762/3
C0018852|T191|PT|0449-3246|CSP|heavy chain disease|9762/3
C0018852|T191|SY|NOCODE|DXP|BALLARD DISEASE|9762/3
C0018852|T191|DI|U000782|DXP|HEAVY CHAIN DISEASE|9762/3
C0018852|T191|SY|NOCODE|DXP|SELIGMANN DISEASE|9762/3
C0018852|T191|AB|C88.2|ICD10CM|Heavy chain disease|9762/3
C0018852|T191|PT|C88.2|ICD10CM|Heavy chain disease|9762/3
C0018852|T191|LLT|10019350|MDR|Heavy chain disease|9762/3
C0018852|T191|PT|10019350|MDR|Heavy chain disease|9762/3
C0018852|T191|PT|33893|MEDCIN|heavy chain disease|9762/3
C0018852|T191|DEV|D006362|MSH|HEAVY CHAIN DIS|9762/3
C0018852|T191|MH|D006362|MSH|Heavy Chain Disease|9762/3
C0018852|T191|PM|D006362|MSH|Heavy Chain Diseases|9762/3
C0018852|T191|PN|NOCODE|MTH|Heavy Chain Disease|9762/3
C0018852|T191|AB|C3082|NCI|HCD|9762/3
C0018852|T191|PT|C3082|NCI|Heavy Chain Disease|9762/3
C0018852|T191|SY|TCGA|NCI|Heavy Chain Disease|9762/3
C0018852|T191|PT|Xa0SM|RCD|Heavy chain disease|9762/3
C0018852|T191|PT|68979007|SNOMEDCT_US|Heavy chain disease|9762/3
C0018852|T191|PT|6381009|SNOMEDCT_US|Heavy chain disease|9762/3
C0018852|T191|IS|68979007|SNOMEDCT_US|Heavy chain disease, NOS|9762/3
C0021071|T191|SY|0000006611|CHV|alpha-chain disease|9764/3
C0021071|T191|SY|0000006611|CHV|chain alpha disease|9764/3
C0021071|T191|PT|0000006611|CHV|ipsid|9764/3
C0021071|T191|SY|NOCODE|DXP|ALPHA CHAIN DISEASE|9764/3
C0021071|T191|SY|NOCODE|DXP|ALPHA HCD|9764/3
C0021071|T191|SY|NOCODE|DXP|ALPHA HEAVY CHAIN DISEASE|9764/3
C0021071|T191|SY|NOCODE|DXP|ALPHA-HEAVY CHAIN DISEASE|9764/3
C0021071|T191|SY|NOCODE|DXP|IGA HEAVY CHAIN DISEASE|9764/3
C0021071|T191|SY|NOCODE|DXP|IMMUNOPROLIFERATIVE SMALL INTESTINE DISEASE|9764/3
C0021071|T191|SY|NOCODE|DXP|IPSID|9764/3
C0021071|T191|ET|HP:0020194|HPO|Alpha heavy chain disease|9764/3
C0021071|T191|PT|C88.1|ICD10|Alpha heavy chain disease|9764/3
C0021071|T191|PT|C88.3|ICD10|Immunoproliferative small intestinal disease|9764/3
C0021071|T191|ET|C88.3|ICD10CM|Alpha heavy chain disease|9764/3
C0021071|T191|PT|C88.3|ICD10CM|Immunoproliferative small intestinal disease|9764/3
C0021071|T191|AB|C88.3|ICD10CM|Immunoproliferative small intestinal disease|9764/3
C0021071|T191|ET|C88.3|ICD10CM|Mediterranean lymphoma|9764/3
C0021071|T191|PT|MTHU005087|ICPC2ICD10ENG|alpha heavy chain; disease|9764/3
C0021071|T191|PT|MTHU004932|ICPC2ICD10ENG|alpha; alpha heavy chain disease|9764/3
C0021071|T191|PT|MTHU023293|ICPC2ICD10ENG|disease; alpha heavy chain|9764/3
C0021071|T191|PT|MTHU033693|ICPC2ICD10ENG|heavy chain alpha|9764/3
C0021071|T191|PT|MTHU090250|ICPC2ICD10ENG|immunoproliferative; disease, small intestine|9764/3
C0021071|T191|PT|MTHU046826|ICPC2ICD10ENG|lymphoma; mediterranean|9764/3
C0021071|T191|PT|MTHU049176|ICPC2ICD10ENG|mediterranean; lymphoma|9764/3
C0021071|T191|PT|351185|MEDCIN|Alpha heavy chain disease|9764/3
C0021071|T191|PT|351186|MEDCIN|Alpha heavy chain disease, enteric form|9764/3
C0021071|T191|SY|351185|MEDCIN|heavy chain disease alpha|9764/3
C0021071|T191|SY|351186|MEDCIN|heavy chain disease alpha, enteric form|9764/3
C0021071|T191|SY|31572|MEDCIN|immunoproliferative intestinal disease|9764/3
C0021071|T191|PT|31572|MEDCIN|immunoproliferative small intestinal disease|9764/3
C0021071|T191|DEV|D007161|MSH|ALPHA CHAIN DIS|9764/3
C0021071|T191|PM|D007161|MSH|alpha Chain Disease|9764/3
C0021071|T191|ET|D007161|MSH|alpha-Chain Disease|9764/3
C0021071|T191|PM|D007161|MSH|alpha-Chain Diseases|9764/3
C0021071|T191|PM|D007161|MSH|Disease, alpha-Chain|9764/3
C0021071|T191|PM|D007161|MSH|Diseases, alpha-Chain|9764/3
C0021071|T191|DEV|D007161|MSH|HEAVY CHAIN DIS IGA TYPE|9764/3
C0021071|T191|ET|D007161|MSH|Heavy Chain Disease, IgA Type|9764/3
C0021071|T191|DEV|D007161|MSH|IMMUNOPROLIFERATIVE SMALL INTESTINAL DIS|9764/3
C0021071|T191|MH|D007161|MSH|Immunoproliferative Small Intestinal Disease|9764/3
C0021071|T191|ET|D007161|MSH|IPSID|9764/3
C0021071|T191|ET|D007161|MSH|Lymphoma, Mediterranean|9764/3
C0021071|T191|PM|D007161|MSH|Mediterranean Lymphoma|9764/3
C0021071|T191|PT|C3132|NCI|Alpha Heavy Chain Disease|9764/3
C0021071|T191|SY|C3132|NCI|Immunoproliferative Small Intestinal Disease|9764/3
C0021071|T191|AB|C3132|NCI|IPSID|9764/3
C0021071|T191|SY|C3132|NCI|Mediterranean Abdominal Lymphoma|9764/3
C0021071|T191|SY|C3132|NCI|Mediterranean Lymphoma|9764/3
C0021071|T191|OP|C3331|RCD|Alpha heavy chain disease|9764/3
C0021071|T191|OP|BBm6.|RCDSY|Alpha heavy chain disease|9764/3
C0021071|T191|OP|BBmG.|RCDSY|Immunoproliferative small intestinal disease|9764/3
C0021071|T191|OA|BBmG.|RCDSY|Imunoprolif smal intest dis|9764/3
C0021071|T191|SY|109982002|SNOMEDCT_US|Alpha heavy chain disease|9764/3
C0021071|T191|OAP|190819007|SNOMEDCT_US|Alpha heavy chain disease|9764/3
C0021071|T191|SY|6381009|SNOMEDCT_US|Alpha heavy chain disease|9764/3
C0021071|T191|OAP|123312002|SNOMEDCT_US|Alpha heavy chain disease|9764/3
C0021071|T191|OF|123312002|SNOMEDCT_US|Alpha heavy chain disease -RETIRED-|9764/3
C0021071|T191|IS|123312002|SNOMEDCT_US|Alpha heavy chain disease -RETIRED-|9764/3
C0021071|T191|PT|123313007|SNOMEDCT_US|Alpha heavy chain disease, enteric form|9764/3
C0021071|T191|SY|27461004|SNOMEDCT_US|Alpha heavy chain disease, enteric form|9764/3
C0021071|T191|IS|123312002|SNOMEDCT_US|Alpha heavy chain disease, NOS|9764/3
C0021071|T191|SY|6381009|SNOMEDCT_US|IgA heavy chain disease|9764/3
C0021071|T191|IS|6381009|SNOMEDCT_US|IgA heavy chain disease, NOS|9764/3
C0021071|T191|IS|123312002|SNOMEDCT_US|IgA heavy chain disease, NOS|9764/3
C0021071|T191|PT|27461004|SNOMEDCT_US|Immunoproliferative small intestinal disease|9764/3
C0021071|T191|SY|109985000|SNOMEDCT_US|Immunoproliferative small intestinal disease|9764/3
C0021071|T191|IS|123313007|SNOMEDCT_US|Immunoproliferative small intestinal disease|9764/3
C0021071|T191|SY|27461004|SNOMEDCT_US|Mediterranean lymphoma|9764/3
C0021071|T191|IS|123313007|SNOMEDCT_US|Mediterranean lymphoma|9764/3
C0026470|T191|PT|0011617|CCPSS|GAMMOPATHY MONOCLONAL BENIGN|9765/1
C0026470|T191|PT|0014467|CCPSS|GAMMOPATHY MONOCLONAL UNCERTAIN SIGNIFICANCE|9765/1
C0026470|T191|SY|0000008234|CHV|benign monoclonal gammapathy|9765/1
C0026470|T191|PT|0000008234|CHV|benign monoclonal gammopathy|9765/1
C0026470|T191|SY|0000027191|CHV|gammopathy monoclonal|9765/1
C0026470|T191|SY|0000027191|CHV|mgus|9765/1
C0026470|T191|PT|0000027191|CHV|monoclonal gammopathy|9765/1
C0026470|T191|PT|U000069|COSTAR|BENIGN MONOCLONAL HYPERGAMMAGLOBUMINEMIA|9765/1
C0026470|T191|DI|U000204|DXP|BENIGN MONOCLONAL GAMMOPATHY|9765/1
C0026470|T191|PT|MTHU030242|ICPC2ICD10ENG|gammopathy; monoclonal, of undetermined significance|9765/1
C0026470|T191|PT|MTHU050302|ICPC2ICD10ENG|monoclonal; gammopathy, of undetermined significance|9765/1
C0026470|T191|LLT|10004293|MDR|Benign monoclonal hypergammaglobulinaemia|9765/1
C0026470|T191|LLT|10060563|MDR|Benign monoclonal hypergammaglobulinemia|9765/1
C0026470|T191|LLT|10020631|MDR|Hypergammaglobulinaemia benign monoclonal|9765/1
C0026470|T191|PT|10020631|MDR|Hypergammaglobulinaemia benign monoclonal|9765/1
C0026470|T191|LLT|10054409|MDR|Hypergammaglobulinemia benign monoclonal|9765/1
C0026470|T191|MTH_PT|10020631|MDR|Hypergammaglobulinemia benign monoclonal|9765/1
C0026470|T191|LLT|10027522|MDR|MGUS|9765/1
C0026470|T191|OL|10027523|MDR|MGUS undetermined|9765/1
C0026470|T191|LLT|10027863|MDR|Monoclonal gammopathy of unknown significance|9765/1
C0026470|T191|PT|31812|MEDCIN|benign monoclonal hypergammaglobulinemia|9765/1
C0026470|T191|PT|276394|MEDCIN|monoclonal gammopathy of undetermined significance|9765/1
C0026470|T191|PM|D008998|MSH|Benign Monoclonal Gammapathies|9765/1
C0026470|T191|PM|D008998|MSH|Benign Monoclonal Gammapathy|9765/1
C0026470|T191|ET|D008998|MSH|Benign Monoclonal Gammopathies|9765/1
C0026470|T191|PM|D008998|MSH|Benign Monoclonal Gammopathy|9765/1
C0026470|T191|ET|D008998|MSH|Monoclonal Gammapathies, Benign|9765/1
C0026470|T191|ET|D008998|MSH|Monoclonal Gammapathy of Undetermined Significance|9765/1
C0026470|T191|PM|D008998|MSH|Monoclonal Gammapathy, Benign|9765/1
C0026470|T191|ET|D008998|MSH|Monoclonal Gammopathies, Benign|9765/1
C0026470|T191|MH|D008998|MSH|Monoclonal Gammopathy of Undetermined Significance|9765/1
C0026470|T191|PM|D008998|MSH|Monoclonal Gammopathy, Benign|9765/1
C0026470|T191|PN|NOCODE|MTH|Monoclonal Gammopathy of Undetermined Significance|9765/1
C0026470|T191|ET|273.1|MTHICD9|Benign monoclonal gammopathy|9765/1
C0026470|T191|ET|273.1|MTHICD9|Benign monoclonal hypergammaglobulinemia|9765/1
C0026470|T191|ET|273.1|MTHICD9|BMH|9765/1
C0026470|T191|AB|C3996|NCI|MGUS|9765/1
C0026470|T191|PT|C3996|NCI|Monoclonal Gammopathy of Undetermined Significance|9765/1
C0026470|T191|SY|TCGA|NCI|Monoclonal Gammopathy of Undetermined Significance|9765/1
C0026470|T191|SY|10020631|NCI_CTEP-SDC|MGUS|9765/1
C0026470|T191|DN|C3996|NCI_CTRP|Monoclonal Gammopathy of Undetermined Significance|9765/1
C0026470|T191|PT|CDR0000411380|NCI_NCI-GLOSS|MGUS|9765/1
C0026470|T191|PT|CDR0000411379|NCI_NCI-GLOSS|monoclonal gammopathy of undetermined significance|9765/1
C0026470|T191|SY|CDR0000040134|PDQ|Benign Monoclonal Gammopathy|9765/1
C0026470|T191|AB|CDR0000040134|PDQ|MGUS|9765/1
C0026470|T191|PT|CDR0000040134|PDQ|monoclonal gammopathy of undetermined significance|9765/1
C0026470|T191|SY|CDR0000040134|PDQ|Monoclonal Gammopathy of Unknown Significance|9765/1
C0026470|T191|SY|CDR0000040134|PDQ|plasma cell neoplasm, monoclonal gammopathy of unknown significance|9765/1
C0026470|T191|SY|Xa0SJ|RCD|MGUS - Monoclonal gammopathy of uncertain significance|9765/1
C0026470|T191|AB|Xa0SJ|RCD|MGUS-Mono gammop uncert signif|9765/1
C0026470|T191|AB|Xa0SJ|RCD|Mono gammop uncert significanc|9765/1
C0026470|T191|PT|Xa0SJ|RCD|Monoclonal gammopathy of uncertain significance|9765/1
C0026470|T191|SY|58648008|SNOMEDCT_US|Asymptomatic monoclonal gammopathy|9765/1
C0026470|T191|PT|58648008|SNOMEDCT_US|Benign monoclonal gammopathy|9765/1
C0026470|T191|SY|35601003|SNOMEDCT_US|MGUS|9765/1
C0026470|T191|SY|277577000|SNOMEDCT_US|MGUS - Monoclonal gammopathy of uncertain significance|9765/1
C0026470|T191|PT|277577000|SNOMEDCT_US|Monoclonal gammopathy of uncertain significance|9765/1
C0026470|T191|PT|35601003|SNOMEDCT_US|Monoclonal gammopathy of undetermined significance|9765/1
C0026470|T191|SY|277577000|SNOMEDCT_US|Monoclonal gammopathy of undetermined significance|9765/1
C0024307|T191|PT|0025295|CCPSS|LYMPHOMATOID GRANULOMATOSIS|9766/1
C0024307|T191|PT|0000007622|CHV|lymphomatoid granulomatosis|9766/1
C0024307|T191|DI|U001122|DXP|LYMPHOMATOID GRANULOMATOSIS|9766/1
C0024307|T191|ET|C83.8|ICD10CM|Lymphoid granulomatosis|9766/1
C0024307|T191|PT|MTHU006354|ICPC2ICD10ENG|angiocentric immunoproliferative; lesion|9766/1
C0024307|T191|PT|MTHU032713|ICPC2ICD10ENG|granulomatosis; lymphoid|9766/1
C0024307|T191|PT|MTHU043372|ICPC2ICD10ENG|lesion; angiocentric immunoproliferative|9766/1
C0024307|T191|PT|MTHU046726|ICPC2ICD10ENG|lymphoid; granulomatosis|9766/1
C0024307|T191|LLT|10025325|MDR|Lymphomatoid granulomatosis|9766/1
C0024307|T191|PT|31832|MEDCIN|lymphomatoid granulomatosis|9766/1
C0024307|T191|PM|D008230|MSH|Granulomatoses, Lymphomatoid|9766/1
C0024307|T191|ET|D008230|MSH|Granulomatosis, Lymphomatoid|9766/1
C0024307|T191|PM|D008230|MSH|Lymphomatoid Granulomatoses|9766/1
C0024307|T191|MH|D008230|MSH|Lymphomatoid Granulomatosis|9766/1
C0024307|T191|PN|NOCODE|MTH|Lymphomatoid Granulomatosis|9766/1
C0024307|T191|AB|C40970|NCI|AIL|9766/1
C0024307|T191|PT|C40970|NCI|Angiocentric Immunoproliferative Lesion|9766/1
C0024307|T191|AB|C7930|NCI|LYG|9766/1
C0024307|T191|PT|C7930|NCI|Lymphomatoid Granulomatosis|9766/1
C0024307|T191|SY|TCGA|NCI|Lymphomatoid Granulomatosis|9766/1
C0024307|T191|PT|10025325|NCI_CTEP-SDC|Lymphomatoid granulomatosis|9766/1
C0024307|T191|PT|CDR0000045766|NCI_NCI-GLOSS|lymphomatoid granulomatosis|9766/1
C0024307|T191|IS|CDR0000039048|PDQ|angiocentric immunoproliferative lesions|9766/1
C0024307|T191|PT|R0121670|QMR|LYMPHOMATOID GRANULOMATOSIS|9766/1
C0024307|T191|AB|X705o|RCD|LG - Lymphomatoid granulomatos|9766/1
C0024307|T191|SY|X705o|RCD|LG - Lymphomatoid granulomatosis|9766/1
C0024307|T191|PT|X705o|RCD|Lymphomatoid granulomatosis|9766/1
C0024307|T191|OA|BBmF.|RCDSY|Angiocent immunoprolif lesn|9766/1
C0024307|T191|OP|BBmF.|RCDSY|Angiocentric immunoproliferative lesion|9766/1
C0024307|T191|PT|41556003|SNOMEDCT_US|Angiocentric immunoproliferative lesion|9766/1
C0024307|T191|SY|239940004|SNOMEDCT_US|LG - Lymphomatoid granulomatosis|9766/1
C0024307|T191|IS|41556003|SNOMEDCT_US|Lymphmatoid granulomatosis|9766/1
C0024307|T191|IS|41556003|SNOMEDCT_US|Lymphoid granulomatosis|9766/1
C0024307|T191|PT|789177000|SNOMEDCT_US|Lymphomatoid granulomatosis|9766/1
C0024307|T191|OAP|60337005|SNOMEDCT_US|Lymphomatoid granulomatosis|9766/1
C0024307|T191|PT|239940004|SNOMEDCT_US|Lymphomatoid granulomatosis|9766/1
C5230382|T191|PT|789178005|SNOMEDCT_US|Lymphomatoid granulomatosis grade 1|9766/1
C5230383|T191|PT|789179002|SNOMEDCT_US|Lymphomatoid granulomatosis grade 2|9766/1
C0020981|T191|SY|0000006589|CHV|aild|9767/1
C0020981|T191|SY|0000006589|CHV|angioblastic lymphadenopathy|9767/1
C0020981|T191|PT|0000006589|CHV|angioimmunoblastic lymphadenopathy|9767/1
C0020981|T191|SY|0000006589|CHV|angioimmunoblastic lymphoma|9767/1
C0020981|T191|SY|0000006589|CHV|immunoblastic lymphadenopathy|9767/1
C0020981|T191|DI|U001112|DXP|LYMPHADENOPATHY, ANGIOIMMUNOBLASTIC, WITH DYSPROTEINEMIA|9767/1
C0020981|T191|SY|NOCODE|DXP|LYMPHADENOPATHY, IMMUNOBLASTIC|9767/1
C0020981|T191|AB|C86.5|ICD10CM|Angioimmunoblastic T-cell lymphoma|9767/1
C0020981|T191|PT|C86.5|ICD10CM|Angioimmunoblastic T-cell lymphoma|9767/1
C0020981|T191|PT|MTHU006365|ICPC2ICD10ENG|angioimmunoblastic; lymphadenopathy|9767/1
C0020981|T191|PT|MTHU006366|ICPC2ICD10ENG|angioimmunoblastic; lymphoma|9767/1
C0020981|T191|PT|MTHU046565|ICPC2ICD10ENG|lymphadenopathy; angioimmunoblastic|9767/1
C0020981|T191|PT|MTHU046737|ICPC2ICD10ENG|lymphoma; angioimmunoblastic|9767/1
C0020981|T191|LLT|10080248|MDR|Angioimmunoblastic lymphadenopathy|9767/1
C0020981|T191|LLT|10079289|MDR|Angioimmunoblastic lymphadenopathy with dysproteinaemia|9767/1
C0020981|T191|LLT|10079282|MDR|Angioimmunoblastic lymphadenopathy with dysproteinemia|9767/1
C0020981|T191|LLT|10002449|MDR|Angioimmunoblastic T-cell lymphoma|9767/1
C0020981|T191|PT|10002449|MDR|Angioimmunoblastic T-cell lymphoma|9767/1
C0020981|T191|LLT|10002451|MDR|Angioimmunoblastic T-cell lymphoma NOS|9767/1
C0020981|T191|HT|10002450|MDR|Angioimmunoblastic T-cell lymphomas|9767/1
C0020981|T191|SY|31466|MEDCIN|AILD|9767/1
C0020981|T191|PT|31466|MEDCIN|angioimmunoblastic T-cell lymphoma|9767/1
C0020981|T191|SY|33782|MEDCIN|immunoblastic lymphadenopathy|9767/1
C0020981|T191|PT|33782|MEDCIN|malignant immunoblastic lymphadenopathy|9767/1
C0020981|T191|PM|D007119|MSH|Angioimmunoblastic Lymphadenopathies|9767/1
C0020981|T191|ET|D007119|MSH|Angioimmunoblastic Lymphadenopathy|9767/1
C0020981|T191|PM|D007119|MSH|Immunoblastic Lymphadenopathies|9767/1
C0020981|T191|MH|D007119|MSH|Immunoblastic Lymphadenopathy|9767/1
C0020981|T191|PM|D007119|MSH|Lymphadenopathies, Angioimmunoblastic|9767/1
C0020981|T191|PM|D007119|MSH|Lymphadenopathies, Immunoblastic|9767/1
C0020981|T191|PM|D007119|MSH|Lymphadenopathy, Angioimmunoblastic|9767/1
C0020981|T191|ET|D007119|MSH|Lymphadenopathy, Immunoblastic|9767/1
C0020981|T191|PN|NOCODE|MTH|Angioimmunoblastic Lymphadenopathy|9767/1
C0020981|T191|AB|C7528|NCI|AILD|9767/1
C0020981|T191|AB|C7528|NCI|AILT|9767/1
C0020981|T191|OP|C7528|NCI|Angioimmunoblastic Lymphadenopathy|9767/1
C0020981|T191|SY|C7528|NCI|Angioimmunoblastic Lymphadenopathy Type T-Cell Lymphoma|9767/1
C0020981|T191|OP|C7528|NCI|Angioimmunoblastic Lymphadenopathy with Dysproteinemia|9767/1
C0020981|T191|PT|C7528|NCI|Angioimmunoblastic T-Cell Lymphoma|9767/1
C0020981|T191|SY|TCGA|NCI|Angioimmunoblastic T-Cell Lymphoma|9767/1
C0020981|T191|PT|C7528|NCI_CPTAC|Angioimmunoblastic T-Cell Lymphoma|9767/1
C0020981|T191|DN|C7528|NCI_CTRP|Angioimmunoblastic T-Cell Lymphoma|9767/1
C0020981|T191|PT|CDR0000346464|NCI_NCI-GLOSS|angioimmunoblastic T-cell lymphoma|9767/1
C0020981|T191|AB|CDR0000042765|PDQ|AILD|9767/1
C0020981|T191|AB|CDR0000042765|PDQ|AILT|9767/1
C0020981|T191|IS|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy|9767/1
C0020981|T191|SY|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy|9767/1
C0020981|T191|SY|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy type T-cell lymphoma|9767/1
C0020981|T191|SY|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy with dysproteinemia|9767/1
C0020981|T191|IS|CDR0000042765|PDQ|angioimmunoblastic lymphadenopathy with dysproteinemia|9767/1
C0020981|T191|PT|CDR0000042765|PDQ|angioimmunoblastic T-cell lymphoma|9767/1
C0020981|T191|PT|Q0300328|QMR|ANGIOIMMUNOBLASTIC LYMPHADENOPATHY|9767/1
C0020981|T191|AB|Xa0Tk|RCD|Angioim lymphadenopy+dysprot|9767/1
C0020981|T191|PT|Xa0Tk|RCD|Angioimmunoblastic lymphadenopathy with dysproteinaemia|9767/1
C0020981|T191|SY|Xa0Tk|RCD|Angioimmunoblastic lymphoma|9767/1
C0020981|T191|PT|Xa0Tk|RCDAE|Angioimmunoblastic lymphadenopathy with dysproteinemia|9767/1
C0020981|T191|OA|BBm8.|RCDSY|Angioimmunoblas lymphadenop|9767/1
C0020981|T191|OP|BBm8.|RCDSY|Angioimmunoblastic lymphadenopathy|9767/1
C0020981|T191|OAS|127216000|SNOMEDCT_US|AILD|9767/1
C0020981|T191|PT|52097008|SNOMEDCT_US|Angioimmunoblastic lymphadenopathy|9767/1
C0020981|T191|OAP|127216000|SNOMEDCT_US|Angioimmunoblastic lymphadenopathy with dysproteinaemia|9767/1
C0020981|T191|OAP|127216000|SNOMEDCT_US|Angioimmunoblastic lymphadenopathy with dysproteinemia|9767/1
C0020981|T191|SY|835009|SNOMEDCT_US|Angioimmunoblastic lymphoma|9767/1
C0020981|T191|PT|413537009|SNOMEDCT_US|Angioimmunoblastic T-cell lymphoma|9767/1
C0020981|T191|PT|835009|SNOMEDCT_US|Angioimmunoblastic T-cell lymphoma|9767/1
C1955861|T191|PT|MTHU046872|ICPC2ICD10ENG|lymphoproliferative; disease, T-gamma|9768/1
C1955861|T191|LLT|10065862|MDR|T-cell large granular lymphocytic leukemia|9768/1
C1955861|T191|SY|392217|MEDCIN|leukemia lymphocytic chronic T-cell large granular|9768/1
C1955861|T191|PT|392217|MEDCIN|T-cell large granular lymphocytic leukemia|9768/1
C1955861|T191|PM|D054066|MSH|Granular Lymphocytoses, Large|9768/1
C1955861|T191|PM|D054066|MSH|Granular Lymphocytosis, Large|9768/1
C1955861|T191|PM|D054066|MSH|Large Granular Lymphocytoses|9768/1
C1955861|T191|ET|D054066|MSH|Large Granular Lymphocytosis|9768/1
C1955861|T191|PM|D054066|MSH|Leukemia, T Cell Large Granular Lymphocytic|9768/1
C1955861|T191|PM|D054066|MSH|Leukemia, T LGL|9768/1
C1955861|T191|PEP|D054066|MSH|Leukemia, T-Cell Large Granular Lymphocytic|9768/1
C1955861|T191|ET|D054066|MSH|Leukemia, T-LGL|9768/1
C1955861|T191|PM|D054066|MSH|Leukemias, T-LGL|9768/1
C1955861|T191|PM|D054066|MSH|Lymphocytoses, Large Granular|9768/1
C1955861|T191|PM|D054066|MSH|Lymphocytosis, Large Granular|9768/1
C1955861|T191|PM|D054066|MSH|T Cell Large Granular Lymphocyte Leukemia|9768/1
C1955861|T191|PM|D054066|MSH|T Cell Large Granular Lymphocytic Leukemia|9768/1
C1955861|T191|PM|D054066|MSH|T LGL Leukemia|9768/1
C1955861|T191|ET|D054066|MSH|T-Cell Large Granular Lymphocyte Leukemia|9768/1
C1955861|T191|ET|D054066|MSH|T-Cell Large Granular Lymphocytic Leukemia|9768/1
C1955861|T191|ET|D054066|MSH|T-LGL Leukemia|9768/1
C1955861|T191|PM|D054066|MSH|T-LGL Leukemias|9768/1
C1955861|T191|PN|NOCODE|MTH|T-Cell Large Granular Lymphocyte Leukemia|9768/1
C1955861|T191|SY|C4664|NCI|Large Cell Granular Lymphogenous Leukemia|9768/1
C1955861|T191|SY|C4664|NCI|Large Cell Granular Lymphoid Leukemia|9768/1
C1955861|T191|SY|C4664|NCI|Large Granular Lymphocytic Leukemia|9768/1
C1955861|T191|SY|C4664|NCI|Large Granular Lymphocytosis|9768/1
C1955861|T191|AB|C4664|NCI|LGLL|9768/1
C1955861|T191|SY|C4664|NCI|T Gamma Lymphoproliferative Disorder|9768/1
C1955861|T191|SY|TCGA|NCI|T-Cell Large Granular Lymphocyte Leukemia|9768/1
C1955861|T191|PT|C4664|NCI|T-Cell Large Granular Lymphocyte Leukemia|9768/1
C1955861|T191|SY|C4664|NCI|T-Cell Large Granular Lymphocytic Leukemia|9768/1
C1955861|T191|SY|C4664|NCI|T-Gamma Lymphoproliferative Disorder|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|Large Cell Granular Lymphogenous Leukemia|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|Large Cell Granular Lymphoid Leukemia|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|Large Granular Lymphocytic Leukemia|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|Large Granular Lymphocytosis|9768/1
C1955861|T191|PT|C4664|NCI_CDISC|LEUKEMIA, LARGE GRANULAR LYMPHOCYTIC, MALIGNANT|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|LGLL|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|T Gamma Lymphoproliferative Disorder|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|T-Cell Large Granular Lymphocytic Leukemia|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|T-Gamma Lymphoproliferative Disorder|9768/1
C1955861|T191|SY|C4664|NCI_CDISC|Tgamma Large Granular Lymphocyte Leukemia|9768/1
C1955861|T191|SY|10065862|NCI_CTEP-SDC|T-cell large gran. lymph. leuk.|9768/1
C1955861|T191|PT|10065862|NCI_CTEP-SDC|T-cell large granular lymphocytic leukemia|9768/1
C1955861|T191|DN|C4664|NCI_CTRP|T-Cell Large Granular Lymphocyte Leukemia|9768/1
C1955861|T191|PT|CDR0000633892|NCI_NCI-GLOSS|T-cell large granular lymphocyte leukemia|9768/1
C1955861|T191|PT|CDR0000633893|NCI_NCI-GLOSS|T-LGL leukemia|9768/1
C1955861|T191|PT|CDR0000039823|PDQ|T-cell large granular lymphocyte leukemia|9768/1
C1955861|T191|OP|CDR0000040442|PDQ|T-gamma lymphoproliferative disorder|9768/1
C1955861|T191|SY|CDR0000039823|PDQ|T-gamma lymphoproliferative disorder|9768/1
C1955861|T191|OA|BBmC.|RCDSY|T-gam lymphoprolif disease|9768/1
C1955861|T191|OP|BBmC.|RCDSY|T-gamma lymphoproliferative disease|9768/1
C1955861|T191|PTGB|699818003|SNOMEDCT_US|T-cell large granular lymphocytic leukaemia|9768/1
C1955861|T191|PTGB|128819001|SNOMEDCT_US|T-cell large granular lymphocytic leukaemia|9768/1
C1955861|T191|PT|699818003|SNOMEDCT_US|T-cell large granular lymphocytic leukemia|9768/1
C1955861|T191|PT|128819001|SNOMEDCT_US|T-cell large granular lymphocytic leukemia|9768/1
C1955861|T191|SY|128819001|SNOMEDCT_US|T-cell large granular lymphocytosis|9768/1
C1955861|T191|PT|55081009|SNOMEDCT_US|T-gamma lymphoproliferative disease|9768/1
C2939462|T191|PN|NOCODE|MTH|Immunoglobulin deposition disease|9769/1
C2939462|T191|SY|C7151|NCI|Immunoglobulin Deposition Disease|9769/1
C2939462|T191|PT|C7151|NCI|Monoclonal Immunoglobulin Deposition Disease|9769/1
C2939462|T191|PT|C7151|NCI_CPTAC|Monoclonal Immunoglobulin Deposition Disease|9769/1
C2939462|T191|DN|C7151|NCI_CTRP|Monoclonal Immunoglobulin Deposition Disease|9769/1
C2939462|T191|SY|CDR0000618304|PDQ|Immunoglobulin Deposition Disease|9769/1
C2939462|T191|PT|CDR0000618304|PDQ|monoclonal immunoglobulin deposition disease|9769/1
C2939462|T191|PT|128817004|SNOMEDCT_US|Immunoglobulin deposition disease|9769/1
C2939462|T191|SY|128817004|SNOMEDCT_US|Primary amyloidosis|9769/1
C2939462|T191|SY|128817004|SNOMEDCT_US|Systemic light chain disease|9769/1
C0023418|T191|ET|0000004617|AOD|leukemia|9800/3
C0023418|T191|PT|BI00316|BI|leukemia|9800/3
C0023418|T191|PT|0051957|CCPSS|LEUKEMIA|9800/3
C0023418|T191|MD|2.10.3|CCS|Leukemias|9800/3
C0023418|T191|SD|39|CCS|Leukemias|9800/3
C0023418|T191|PT|0000049549|CHV|all types of leukemia|9800/3
C0023418|T191|SY|0000007330|CHV|leukaemia|9800/3
C0023418|T191|SY|0000007330|CHV|leukaemias|9800/3
C0023418|T191|PT|0000007330|CHV|leukemia|9800/3
C0023418|T191|SY|0000049549|CHV|leukemia type|9800/3
C0023418|T191|SY|0000049549|CHV|leukemia types|9800/3
C0023418|T191|SY|0000007330|CHV|leukemias|9800/3
C0023418|T191|SY|0000049549|CHV|leukemias types|9800/3
C0023418|T191|SY|0000049549|CHV|type leukemia|9800/3
C0023418|T191|SY|0000049549|CHV|types leukemia|9800/3
C0023418|T191|PT|U000412|COSTAR|LEUKEMIA|9800/3
C0023418|T191|PT|2004-1566|CSP|leukemia|9800/3
C0023418|T191|GT|LEUKEMIA|CST|LEUKAEMIA|9800/3
C0023418|T191|PT|LEUKEMIA|CST|LEUKEMIA|9800/3
C0023418|T191|FI|U002348|DXP|LEUKEMIA|9800/3
C0023418|T191|PT|HP:0001909|HPO|Leukemia|9800/3
C0023418|T191|HT|C95|ICD10|Leukaemia of unspecified cell type|9800/3
C0023418|T191|PT|C95.9|ICD10|Leukaemia, unspecified|9800/3
C0023418|T191|HT|C95|ICD10AE|Leukemia of unspecified cell type|9800/3
C0023418|T191|PT|C95.9|ICD10AE|Leukemia, unspecified|9800/3
C0023418|T191|ET|C95.90|ICD10CM|Leukemia NOS|9800/3
C0023418|T191|AB|C95|ICD10CM|Leukemia of unspecified cell type|9800/3
C0023418|T191|HT|C95|ICD10CM|Leukemia of unspecified cell type|9800/3
C0023418|T191|AB|C95.9|ICD10CM|Leukemia, unspecified|9800/3
C0023418|T191|HT|C95.9|ICD10CM|Leukemia, unspecified|9800/3
C0023418|T191|HT|208|ICD9CM|Leukemia of unspecified cell type|9800/3
C0023418|T191|HT|208.9|ICD9CM|Unspecified leukemia|9800/3
C0023418|T191|PT|B73|ICPC|Leukemia|9800/3
C0023418|T191|AB|B73|ICPC2EENG|Leukaemia|9800/3
C0023418|T191|PT|B73|ICPC2EENG|Leukaemia|9800/3
C0023418|T191|PT|MTHU044737|ICPC2ICD10ENG|leukemia|9800/3
C0023418|T191|PTN|B73001|ICPC2P|leukaemia|9800/3
C0023418|T191|PT|B73001|ICPC2P|Leukaemia|9800/3
C0023418|T191|MTH_PT|B73001|ICPC2P|Leukemia|9800/3
C0023418|T191|MTH_PTN|B73001|ICPC2P|leukemia|9800/3
C0023418|T191|PT|U002665|LCH|Leukemia|9800/3
C0023418|T191|PT|sh85076285|LCH_NW|Leukemia|9800/3
C0023418|T191|LA|LA10545-4|LNC|Leukemia|9800/3
C0023418|T191|PT|10024288|MDR|Leukaemia|9800/3
C0023418|T191|LLT|10024288|MDR|Leukaemia|9800/3
C0023418|T191|LLT|10024312|MDR|Leukaemia NOS|9800/3
C0023418|T191|LLT|10024314|MDR|Leukaemia of unspecified cell type|9800/3
C0023418|T191|LLT|10024323|MDR|Leukaemia unspecified|9800/3
C0023418|T191|HG|10024324|MDR|Leukaemias|9800/3
C0023418|T191|LLT|10024329|MDR|Leukemia|9800/3
C0023418|T191|MTH_PT|10024288|MDR|Leukemia|9800/3
C0023418|T191|LLT|10024351|MDR|Leukemia NOS|9800/3
C0023418|T191|LLT|10024352|MDR|Leukemia of unspecified cell type|9800/3
C0023418|T191|LLT|10060500|MDR|Leukemia unspecified|9800/3
C0023418|T191|MTH_HG|10024324|MDR|Leukemias|9800/3
C0023418|T191|LLT|10045991|MDR|Unspecified leukaemia|9800/3
C0023418|T191|LLT|10060430|MDR|Unspecified leukaemia without mention of remission|9800/3
C0023418|T191|LLT|10045992|MDR|Unspecified leukemia|9800/3
C0023418|T191|LLT|10045994|MDR|Unspecified leukemia without mention of remission|9800/3
C0023418|T191|PT|31470|MEDCIN|leukemia|9800/3
C0023418|T191|PT|5620|MEDLINEPLUS|Leukemia|9800/3
C0023418|T191|ET|D007938|MSH|Leucocythaemia|9800/3
C0023418|T191|PM|D007938|MSH|Leucocythaemias|9800/3
C0023418|T191|ET|D007938|MSH|Leucocythemia|9800/3
C0023418|T191|PM|D007938|MSH|Leucocythemias|9800/3
C0023418|T191|MH|D007938|MSH|Leukemia|9800/3
C0023418|T191|PM|D007938|MSH|Leukemias|9800/3
C0023418|T191|SY|NOCODE|MTH|LEUKEMIA|9800/3
C0023418|T191|PN|NOCODE|MTH|leukemia|9800/3
C0023418|T191|ET|208.9|MTHICD9|Leukemia NOS|9800/3
C0023418|T191|PT|C3161|NCI|Leukemia|9800/3
C0023418|T191|SY|TCGA|NCI|Leukemia|9800/3
C0023418|T191|SY|C3161|NCI_CDISC|Leukemia NOS|9800/3
C0023418|T191|PT|C3161|NCI_CDISC|LEUKEMIA, MALIGNANT|9800/3
C0023418|T191|SY|C3161|NCI_CDISC|Leukemias|9800/3
C0023418|T191|SY|C3161|NCI_CDISC|Leukemias, General|9800/3
C0023418|T191|PT|C3161|NCI_CPTAC|Leukemia|9800/3
C0023418|T191|PT|10024312|NCI_CTEP-SDC|Leukemia, NOS|9800/3
C0023418|T191|PT|C3161|NCI_CTRP|Leukemia|9800/3
C0023418|T191|DN|C3161|NCI_CTRP|Leukemia|9800/3
C0023418|T191|PT|CDR0000045343|NCI_NCI-GLOSS|leukemia|9800/3
C0023418|T191|PT|C3161|NCI_NICHD|Leukemia|9800/3
C0023418|T191|SY|C3161|NCI_NICHD|Leukemia, Disease|9800/3
C0023418|T191|PT|CDR0000041186|PDQ|leukemia|9800/3
C0023418|T191|SY|CDR0000041186|PDQ|Leukemias|9800/3
C0023418|T191|SY|CDR0000041186|PDQ|Leukemias, General|9800/3
C0023418|T191|PT|28260|PSY|Leukemias|9800/3
C0023418|T191|OP|X78e2|RCD|Leukaemia|9800/3
C0023418|T191|PT|BBr..|RCD|Leukaemia morphology|9800/3
C0023418|T191|OP|B68z.|RCD|Leukaemia NOS|9800/3
C0023418|T191|OP|B68..|RCD|Leukaemia of unspecified cell type|9800/3
C0023418|T191|OA|B68..|RCD|Unspecif. cell type leukaemia|9800/3
C0023418|T191|OP|X78e2|RCDAE|Leukemia|9800/3
C0023418|T191|PT|BBr..|RCDAE|Leukemia morphology|9800/3
C0023418|T191|OP|B68z.|RCDAE|Leukemia NOS|9800/3
C0023418|T191|OP|B68..|RCDAE|Leukemia of unspecified cell type|9800/3
C0023418|T191|OA|B68..|RCDAE|Unspecif. cell type leukemia|9800/3
C0023418|T191|OP|BBr00|RCDSA|Leukemia NOS|9800/3
C0023418|T191|OP|BBr0z|RCDSA|Leukemia unspecified, NOS|9800/3
C0023418|T191|OP|BBr0.|RCDSA|Leukemias unspecified|9800/3
C0023418|T191|OP|BBr00|RCDSY|Leukaemia NOS|9800/3
C0023418|T191|OP|BBr0z|RCDSY|Leukaemia unspecified, NOS|9800/3
C0023418|T191|OP|BBr0.|RCDSY|Leukaemias unspecified|9800/3
C0023418|T191|PTGB|93143009|SNOMEDCT_US|Leukaemia|9800/3
C0023418|T191|PTGB|87163000|SNOMEDCT_US|Leukaemia|9800/3
C0023418|T191|OAP|255049003|SNOMEDCT_US|Leukaemia|9800/3
C1292766|T191|SYGB|128931003|SNOMEDCT_US|Leukaemia - category|9800/3
C0023418|T191|SYGB|87163000|SNOMEDCT_US|Leukaemia morphology|9800/3
C0023418|T191|OAP|188767008|SNOMEDCT_US|Leukaemia NOS|9800/3
C0023418|T191|OF|154598008|SNOMEDCT_US|Leukaemia of unspecified cell type|9800/3
C0023418|T191|OAP|154598008|SNOMEDCT_US|Leukaemia of unspecified cell type|9800/3
C0023418|T191|OAP|188762002|SNOMEDCT_US|Leukaemia of unspecified cell type|9800/3
C0023418|T191|SYGB|93143009|SNOMEDCT_US|Leukaemia, disease|9800/3
C0023418|T191|SYGB|87163000|SNOMEDCT_US|Leukaemia, no ICD-O subtype|9800/3
C0023418|T191|IS|87163000|SNOMEDCT_US|Leukaemia, NOS|9800/3
C0023418|T191|IS|93143009|SNOMEDCT_US|Leukaemia, NOS, without mention of remission|9800/3
C0023418|T191|OAP|255049003|SNOMEDCT_US|Leukemia|9800/3
C0023418|T191|PT|87163000|SNOMEDCT_US|Leukemia|9800/3
C0023418|T191|PT|93143009|SNOMEDCT_US|Leukemia|9800/3
C1292766|T191|SY|128931003|SNOMEDCT_US|Leukemia - category|9800/3
C0023418|T191|SY|87163000|SNOMEDCT_US|Leukemia morphology|9800/3
C0023418|T191|OAP|188767008|SNOMEDCT_US|Leukemia NOS|9800/3
C0023418|T191|OAP|154598008|SNOMEDCT_US|Leukemia of unspecified cell type|9800/3
C0023418|T191|OAP|188762002|SNOMEDCT_US|Leukemia of unspecified cell type|9800/3
C0023418|T191|SY|93143009|SNOMEDCT_US|Leukemia, disease|9800/3
C0023418|T191|SY|87163000|SNOMEDCT_US|Leukemia, no ICD-O subtype|9800/3
C0023418|T191|SY|87163000|SNOMEDCT_US|Leukemia, no International Classification of Diseases for Oncology subtype|9800/3
C0023418|T191|IS|87163000|SNOMEDCT_US|Leukemia, NOS|9800/3
C0023418|T191|IS|93143009|SNOMEDCT_US|Leukemia, NOS, without mention of remission|9800/3
C0023418|T191|HT|0573|WHO|LEUKAEMIA|9800/3
C0085669|T191|PT|0025555|CCPSS|LEUKEMIA ACUTE|9801/3
C0085669|T191|SY|0000015724|CHV|acute leukaemia|9801/3
C0085669|T191|SY|0000015724|CHV|acute leukaemias|9801/3
C0085669|T191|PT|0000015724|CHV|acute leukemia|9801/3
C0085669|T191|SY|0000015724|CHV|acute leukemias|9801/3
C0085669|T191|PT|U000010|COSTAR|ACUTE LEUKEMIA|9801/3
C0085669|T191|PT|2004-1600|CSP|acute leukemia|9801/3
C0085669|T191|PT|LEUKEMIA ACUTE|CST|ACUTE LEUKEMIA|9801/3
C0085669|T191|GT|LEUKEMIA ACUTE|CST|LEUKAEMIA ACUTE|9801/3
C0085669|T191|GT|LEUKEMIA ACUTE|CST|LEUKEMIA ACUTE|9801/3
C0085669|T191|PT|HP:0002488|HPO|Acute leukemia|9801/3
C0085669|T191|SY|HP:0002488|HPO|Acute leukemias|9801/3
C0085669|T191|PT|C95.0|ICD10|Acute leukaemia of unspecified cell type|9801/3
C0085669|T191|PT|C95.0|ICD10AE|Acute leukemia of unspecified cell type|9801/3
C0085669|T191|ET|C95.00|ICD10CM|Acute leukemia NOS|9801/3
C0085669|T191|AB|C95.0|ICD10CM|Acute leukemia of unspecified cell type|9801/3
C0085669|T191|HT|C95.0|ICD10CM|Acute leukemia of unspecified cell type|9801/3
C0085669|T191|HT|208.0|ICD9CM|Leukemia of unspecified cell type, acute|9801/3
C0085669|T191|PT|MTHU003149|ICPC2ICD10ENG|acute; leukemia|9801/3
C0085669|T191|PT|MTHU044738|ICPC2ICD10ENG|leukemia; acute|9801/3
C0085669|T191|LLT|10000830|MDR|Acute leukaemia|9801/3
C0085669|T191|PT|10000830|MDR|Acute leukaemia|9801/3
C0085669|T191|LLT|10000831|MDR|Acute leukaemia NOS|9801/3
C0085669|T191|LLT|10000833|MDR|Acute leukaemia of unspecified cell type|9801/3
C0085669|T191|MTH_PT|10000830|MDR|Acute leukemia|9801/3
C0085669|T191|LLT|10000835|MDR|Acute leukemia|9801/3
C0085669|T191|LLT|10000836|MDR|Acute leukemia NOS|9801/3
C0085669|T191|LLT|10060554|MDR|Acute leukemia of unspecified cell type|9801/3
C0085669|T191|LLT|10024289|MDR|Leukaemia acute|9801/3
C0085669|T191|LLT|10024315|MDR|Leukaemia of unspecified cell type, acute|9801/3
C0085669|T191|LLT|10024330|MDR|Leukemia acute|9801/3
C0085669|T191|LLT|10024353|MDR|Leukemia of unspecified cell type, acute|9801/3
C0085669|T191|PT|36061|MEDCIN|acute leukemia|9801/3
C1301357|T191|PT|366678|MEDCIN|Acute leukemia of ambiguous lineage|9801/3
C0085669|T191|SY|36061|MEDCIN|leukemia acute|9801/3
C1301357|T191|SY|366678|MEDCIN|leukemia acute ambiguous lineage|9801/3
C0085669|T191|PN|NOCODE|MTH|Acute leukemia|9801/3
C1301357|T191|PN|NOCODE|MTH|Acute Leukemia of Ambiguous Lineage|9801/3
C0085669|T191|SY|NOCODE|MTH|LEUKEMIA ACUTE|9801/3
C0085669|T191|ET|208.0|MTHICD9|Acute leukemia NOS|9801/3
C0085669|T191|PT|C9300|NCI|Acute Leukemia|9801/3
C1301357|T191|PT|C7464|NCI|Acute Leukemia of Ambiguous Lineage|9801/3
C1301357|T191|SY|TCGA|NCI|Acute Leukemia of Ambiguous Lineage|9801/3
C1301357|T191|SY|C7464|NCI|Acute Leukemia of Indeterminate Lineage|9801/3
C0085669|T191|PT|C9300|NCI_CPTAC|Acute Leukemia|9801/3
C0085669|T191|DN|C9300|NCI_CTRP|Acute Leukemia|9801/3
C1301357|T191|DN|C7464|NCI_CTRP|Acute Leukemia of Ambiguous Lineage|9801/3
C0085669|T191|PT|CDR0000045145|NCI_NCI-GLOSS|acute leukemia|9801/3
C1301357|T191|PT|C7464|NCI_NICHD|Acute Leukemia of Ambiguous Lineage|9801/3
C1301357|T191|SY|C7464|NCI_NICHD|Acute Leukemia of Indeterminate Lineage|9801/3
C0085669|T191|PT|CDR0000038952|PDQ|acute leukemia|9801/3
C0085669|T191|SY|CDR0000040510|PDQ|acute leukemia not otherwise specified|9801/3
C0085669|T191|SY|CDR0000040510|PDQ|acute leukemia, NOS|9801/3
C1301357|T191|PT|CDR0000670794|PDQ|acute leukemias of ambiguous lineage|9801/3
C0085669|T191|SY|CDR0000038952|PDQ|leukemia, acute|9801/3
C0085669|T191|SY|CDR0000040510|PDQ|stem cell acute leukemia|9801/3
C0085669|T191|PT|Xa9AM|RCD|Acute leukaemia|9801/3
C0085669|T191|OP|B680.|RCD|Acute leukaemia NOS|9801/3
C0085669|T191|PT|Xa9AM|RCDAE|Acute leukemia|9801/3
C0085669|T191|OP|B680.|RCDAE|Acute leukemia NOS|9801/3
C0085669|T191|OP|BBr01|RCDSA|Acute leukemia NOS|9801/3
C0085669|T191|OP|BBr01|RCDSY|Acute leukaemia NOS|9801/3
C0085669|T191|PTGB|24072005|SNOMEDCT_US|Acute leukaemia|9801/3
C0085669|T191|PTGB|91855006|SNOMEDCT_US|Acute leukaemia|9801/3
C1292764|T191|SYGB|128932005|SNOMEDCT_US|Acute leukaemia - category|9801/3
C0085669|T191|OAP|154599000|SNOMEDCT_US|Acute leukaemia NOS|9801/3
C0085669|T191|OAP|188763007|SNOMEDCT_US|Acute leukaemia NOS|9801/3
C0085669|T191|OF|154599000|SNOMEDCT_US|Acute leukaemia NOS|9801/3
C1301357|T191|PTGB|721308005|SNOMEDCT_US|Acute leukaemia of ambiguous lineage|9801/3
C1301357|T191|PTGB|397345009|SNOMEDCT_US|Acute leukaemia of ambiguous lineage|9801/3
C0085669|T191|SYGB|91855006|SNOMEDCT_US|Acute leukaemia, disease|9801/3
C0085669|T191|SYGB|24072005|SNOMEDCT_US|Acute leukaemia, morphology, including blast cell OR undifferentiated leukaemia|9801/3
C0085669|T191|PT|24072005|SNOMEDCT_US|Acute leukemia|9801/3
C0085669|T191|PT|91855006|SNOMEDCT_US|Acute leukemia|9801/3
C1292764|T191|SY|128932005|SNOMEDCT_US|Acute leukemia - category|9801/3
C0085669|T191|OAP|154599000|SNOMEDCT_US|Acute leukemia NOS|9801/3
C0085669|T191|OAP|188763007|SNOMEDCT_US|Acute leukemia NOS|9801/3
C1301357|T191|PT|721308005|SNOMEDCT_US|Acute leukemia of ambiguous lineage|9801/3
C1301357|T191|PT|397345009|SNOMEDCT_US|Acute leukemia of ambiguous lineage|9801/3
C0085669|T191|SY|91855006|SNOMEDCT_US|Acute leukemia, disease|9801/3
C0085669|T191|SY|24072005|SNOMEDCT_US|Acute leukemia, morphology, including blast cell OR undifferentiated leukemia|9801/3
C0085669|T191|IS|24072005|SNOMEDCT_US|Acute leukemia, NOS|9801/3
C0085669|T191|PT|0574|WHO|LEUKAEMIA ACUTE|9801/3
C0023464|T191|SY|HP:0005531|HPO|Acute biphenotypic leukemia|9805/3
C0023464|T191|PT|HP:0005531|HPO|Biphenotypic acute leukaemia|9805/3
C0023464|T191|SY|HP:0005531|HPO|Myeloid/lymphoid leukemia|9805/3
C0023464|T191|ET|C95.0|ICD10CM|Acute mixed lineage leukemia|9805/3
C0023464|T191|ET|C95.0|ICD10CM|Biphenotypic acute leukemia|9805/3
C0023464|T191|PT|10067399|MDR|Acute biphenotypic leukaemia|9805/3
C0023464|T191|LLT|10067399|MDR|Acute biphenotypic leukaemia|9805/3
C0023464|T191|LLT|10067837|MDR|Acute biphenotypic leukemia|9805/3
C0023464|T191|MTH_PT|10067399|MDR|Acute biphenotypic leukemia|9805/3
C0023464|T191|PT|230904|MEDCIN|acute biphenotypic leukemia|9805/3
C0023464|T191|SY|230904|MEDCIN|leukemia acute biphenotypic|9805/3
C0023464|T191|ET|D015456|MSH|Acute Biphenotypic Leukemia|9805/3
C0023464|T191|PM|D015456|MSH|Acute Biphenotypic Leukemias|9805/3
C0023464|T191|PM|D015456|MSH|Acute Leukemia, Biphenotypic|9805/3
C0023464|T191|PM|D015456|MSH|Acute Leukemia, Hybrid|9805/3
C0023464|T191|PM|D015456|MSH|Acute Leukemia, Mixed-Lineage|9805/3
C0023464|T191|PM|D015456|MSH|Acute Leukemias, Biphenotypic|9805/3
C0023464|T191|PM|D015456|MSH|Acute Leukemias, Hybrid|9805/3
C0023464|T191|PM|D015456|MSH|Acute Leukemias, Mixed-Lineage|9805/3
C0023464|T191|DSV|D015456|MSH|B AND T CELL ACUTE LYMPHOBLASTIC LEUKEMIA|9805/3
C0023464|T191|ET|D015456|MSH|B and T Cell Acute Lymphoblastic Leukemia|9805/3
C0023464|T191|DSV|D015456|MSH|B AND T CELL LEUKEMIA ACUTE|9805/3
C0023464|T191|ET|D015456|MSH|B and T Cell Leukemia, Acute|9805/3
C0023464|T191|ET|D015456|MSH|B- and T-Cell Acute Lymphoblastic Leukemia|9805/3
C0023464|T191|ET|D015456|MSH|B- and T-Cell Leukemia, Acute|9805/3
C0023464|T191|ET|D015456|MSH|Biphenotypic Acute Leukemia|9805/3
C0023464|T191|PM|D015456|MSH|Biphenotypic Acute Leukemias|9805/3
C0023464|T191|PM|D015456|MSH|Biphenotypic Leukemia, Acute|9805/3
C0023464|T191|PM|D015456|MSH|Biphenotypic Leukemias, Acute|9805/3
C0023464|T191|PM|D015456|MSH|Hybrid Acute Leukemia|9805/3
C0023464|T191|ET|D015456|MSH|Hybrid Acute Leukemias|9805/3
C0023464|T191|DSV|D015456|MSH|LEUKEMIA MIXED B AND T CELL|9805/3
C0023464|T191|PM|D015456|MSH|Leukemia, Acute Biphenotypic|9805/3
C0023464|T191|PM|D015456|MSH|Leukemia, Biphenotypic Acute|9805/3
C0023464|T191|MH|D015456|MSH|Leukemia, Biphenotypic, Acute|9805/3
C0023464|T191|PM|D015456|MSH|Leukemia, Hybrid Acute|9805/3
C0023464|T191|ET|D015456|MSH|Leukemia, Lymphocytic, Acute, Mixed Cell|9805/3
C0023464|T191|ET|D015456|MSH|Leukemia, Lymphocytic, Acute, Mixed-Cell|9805/3
C0023464|T191|PM|D015456|MSH|Leukemia, Mixed Cell|9805/3
C0023464|T191|ET|D015456|MSH|Leukemia, Mixed-Cell|9805/3
C0023464|T191|PM|D015456|MSH|Leukemia, Mixed-Lineage Acute|9805/3
C0023464|T191|ET|D015456|MSH|Leukemia, Mixed, B and T Cell|9805/3
C0023464|T191|ET|D015456|MSH|Leukemia, Mixed, B- and T-Cell|9805/3
C0023464|T191|PM|D015456|MSH|Leukemias, Acute Biphenotypic|9805/3
C0023464|T191|PM|D015456|MSH|Leukemias, Biphenotypic Acute|9805/3
C0023464|T191|PM|D015456|MSH|Leukemias, Hybrid Acute|9805/3
C0023464|T191|PM|D015456|MSH|Leukemias, Mixed-Cell|9805/3
C0023464|T191|PM|D015456|MSH|Leukemias, Mixed-Lineage Acute|9805/3
C0023464|T191|DSV|D015456|MSH|LYMPHOCYTIC LEUKEMIA ACUTE B AND T CELL|9805/3
C0023464|T191|ET|D015456|MSH|Lymphocytic Leukemia, Acute, B and T Cell|9805/3
C0023464|T191|ET|D015456|MSH|Lymphocytic Leukemia, Acute, B- and T-Cell|9805/3
C0023464|T191|PM|D015456|MSH|Mixed Lineage Acute Leukemias|9805/3
C0023464|T191|PM|D015456|MSH|Mixed-Cell Leukemia|9805/3
C0023464|T191|PM|D015456|MSH|Mixed-Cell Leukemias|9805/3
C0023464|T191|PM|D015456|MSH|Mixed-Lineage Acute Leukemia|9805/3
C0023464|T191|ET|D015456|MSH|Mixed-Lineage Acute Leukemias|9805/3
C0023464|T191|PN|NOCODE|MTH|Acute biphenotypic leukemia|9805/3
C2826025|T191|PN|NOCODE|MTH|Mixed phenotype acute leukemia|9805/3
C0023464|T191|PT|C4673|NCI|Acute Biphenotypic Leukemia|9805/3
C0023464|T191|SY|TCGA|NCI|Acute Biphenotypic Leukemia|9805/3
C2826025|T191|PT|C82179|NCI|Mixed Phenotype Acute Leukemia|9805/3
C2826025|T191|AB|C82179|NCI|MPAL|9805/3
C0023464|T191|DN|C4673|NCI_CTRP|Acute Biphenotypic Leukemia|9805/3
C2826025|T191|DN|C82179|NCI_CTRP|Mixed Phenotype Acute Leukemia|9805/3
C0023464|T191|PT|C4673|NCI_NICHD|Acute Biphenotypic Leukemia|9805/3
C2826025|T191|PT|C82179|NCI_NICHD|Mixed Phenotype Acute Leukemia|9805/3
C2826025|T191|SY|C82179|NCI_NICHD|MPAL|9805/3
C0023464|T191|PT|Xa0jn|RCD|Acute biphenotypic leukaemia|9805/3
C0023464|T191|PT|Xa0jn|RCDAE|Acute biphenotypic leukemia|9805/3
C0023464|T191|PTGB|278453007|SNOMEDCT_US|Acute biphenotypic leukaemia|9805/3
C0023464|T191|PTGB|128818009|SNOMEDCT_US|Acute biphenotypic leukaemia|9805/3
C0023464|T191|PT|128818009|SNOMEDCT_US|Acute biphenotypic leukemia|9805/3
C0023464|T191|PT|278453007|SNOMEDCT_US|Acute biphenotypic leukemia|9805/3
C0023464|T191|IS|128818009|SNOMEDCT_US|Acute mixed lineage leukaemia|9805/3
C2826025|T191|SYGB|450913003|SNOMEDCT_US|Acute mixed lineage leukaemia|9805/3
C2826025|T191|SY|450913003|SNOMEDCT_US|Acute mixed lineage leukemia|9805/3
C0023464|T191|IS|128818009|SNOMEDCT_US|Acute mixed lineage leukemia|9805/3
C2826025|T191|PTGB|450913003|SNOMEDCT_US|Mixed phenotype acute leukaemia|9805/3
C2826025|T191|PT|450913003|SNOMEDCT_US|Mixed phenotype acute leukemia|9805/3
C3472616|T191|SY|C82212|NCI|Mixed Phenotype Acute Leukemia, B/Myeloid, NOS|9808/3
C3472616|T191|PT|C82212|NCI|Mixed Phenotype Acute Leukemia, B/Myeloid, Not Otherwise Specified|9808/3
C3472616|T191|OP|450916006|SNOMEDCT_US|Mixed phenotype acute leukaemia B/lymphoid|9808/3
C3472616|T191|PTGB|450916006|SNOMEDCT_US|Mixed phenotype acute leukaemia B/myeloid|9808/3
C3472616|T191|SYGB|450916006|SNOMEDCT_US|Mixed phenotype acute leukaemia with myeloid and B-cell lymphoid phenotypes|9808/3
C3472616|T191|OP|450916006|SNOMEDCT_US|Mixed phenotype acute leukemia B/lymphoid|9808/3
C3472616|T191|PT|450916006|SNOMEDCT_US|Mixed phenotype acute leukemia B/myeloid|9808/3
C3472616|T191|SY|450916006|SNOMEDCT_US|Mixed phenotype acute leukemia with myeloid and B-cell lymphoid phenotypes|9808/3
C2826055|T191|SY|C82213|NCI|Mixed Phenotype Acute Leukemia, T/Myeloid, NOS|9809/3
C2826055|T191|PT|C82213|NCI|Mixed Phenotype Acute Leukemia, T/Myeloid, Not Otherwise Specified|9809/3
C2826055|T191|PTGB|450917002|SNOMEDCT_US|Mixed phenotype acute leukaemia T/myeloid|9809/3
C2826055|T191|SYGB|450917002|SNOMEDCT_US|Mixed phenotype acute leukaemia with myeloid and T-cell lymphoid pheotypes|9809/3
C2826055|T191|PT|450917002|SNOMEDCT_US|Mixed phenotype acute leukemia T/myeloid|9809/3
C2826055|T191|SY|450917002|SNOMEDCT_US|Mixed phenotype acute leukemia with myeloid and T-cell lymphoid phenotypes|9809/3
C0023448|T191|ET|0000004619|AOD|lymphocytic leukemia|981-983
C0023448|T191|SY|0000007336|CHV|leukemia lymphoblastic|981-983
C0023448|T191|SY|0000007336|CHV|leukemia lymphocytic|981-983
C0023448|T191|SY|0000007336|CHV|leukemia lymphoid|981-983
C0023448|T191|SY|0000007336|CHV|lymphatic leukaemia|981-983
C0023448|T191|SY|0000007336|CHV|lymphatic leukemia|981-983
C0023448|T191|SY|0000007336|CHV|lymphoblastic leukemia|981-983
C0023448|T191|SY|0000007336|CHV|lymphocytic leukaemia|981-983
C0023448|T191|PT|0000007336|CHV|lymphocytic leukemia|981-983
C0023448|T191|SY|0000007336|CHV|lymphoid leukaemia|981-983
C0023448|T191|SY|0000007336|CHV|lymphoid leukemia|981-983
C0023448|T191|PT|U000428|COSTAR|LYMPHOCYTIC LEUKEMIA|981-983
C0023448|T191|ET|2004-2462|CSP|lymphatic leukemia|981-983
C0023448|T191|ET|2004-2462|CSP|lymphoblastic leukemia|981-983
C0023448|T191|PT|2004-2462|CSP|lymphocytic leukemia|981-983
C0023448|T191|ET|2004-2462|CSP|lymphogenous leukemia|981-983
C0023448|T191|ET|2004-2462|CSP|lymphoid leukemia|981-983
C0023448|T191|GT|LEUKEMIA CHRON LYMPHO|CST|LEUKAEMIA LYMPHOCYTIC|981-983
C0023448|T191|GT|LEUKEMIA CHRON LYMPHO|CST|LEUKEMIA LYMPHATIC|981-983
C0023448|T191|GT|LEUKEMIA CHRON LYMPHO|CST|LEUKEMIA LYMPHOID|981-983
C0023448|T191|PT|HP:0005526|HPO|Lymphoid leukemia|981-983
C0023448|T191|HT|C91|ICD10|Lymphoid leukaemia|981-983
C0023448|T191|PT|C91.9|ICD10|Lymphoid leukaemia, unspecified|981-983
C0023448|T191|HT|C91|ICD10AE|Lymphoid leukemia|981-983
C0023448|T191|PT|C91.9|ICD10AE|Lymphoid leukemia, unspecified|981-983
C0023448|T191|HT|C91|ICD10CM|Lymphoid leukemia|981-983
C0023448|T191|AB|C91|ICD10CM|Lymphoid leukemia|981-983
C0023448|T191|ET|C91.90|ICD10CM|Lymphoid leukemia NOS|981-983
C0023448|T191|AB|C91.9|ICD10CM|Lymphoid leukemia, unspecified|981-983
C0023448|T191|HT|C91.9|ICD10CM|Lymphoid leukemia, unspecified|981-983
C0023448|T191|HT|204|ICD9CM|Lymphoid leukemia|981-983
C0023448|T191|HT|204.9|ICD9CM|Unspecified lymphoid leukemia|981-983
C0023448|T191|PT|MTHU044761|ICPC2ICD10ENG|leukemia; lymphatic|981-983
C0023448|T191|PT|MTHU044766|ICPC2ICD10ENG|leukemia; lymphoblastic|981-983
C0023448|T191|PT|MTHU046611|ICPC2ICD10ENG|lymphatic; leukemia|981-983
C0023448|T191|PT|MTHU046684|ICPC2ICD10ENG|lymphoblastic; leukemia|981-983
C0023448|T191|PT|sh85079150|LCH_NW|Lymphocytic leukemia|981-983
C0023448|T191|LLT|10024301|MDR|Leukaemia lymphatic|981-983
C0023448|T191|LLT|10024302|MDR|Leukaemia lymphocytic|981-983
C0023448|T191|LLT|10024304|MDR|Leukaemia lymphoid|981-983
C0023448|T191|LLT|10024337|MDR|Leukemia lymphatic|981-983
C0023448|T191|LLT|10024339|MDR|Leukemia lymphocytic|981-983
C0023448|T191|LLT|10024341|MDR|Leukemia lymphoid|981-983
C0023448|T191|LLT|10060397|MDR|Lymphatic leukaemia|981-983
C0023448|T191|LLT|10025230|MDR|Lymphatic leukemia|981-983
C0023448|T191|LLT|10025234|MDR|Lymphoblastic leukaemia NOS|981-983
C0023448|T191|LLT|10025235|MDR|Lymphoblastic leukemia NOS|981-983
C0023448|T191|PT|10025270|MDR|Lymphocytic leukaemia|981-983
C0023448|T191|LLT|10025270|MDR|Lymphocytic leukaemia|981-983
C0023448|T191|LLT|10025271|MDR|Lymphocytic leukemia|981-983
C0023448|T191|MTH_PT|10025270|MDR|Lymphocytic leukemia|981-983
C0023448|T191|LLT|10025299|MDR|Lymphoid leukaemia|981-983
C0023448|T191|LLT|10025304|MDR|Lymphoid leukemia|981-983
C0023448|T191|LLT|10045996|MDR|Unspecified lymphoid leukaemia|981-983
C0023448|T191|LLT|10045997|MDR|Unspecified lymphoid leukemia|981-983
C0023448|T191|SY|99743|MEDCIN|leukemia lymphocytic|981-983
C0023448|T191|PT|99743|MEDCIN|lymphocytic leukemia|981-983
C0023448|T191|ET|D007945|MSH|Leukemia, Lymphocytic|981-983
C0023448|T191|MH|D007945|MSH|Leukemia, Lymphoid|981-983
C0023448|T191|PM|D007945|MSH|Leukemias, Lymphocytic|981-983
C0023448|T191|PM|D007945|MSH|Leukemias, Lymphoid|981-983
C0023448|T191|ET|D007945|MSH|Lymphocytic Leukemia|981-983
C0023448|T191|PM|D007945|MSH|Lymphocytic Leukemias|981-983
C0023448|T191|ET|D007945|MSH|Lymphoid Leukemia|981-983
C0023448|T191|PM|D007945|MSH|Lymphoid Leukemias|981-983
C0023448|T191|SY|NOCODE|MTH|LEUKEMIA LYMPHATIC|981-983
C0023448|T191|SY|NOCODE|MTH|LEUKEMIA LYMPHOCYTIC|981-983
C0023448|T191|SY|NOCODE|MTH|LEUKEMIA LYMPHOID|981-983
C0023448|T191|PN|NOCODE|MTH|Lymphoid leukemia|981-983
C0023448|T191|SY|C7539|NCI|Lymphocytic Leukemia|981-983
C0023448|T191|SY|C7539|NCI|Lymphogenous Leukemia|981-983
C0023448|T191|PT|C7539|NCI|Lymphoid Leukemia|981-983
C0023448|T191|PT|C7539|NCI_CDISC|LEUKEMIA, LYMPHOCYTIC, MALIGNANT|981-983
C0023448|T191|SY|C7539|NCI_CDISC|Lymphocytic Leukemia|981-983
C0023448|T191|SY|C7539|NCI_CDISC|Lymphogenous Leukemia|981-983
C0023448|T191|PT|C7539|NCI_CPTAC|Lymphoid Leukemia|981-983
C0023448|T191|PT|C7539|NCI_CTRP|Lymphoid Leukemia|981-983
C0023448|T191|DN|C7539|NCI_CTRP|Lymphoid Leukemia|981-983
C0023448|T191|PT|CDR0000330173|NCI_NCI-GLOSS|lymphocytic leukemia|981-983
C0023448|T191|SY|B64..|RCD|Lymphatic leukaemia|981-983
C0023448|T191|PT|B64..|RCD|Lymphoid leukaemia|981-983
C0023448|T191|OP|B64z.|RCD|Lymphoid leukaemia NOS|981-983
C0023448|T191|SY|B64..|RCDAE|Lymphatic leukemia|981-983
C0023448|T191|PT|B64..|RCDAE|Lymphoid leukemia|981-983
C0023448|T191|OP|B64z.|RCDAE|Lymphoid leukemia NOS|981-983
C0023448|T191|OP|BBr20|RCDSA|Lymphoid leukemia NOS|981-983
C0023448|T191|PT|BBr2.|RCDSA|Lymphoid leukemias|981-983
C0023448|T191|OP|BBr20|RCDSY|Lymphoid leukaemia NOS|981-983
C0023448|T191|PT|BBr2.|RCDSY|Lymphoid leukaemias|981-983
C0023448|T191|SYGB|32280000|SNOMEDCT_US|Lymphatic leukaemia|981-983
C0023448|T191|SYGB|188725004|SNOMEDCT_US|Lymphatic leukaemia|981-983
C0023448|T191|SY|32280000|SNOMEDCT_US|Lymphatic leukemia|981-983
C0023448|T191|SY|188725004|SNOMEDCT_US|Lymphatic leukemia|981-983
C0023448|T191|IS|32280000|SNOMEDCT_US|Lymphatic leukemia, NOS|981-983
C0023448|T191|SYGB|32280000|SNOMEDCT_US|Lymphocytic leukaemia|981-983
C0023448|T191|SY|32280000|SNOMEDCT_US|Lymphocytic leukemia|981-983
C0023448|T191|IS|32280000|SNOMEDCT_US|Lymphocytic leukemia, NOS|981-983
C0023448|T191|OAP|93170002|SNOMEDCT_US|Lymphoid leukaemia|981-983
C0023448|T191|OAS|269631008|SNOMEDCT_US|Lymphoid leukaemia|981-983
C0023448|T191|OAS|154587007|SNOMEDCT_US|Lymphoid leukaemia|981-983
C0023448|T191|PTGB|32280000|SNOMEDCT_US|Lymphoid leukaemia|981-983
C0023448|T191|PTGB|188725004|SNOMEDCT_US|Lymphoid leukaemia|981-983
C0023448|T191|OAP|188731001|SNOMEDCT_US|Lymphoid leukaemia NOS|981-983
C0023448|T191|SYGB|32280000|SNOMEDCT_US|Lymphoid leukaemia, no ICD-O subtype|981-983
C0023448|T191|PT|188725004|SNOMEDCT_US|Lymphoid leukemia|981-983
C0023448|T191|PT|32280000|SNOMEDCT_US|Lymphoid leukemia|981-983
C0023448|T191|OAP|93170002|SNOMEDCT_US|Lymphoid leukemia|981-983
C0023448|T191|OAS|154587007|SNOMEDCT_US|Lymphoid leukemia|981-983
C0023448|T191|OAS|269631008|SNOMEDCT_US|Lymphoid leukemia|981-983
C0023448|T191|OAP|188731001|SNOMEDCT_US|Lymphoid leukemia NOS|981-983
C0023448|T191|SY|32280000|SNOMEDCT_US|Lymphoid leukemia, no ICD-O subtype|981-983
C0023448|T191|SY|32280000|SNOMEDCT_US|Lymphoid leukemia, no International Classification of Diseases for Oncology subtype|981-983
C0023448|T191|IS|32280000|SNOMEDCT_US|Lymphoid leukemia, NOS|981-983
C0023448|T191|IT|0176|WHO|LEUKAEMIA LYMPHATIC|981-983
C0023448|T191|PT|0176|WHO|LEUKAEMIA LYMPHOCYTIC|981-983
C0023448|T191|IT|0176|WHO|LEUKAEMIA LYMPHOID|981-983
C2698310|T191|SY|C80326|NCI|B Lymphoblastic Leukemia/Lymphoma, NOS|9811/3
C2698310|T191|PT|C80326|NCI|B Lymphoblastic Leukemia/Lymphoma, Not Otherwise Specified|9811/3
C4329384|T191|SY|C130039|NCI|B-Lymphoblastic Leukemia/Lymphoma with iAMP21|9811/3
C4329384|T191|PT|C130039|NCI|B-Lymphoblastic Leukemia/Lymphoma with Intrachromosomal Amplification of Chromosome 21|9811/3
C2698310|T191|SY|C80326|NCI|B-Lymphoblastic Leukemia/Lymphoma, Not Otherwise Specified|9811/3
C4329384|T191|PTGB|785825000|SNOMEDCT_US|B lymphoblastic leukaemia lymphoma with iAMP21|9811/3
C4329384|T191|SYGB|785825000|SNOMEDCT_US|B lymphoblastic leukaemia lymphoma with intrachromosomal amplification of chromosome 21|9811/3
C3472624|T191|PTGB|450949002|SNOMEDCT_US|B lymphoblastic leukaemia lymphoma, no ICD-O subtype|9811/3
C4329384|T191|PT|785825000|SNOMEDCT_US|B lymphoblastic leukemia lymphoma with iAMP21|9811/3
C4329384|T191|SY|785825000|SNOMEDCT_US|B lymphoblastic leukemia lymphoma with intrachromosomal amplification of chromosome 21|9811/3
C3472624|T191|PT|450949002|SNOMEDCT_US|B lymphoblastic leukemia lymphoma, no ICD-O subtype|9811/3
C3472624|T191|SY|450949002|SNOMEDCT_US|B lymphoblastic leukemia lymphoma, no International Classification of Diseases for Oncology subtype|9811/3
C1709527|T191|PT|HP:0004848|HPO|Ph-positive acute lymphoblastic leukemia|9812/3
C1709527|T191|SY|HP:0004848|HPO|Philadelphia-positive acute lymphoblastic leukemia|9812/3
C1709527|T191|SY|339905|MEDCIN|leukemia lymphocytic acute philadelphia chromosome-positive lymphoblastic|9812/3
C1709527|T191|PT|339905|MEDCIN|Philadelphia chromosome-positive acute lymphoblastic leukemia|9812/3
C1709527|T191|SY|C36312|NCI|Acute Lymphoblastic Leukemia, Philadelphia Chromosome Positive|9812/3
C1709527|T191|SY|C36312|NCI|Philadelphia Positive Acute Lymphoblastic Leukemia|9812/3
C1709527|T191|SY|C36312|NCI|Philadelphia Positive Precursor Lymphoblastic Leukemia|9812/3
C1709527|T191|SY|425688002|SNOMEDCT_US|Ph positive ALL|9812/3
C1709527|T191|SY|426955004|SNOMEDCT_US|Ph positive ALL|9812/3
C1709527|T191|SYGB|426955004|SNOMEDCT_US|Ph+ acute lymphoblastic leukaemia|9812/3
C1709527|T191|SYGB|425688002|SNOMEDCT_US|Ph+ acute lymphoblastic leukaemia|9812/3
C1709527|T191|SY|425688002|SNOMEDCT_US|Ph+ acute lymphoblastic leukemia|9812/3
C1709527|T191|SY|426955004|SNOMEDCT_US|Ph+ acute lymphoblastic leukemia|9812/3
C1709527|T191|SY|426955004|SNOMEDCT_US|Ph+ ALL|9812/3
C1709527|T191|SY|425688002|SNOMEDCT_US|Ph+ ALL|9812/3
C1709527|T191|PTGB|426955004|SNOMEDCT_US|Philadelphia chromosome-positive acute lymphoblastic leukaemia|9812/3
C1709527|T191|PTGB|425688002|SNOMEDCT_US|Philadelphia chromosome-positive acute lymphoblastic leukaemia|9812/3
C1709527|T191|PT|426955004|SNOMEDCT_US|Philadelphia chromosome-positive acute lymphoblastic leukemia|9812/3
C1709527|T191|PT|425688002|SNOMEDCT_US|Philadelphia chromosome-positive acute lymphoblastic leukemia|9812/3
C2698311|T191|PT|C80335|NCI|B Lymphoblastic Leukemia/Lymphoma with Hyperdiploidy|9815/3
C2698311|T191|SY|C80335|NCI|B-Lymphoblastic Leukemia/Lymphoma with Hyperdiploidy|9815/3
C2698311|T191|PTGB|450953000|SNOMEDCT_US|B lymphoblastic leukaemia lymphoma with hyperdiploidy|9815/3
C2698311|T191|PT|450953000|SNOMEDCT_US|B lymphoblastic leukemia lymphoma with hyperdiploidy|9815/3
C2698312|T191|PT|C80338|NCI|B Lymphoblastic Leukemia/Lymphoma with Hypodiploidy|9816/3
C2698312|T191|SY|C80338|NCI|B-Lymphoblastic Leukemia/Lymphoma with Hypodiploidy|9816/3
C0023448|T191|ET|0000004619|AOD|lymphocytic leukemia|9820/3
C0023448|T191|SY|0000007336|CHV|leukemia lymphoblastic|9820/3
C0023448|T191|SY|0000007336|CHV|leukemia lymphocytic|9820/3
C0023448|T191|SY|0000007336|CHV|leukemia lymphoid|9820/3
C0023448|T191|SY|0000007336|CHV|lymphatic leukaemia|9820/3
C0023448|T191|SY|0000007336|CHV|lymphatic leukemia|9820/3
C0023448|T191|SY|0000007336|CHV|lymphoblastic leukemia|9820/3
C0023448|T191|SY|0000007336|CHV|lymphocytic leukaemia|9820/3
C0023448|T191|PT|0000007336|CHV|lymphocytic leukemia|9820/3
C0023448|T191|SY|0000007336|CHV|lymphoid leukaemia|9820/3
C0023448|T191|SY|0000007336|CHV|lymphoid leukemia|9820/3
C0023448|T191|PT|U000428|COSTAR|LYMPHOCYTIC LEUKEMIA|9820/3
C0023448|T191|ET|2004-2462|CSP|lymphatic leukemia|9820/3
C0023448|T191|ET|2004-2462|CSP|lymphoblastic leukemia|9820/3
C0023448|T191|PT|2004-2462|CSP|lymphocytic leukemia|9820/3
C0023448|T191|ET|2004-2462|CSP|lymphogenous leukemia|9820/3
C0023448|T191|ET|2004-2462|CSP|lymphoid leukemia|9820/3
C0023448|T191|GT|LEUKEMIA CHRON LYMPHO|CST|LEUKAEMIA LYMPHOCYTIC|9820/3
C0023448|T191|GT|LEUKEMIA CHRON LYMPHO|CST|LEUKEMIA LYMPHATIC|9820/3
C0023448|T191|GT|LEUKEMIA CHRON LYMPHO|CST|LEUKEMIA LYMPHOID|9820/3
C0023448|T191|PT|HP:0005526|HPO|Lymphoid leukemia|9820/3
C0023448|T191|HT|C91|ICD10|Lymphoid leukaemia|9820/3
C0023448|T191|PT|C91.9|ICD10|Lymphoid leukaemia, unspecified|9820/3
C0023448|T191|HT|C91|ICD10AE|Lymphoid leukemia|9820/3
C0023448|T191|PT|C91.9|ICD10AE|Lymphoid leukemia, unspecified|9820/3
C0023448|T191|AB|C91|ICD10CM|Lymphoid leukemia|9820/3
C0023448|T191|HT|C91|ICD10CM|Lymphoid leukemia|9820/3
C0023448|T191|ET|C91.90|ICD10CM|Lymphoid leukemia NOS|9820/3
C0023448|T191|AB|C91.9|ICD10CM|Lymphoid leukemia, unspecified|9820/3
C0023448|T191|HT|C91.9|ICD10CM|Lymphoid leukemia, unspecified|9820/3
C0023448|T191|HT|204|ICD9CM|Lymphoid leukemia|9820/3
C0023448|T191|HT|204.9|ICD9CM|Unspecified lymphoid leukemia|9820/3
C0023448|T191|PT|MTHU044761|ICPC2ICD10ENG|leukemia; lymphatic|9820/3
C0023448|T191|PT|MTHU044766|ICPC2ICD10ENG|leukemia; lymphoblastic|9820/3
C0023448|T191|PT|MTHU046611|ICPC2ICD10ENG|lymphatic; leukemia|9820/3
C0023448|T191|PT|MTHU046684|ICPC2ICD10ENG|lymphoblastic; leukemia|9820/3
C0023448|T191|PT|sh85079150|LCH_NW|Lymphocytic leukemia|9820/3
C0023448|T191|LLT|10024301|MDR|Leukaemia lymphatic|9820/3
C0023448|T191|LLT|10024302|MDR|Leukaemia lymphocytic|9820/3
C0023448|T191|LLT|10024304|MDR|Leukaemia lymphoid|9820/3
C0023448|T191|LLT|10024337|MDR|Leukemia lymphatic|9820/3
C0023448|T191|LLT|10024339|MDR|Leukemia lymphocytic|9820/3
C0023448|T191|LLT|10024341|MDR|Leukemia lymphoid|9820/3
C0023448|T191|LLT|10060397|MDR|Lymphatic leukaemia|9820/3
C0023448|T191|LLT|10025230|MDR|Lymphatic leukemia|9820/3
C0023448|T191|LLT|10025234|MDR|Lymphoblastic leukaemia NOS|9820/3
C0023448|T191|LLT|10025235|MDR|Lymphoblastic leukemia NOS|9820/3
C0023448|T191|LLT|10025270|MDR|Lymphocytic leukaemia|9820/3
C0023448|T191|PT|10025270|MDR|Lymphocytic leukaemia|9820/3
C0023448|T191|LLT|10025271|MDR|Lymphocytic leukemia|9820/3
C0023448|T191|MTH_PT|10025270|MDR|Lymphocytic leukemia|9820/3
C0023448|T191|LLT|10025299|MDR|Lymphoid leukaemia|9820/3
C0023448|T191|LLT|10025304|MDR|Lymphoid leukemia|9820/3
C0023448|T191|LLT|10045996|MDR|Unspecified lymphoid leukaemia|9820/3
C0023448|T191|LLT|10045997|MDR|Unspecified lymphoid leukemia|9820/3
C0023448|T191|SY|99743|MEDCIN|leukemia lymphocytic|9820/3
C0023448|T191|PT|99743|MEDCIN|lymphocytic leukemia|9820/3
C0023448|T191|ET|D007945|MSH|Leukemia, Lymphocytic|9820/3
C0023448|T191|MH|D007945|MSH|Leukemia, Lymphoid|9820/3
C0023448|T191|PM|D007945|MSH|Leukemias, Lymphocytic|9820/3
C0023448|T191|PM|D007945|MSH|Leukemias, Lymphoid|9820/3
C0023448|T191|ET|D007945|MSH|Lymphocytic Leukemia|9820/3
C0023448|T191|PM|D007945|MSH|Lymphocytic Leukemias|9820/3
C0023448|T191|ET|D007945|MSH|Lymphoid Leukemia|9820/3
C0023448|T191|PM|D007945|MSH|Lymphoid Leukemias|9820/3
C0023448|T191|SY|NOCODE|MTH|LEUKEMIA LYMPHATIC|9820/3
C0023448|T191|SY|NOCODE|MTH|LEUKEMIA LYMPHOCYTIC|9820/3
C0023448|T191|SY|NOCODE|MTH|LEUKEMIA LYMPHOID|9820/3
C0023448|T191|PN|NOCODE|MTH|Lymphoid leukemia|9820/3
C0023448|T191|SY|C7539|NCI|Lymphocytic Leukemia|9820/3
C0023448|T191|SY|C7539|NCI|Lymphogenous Leukemia|9820/3
C0023448|T191|PT|C7539|NCI|Lymphoid Leukemia|9820/3
C0023448|T191|PT|C7539|NCI_CDISC|LEUKEMIA, LYMPHOCYTIC, MALIGNANT|9820/3
C0023448|T191|SY|C7539|NCI_CDISC|Lymphocytic Leukemia|9820/3
C0023448|T191|SY|C7539|NCI_CDISC|Lymphogenous Leukemia|9820/3
C0023448|T191|PT|C7539|NCI_CPTAC|Lymphoid Leukemia|9820/3
C0023448|T191|PT|C7539|NCI_CTRP|Lymphoid Leukemia|9820/3
C0023448|T191|DN|C7539|NCI_CTRP|Lymphoid Leukemia|9820/3
C0023448|T191|PT|CDR0000330173|NCI_NCI-GLOSS|lymphocytic leukemia|9820/3
C0023448|T191|SY|B64..|RCD|Lymphatic leukaemia|9820/3
C0023448|T191|PT|B64..|RCD|Lymphoid leukaemia|9820/3
C0023448|T191|OP|B64z.|RCD|Lymphoid leukaemia NOS|9820/3
C0023448|T191|SY|B64..|RCDAE|Lymphatic leukemia|9820/3
C0023448|T191|PT|B64..|RCDAE|Lymphoid leukemia|9820/3
C0023448|T191|OP|B64z.|RCDAE|Lymphoid leukemia NOS|9820/3
C0023448|T191|OP|BBr20|RCDSA|Lymphoid leukemia NOS|9820/3
C0023448|T191|PT|BBr2.|RCDSA|Lymphoid leukemias|9820/3
C0023448|T191|OP|BBr20|RCDSY|Lymphoid leukaemia NOS|9820/3
C0023448|T191|PT|BBr2.|RCDSY|Lymphoid leukaemias|9820/3
C0023448|T191|SYGB|188725004|SNOMEDCT_US|Lymphatic leukaemia|9820/3
C0023448|T191|SYGB|32280000|SNOMEDCT_US|Lymphatic leukaemia|9820/3
C0023448|T191|SY|32280000|SNOMEDCT_US|Lymphatic leukemia|9820/3
C0023448|T191|SY|188725004|SNOMEDCT_US|Lymphatic leukemia|9820/3
C0023448|T191|IS|32280000|SNOMEDCT_US|Lymphatic leukemia, NOS|9820/3
C0023448|T191|SYGB|32280000|SNOMEDCT_US|Lymphocytic leukaemia|9820/3
C0023448|T191|SY|32280000|SNOMEDCT_US|Lymphocytic leukemia|9820/3
C0023448|T191|IS|32280000|SNOMEDCT_US|Lymphocytic leukemia, NOS|9820/3
C0023448|T191|PTGB|32280000|SNOMEDCT_US|Lymphoid leukaemia|9820/3
C0023448|T191|PTGB|188725004|SNOMEDCT_US|Lymphoid leukaemia|9820/3
C0023448|T191|OAP|93170002|SNOMEDCT_US|Lymphoid leukaemia|9820/3
C0023448|T191|OAS|269631008|SNOMEDCT_US|Lymphoid leukaemia|9820/3
C0023448|T191|OAS|154587007|SNOMEDCT_US|Lymphoid leukaemia|9820/3
C1292765|T185|SYGB|128935007|SNOMEDCT_US|Lymphoid leukaemia - category|9820/3
C0023448|T191|OAP|188731001|SNOMEDCT_US|Lymphoid leukaemia NOS|9820/3
C0023448|T191|SYGB|32280000|SNOMEDCT_US|Lymphoid leukaemia, no ICD-O subtype|9820/3
C0023448|T191|PT|32280000|SNOMEDCT_US|Lymphoid leukemia|9820/3
C0023448|T191|OAP|93170002|SNOMEDCT_US|Lymphoid leukemia|9820/3
C0023448|T191|OAS|154587007|SNOMEDCT_US|Lymphoid leukemia|9820/3
C0023448|T191|OAS|269631008|SNOMEDCT_US|Lymphoid leukemia|9820/3
C0023448|T191|PT|188725004|SNOMEDCT_US|Lymphoid leukemia|9820/3
C1292765|T185|SY|128935007|SNOMEDCT_US|Lymphoid leukemia - category|9820/3
C0023448|T191|OAP|188731001|SNOMEDCT_US|Lymphoid leukemia NOS|9820/3
C0023448|T191|SY|32280000|SNOMEDCT_US|Lymphoid leukemia, no ICD-O subtype|9820/3
C0023448|T191|SY|32280000|SNOMEDCT_US|Lymphoid leukemia, no International Classification of Diseases for Oncology subtype|9820/3
C0023448|T191|IS|32280000|SNOMEDCT_US|Lymphoid leukemia, NOS|9820/3
C0023448|T191|IT|0176|WHO|LEUKAEMIA LYMPHATIC|9820/3
C0023448|T191|PT|0176|WHO|LEUKAEMIA LYMPHOCYTIC|9820/3
C0023448|T191|IT|0176|WHO|LEUKAEMIA LYMPHOID|9820/3
C0023434|T191|PT|BI00303|BI|chronic lymphocytic leukemia|9823/3
C0023434|T191|AB|BI00303|BI|cll|9823/3
C0023434|T191|PT|0052930|CCPSS|LEUKEMIA CHRONIC LYMPHOCYTIC|9823/3
C0023434|T191|SY|0000007331|CHV|b cell leukemia|9823/3
C0023434|T191|SY|0000007331|CHV|b cell lymphocytic leukemia|9823/3
C0023434|T191|SY|0000007333|CHV|b chronic lymphocytic leukemia|9823/3
C0023434|T191|PT|0000007333|CHV|b-cell cll|9823/3
C0023434|T191|PT|0000007331|CHV|b-cell leukemia|9823/3
C0023434|T191|SY|0000007339|CHV|chronic leukemia lymphocytic|9823/3
C0023434|T191|SY|0000007339|CHV|chronic lymphatic leukaemia|9823/3
C0023434|T191|SY|0000007339|CHV|chronic lymphatic leukemia|9823/3
C0023434|T191|SY|0000007339|CHV|chronic lymphoblastic leukemia|9823/3
C0023434|T191|SY|0000007339|CHV|chronic lymphocytic leukaemia|9823/3
C0023434|T191|SY|0000007339|CHV|chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|0000007339|CHV|chronic lymphogenous leukemia|9823/3
C0023434|T191|SY|0000007339|CHV|chronic lymphoid leukemia|9823/3
C0023434|T191|SY|0000007339|CHV|cll|9823/3
C0023434|T191|SY|0000007339|CHV|cll chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|0000007339|CHV|clls|9823/3
C0023434|T191|SY|0000007331|CHV|leukemia b cell|9823/3
C0023434|T191|SY|0000007339|CHV|leukemia chronic lymphocytic|9823/3
C0023434|T191|SY|0000007339|CHV|lymphocytic leukemia chronic|9823/3
C0023434|T191|PT|183|COSTAR|CHRONIC LYMPHOCYTIC LEUKEMIA|9823/3
C0023434|T191|ET|4005-0012|CSP|chronic lymphatic leukemia|9823/3
C0023434|T191|PT|4005-0012|CSP|chronic lymphocytic leukemia|9823/3
C0023434|T191|ET|4005-0012|CSP|chronic lymphogenous leukemia|9823/3
C0023434|T191|ET|4005-0012|CSP|chronic lymphoid leukemia|9823/3
C0023434|T191|ET|4005-0012|CSP|CLL|9823/3
C0023434|T191|PT|LEUKEMIA CHRON LYMPHO|CST|CHRONIC LYMPHOCYTIC LEUKEMIA|9823/3
C0023434|T191|GT|LEUKEMIA CHRON LYMPHO|CST|LEUKEMIA LYMPHOCYTIC CHRONIC|9823/3
C0023434|T191|SY|NOCODE|DXP|CLL|9823/3
C0023434|T191|DI|U001048|DXP|LEUKEMIA, LYMPHOCYTIC, CHRONIC|9823/3
C0023434|T191|PT|HP:0005550|HPO|Chronic lymphatic leukemia|9823/3
C0023434|T191|SY|HP:0005550|HPO|Chronic lymphocytic leukemia|9823/3
C0023434|T191|PT|C91.1|ICD10|Chronic lymphocytic leukaemia|9823/3
C0023434|T191|PT|C91.1|ICD10AE|Chronic lymphocytic leukemia|9823/3
C0023434|T191|AB|C91.1|ICD10CM|Chronic lymphocytic leukemia of B-cell type|9823/3
C0023434|T191|HT|C91.1|ICD10CM|Chronic lymphocytic leukemia of B-cell type|9823/3
C0023434|T191|ET|C91.10|ICD10CM|Chronic lymphocytic leukemia of B-cell type NOS|9823/3
C0023434|T191|HT|204.1|ICD9CM|Lymphoid leukemia, chronic|9823/3
C0023434|T191|PT|MTHU044764|ICPC2ICD10ENG|leukemia; lymphatic, chronic|9823/3
C0023434|T191|PT|MTHU046614|ICPC2ICD10ENG|lymphatic; leukemia, chronic|9823/3
C0023434|T191|PTN|B73004|ICPC2P|chronic lymphocytic leukaemia|9823/3
C0023434|T191|MTH_PTN|B73004|ICPC2P|chronic lymphocytic leukemia|9823/3
C0023434|T191|PT|B73004|ICPC2P|Leukaemia;chronic lymphocytic|9823/3
C0023434|T191|MTH_PT|B73004|ICPC2P|Leukemia;chronic lymphocytic|9823/3
C0023434|T191|PT|sh87004460|LCH_NW|Chronic lymphocytic leukemia|9823/3
C0023434|T191|LPN|LP208602-5|LNC|Chronic lymphocytic leukemia|9823/3
C1302547|T191|LA|LA26790-8|LNC|Chronic lymphocytic leukemia/small lymphocytic lymphoma|9823/3
C0023434|T191|LPN|LP34550-1|LNC|CLL|9823/3
C0023434|T191|LLT|10008956|MDR|Chronic lymphatic leukaemia|9823/3
C0023434|T191|LLT|10008957|MDR|Chronic lymphatic leukemia|9823/3
C0023434|T191|PT|10008958|MDR|Chronic lymphocytic leukaemia|9823/3
C0023434|T191|LLT|10008958|MDR|Chronic lymphocytic leukaemia|9823/3
C0023434|T191|LLT|10008960|MDR|Chronic lymphocytic leukaemia NOS|9823/3
C0023434|T191|LLT|10008976|MDR|Chronic lymphocytic leukemia|9823/3
C0023434|T191|MTH_PT|10008958|MDR|Chronic lymphocytic leukemia|9823/3
C0023434|T191|MTH_LLT|10008960|MDR|Chronic lymphocytic leukemia NOS|9823/3
C0023434|T191|LLT|10008993|MDR|Chronic lymphoid leukaemia|9823/3
C0023434|T191|LLT|10060576|MDR|Chronic lymphoid leukemia|9823/3
C0023434|T191|LLT|10009310|MDR|CLL|9823/3
C0023434|T191|LLT|10060391|MDR|Leukaemia lymphocytic chronic|9823/3
C0023434|T191|HT|10024295|MDR|Leukaemias chronic lymphocytic|9823/3
C0023434|T191|LLT|10024340|MDR|Leukemia lymphocytic chronic|9823/3
C0023434|T191|MTH_HT|10024295|MDR|Leukemias chronic lymphocytic|9823/3
C0023434|T191|LLT|10025302|MDR|Lymphoid leukaemia, chronic|9823/3
C0023434|T191|LLT|10025306|MDR|Lymphoid leukemia, chronic|9823/3
C0023434|T191|SY|230905|MEDCIN|B-cell chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|230905|MEDCIN|B-cell CLL|9823/3
C0023434|T191|PT|230905|MEDCIN|chronic B-cell lymphocytic leukemia|9823/3
C0023434|T191|PT|31473|MEDCIN|chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|31473|MEDCIN|CLL|9823/3
C0023434|T191|PT|87|MEDLINEPLUS|Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|ET|87|MEDLINEPLUS|CLL|9823/3
C0023434|T191|SY|87|MEDLINEPLUS|CLL|9823/3
C0023434|T191|ET|87|MEDLINEPLUS|Leukemia, Chronic Lymphocytic|9823/3
C0023434|T191|PM|D015451|MSH|B Cell Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|PM|D015451|MSH|B Cell Leukemia, Chronic|9823/3
C0023434|T191|PM|D015451|MSH|B Lymphocytic Leukemia, Chronic|9823/3
C0023434|T191|ET|D015451|MSH|B-Cell Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|ET|D015451|MSH|B-Cell Leukemia, Chronic|9823/3
C0023434|T191|PM|D015451|MSH|B-Cell Leukemias, Chronic|9823/3
C0023434|T191|ET|D015451|MSH|B-Cell Malignancy, Low-Grade|9823/3
C0023434|T191|ET|D015451|MSH|B-Lymphocytic Leukemia, Chronic|9823/3
C0023434|T191|PM|D015451|MSH|B-Lymphocytic Leukemias, Chronic|9823/3
C0023434|T191|PM|D015451|MSH|Chronic B-Cell Leukemia|9823/3
C0023434|T191|PM|D015451|MSH|Chronic B-Cell Leukemias|9823/3
C0023434|T191|PM|D015451|MSH|Chronic B-Lymphocytic Leukemia|9823/3
C0023434|T191|PM|D015451|MSH|Chronic B-Lymphocytic Leukemias|9823/3
C0023434|T191|PM|D015451|MSH|Chronic Lymphoblastic Leukemia|9823/3
C0023434|T191|PM|D015451|MSH|Chronic Lymphoblastic Leukemias|9823/3
C0023434|T191|ET|D015451|MSH|Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|PM|D015451|MSH|Chronic Lymphocytic Leukemias|9823/3
C0023434|T191|PM|D015451|MSH|CLL Lymphoplasmacytoid Lymphoma|9823/3
C0023434|T191|PM|D015451|MSH|CLL Lymphoplasmacytoid Lymphomas|9823/3
C0023434|T191|DEV|D015451|MSH|DIFFUSE WELL DIFFER LYMPHOCYTIC LYMPHOMA|9823/3
C0023434|T191|PM|D015451|MSH|Diffuse Well Differentiated Lymphocytic Lymphoma|9823/3
C0023434|T191|ET|D015451|MSH|Diffuse Well-Differentiated Lymphocytic Lymphoma|9823/3
C0023434|T191|ET|D015451|MSH|Disrupted In B-Cell Malignancy|9823/3
C0023434|T191|ET|D015451|MSH|Leukemia, B Cell, Chronic|9823/3
C0023434|T191|ET|D015451|MSH|Leukemia, B-Cell, Chronic|9823/3
C0023434|T191|PM|D015451|MSH|Leukemia, Chronic B-Cell|9823/3
C0023434|T191|PM|D015451|MSH|Leukemia, Chronic B-Lymphocytic|9823/3
C0023434|T191|ET|D015451|MSH|Leukemia, Chronic Lymphatic|9823/3
C0023434|T191|ET|D015451|MSH|Leukemia, Chronic Lymphocytic|9823/3
C0023434|T191|ET|D015451|MSH|Leukemia, Chronic Lymphocytic, B-Cell|9823/3
C0023434|T191|ET|D015451|MSH|Leukemia, Lymphoblastic, Chronic|9823/3
C0023434|T191|ET|D015451|MSH|Leukemia, Lymphocytic, Chronic|9823/3
C0023434|T191|ET|D015451|MSH|Leukemia, Lymphocytic, Chronic, B Cell|9823/3
C0023434|T191|MH|D015451|MSH|Leukemia, Lymphocytic, Chronic, B-Cell|9823/3
C0023434|T191|PM|D015451|MSH|Leukemias, Chronic B-Cell|9823/3
C0023434|T191|PM|D015451|MSH|Leukemias, Chronic B-Lymphocytic|9823/3
C0023434|T191|PM|D015451|MSH|Leukemias, Chronic Lymphoblastic|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoblastic Leukemia, Chronic|9823/3
C0023434|T191|PM|D015451|MSH|Lymphoblastic Leukemias, Chronic|9823/3
C0023434|T191|DSV|D015451|MSH|LYMPHOCYTIC LEUKEMIA CHRONIC B|9823/3
C0023434|T191|ET|D015451|MSH|Lymphocytic Leukemia, Chronic|9823/3
C0023434|T191|ET|D015451|MSH|Lymphocytic Leukemia, Chronic, B Cell|9823/3
C0023434|T191|ET|D015451|MSH|Lymphocytic Leukemia, Chronic, B-Cell|9823/3
C0023434|T191|PM|D015451|MSH|Lymphocytic Leukemias, Chronic|9823/3
C0023434|T191|ET|D015451|MSH|Lymphocytic Lymphoma|9823/3
C0023434|T191|DEV|D015451|MSH|LYMPHOCYTIC LYMPHOMA DIFFUSE WELL DIFFER|9823/3
C0023434|T191|DEV|D015451|MSH|LYMPHOCYTIC LYMPHOMA WELL DIFFER|9823/3
C0023434|T191|ET|D015451|MSH|Lymphocytic Lymphoma, Diffuse, Well Differentiated|9823/3
C0023434|T191|ET|D015451|MSH|Lymphocytic Lymphoma, Diffuse, Well-Differentiated|9823/3
C0023434|T191|PM|D015451|MSH|Lymphocytic Lymphoma, Small|9823/3
C0023434|T191|ET|D015451|MSH|Lymphocytic Lymphoma, Well Differentiated|9823/3
C0023434|T191|ET|D015451|MSH|Lymphocytic Lymphoma, Well-Differentiated|9823/3
C0023434|T191|PM|D015451|MSH|Lymphocytic Lymphomas|9823/3
C0023434|T191|PM|D015451|MSH|Lymphocytic Lymphomas, Small|9823/3
C0023434|T191|PM|D015451|MSH|Lymphocytic Lymphomas, Well-Differentiated|9823/3
C0023434|T191|DEV|D015451|MSH|LYMPHOMA LYMPHOCYTIC DIFFUSE WELL DIFFER|9823/3
C0023434|T191|DEV|D015451|MSH|LYMPHOMA LYMPHOCYTIC WELL DIFFER|9823/3
C0023434|T191|DEV|D015451|MSH|LYMPHOMA SMALL|9823/3
C0023434|T191|PM|D015451|MSH|Lymphoma, CLL Lymphoplasmacytoid|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Lymphocytic|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Lymphocytic, Diffuse, Well Differentiated|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Lymphocytic, Diffuse, Well-Differentiated|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Lymphocytic, Well Differentiated|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Lymphocytic, Well-Differentiated|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Lymphoplasmacytoid, CLL|9823/3
C0023434|T191|PM|D015451|MSH|Lymphoma, Small Cell|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Small Lymphocytic|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Small Lymphocytic, Plasmacytoid|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoma, Small-Cell|9823/3
C0023434|T191|PM|D015451|MSH|Lymphoma, Well-Differentiated Lymphocytic|9823/3
C0023434|T191|PM|D015451|MSH|Lymphomas, CLL Lymphoplasmacytoid|9823/3
C0023434|T191|PM|D015451|MSH|Lymphomas, Lymphocytic|9823/3
C0023434|T191|PM|D015451|MSH|Lymphomas, Small Lymphocytic|9823/3
C0023434|T191|PM|D015451|MSH|Lymphomas, Small-Cell|9823/3
C0023434|T191|PM|D015451|MSH|Lymphomas, Well-Differentiated Lymphocytic|9823/3
C0023434|T191|ET|D015451|MSH|Lymphoplasmacytoid Lymphoma, CLL|9823/3
C0023434|T191|PM|D015451|MSH|Lymphoplasmacytoid Lymphomas, CLL|9823/3
C0023434|T191|PM|D015451|MSH|Small Cell Lymphoma|9823/3
C0023434|T191|PM|D015451|MSH|Small Lymphocytic Lymphoma|9823/3
C0023434|T191|PM|D015451|MSH|Small Lymphocytic Lymphomas|9823/3
C0023434|T191|DEV|D015451|MSH|SMALL LYMPHOMA|9823/3
C0023434|T191|ET|D015451|MSH|Small-Cell Lymphoma|9823/3
C0023434|T191|PM|D015451|MSH|Small-Cell Lymphomas|9823/3
C0023434|T191|PM|D015451|MSH|Well-Differentiated Lymphocytic Lymphoma|9823/3
C0023434|T191|PM|D015451|MSH|Well-Differentiated Lymphocytic Lymphomas|9823/3
C0023434|T191|PN|NOCODE|MTH|Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|SY|C3163|NCI|B Cell Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|SY|C3163|NCI|B Cell CLL|9823/3
C0023434|T191|SY|C3163|NCI|B Cell Lymphocytic Leukemia|9823/3
C0023434|T191|SY|C3163|NCI|B-Cell Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|SY|C3163|NCI|B-Cell Chronic Lymphogenous Leukemia|9823/3
C0023434|T191|SY|C3163|NCI|B-Cell Chronic Lymphoid Leukemia|9823/3
C0023434|T191|SY|C3163|NCI|B-Cell CLL|9823/3
C0023434|T191|SY|C3163|NCI|B-Cell Lymphocytic Leukemia|9823/3
C0023434|T191|AB|C3163|NCI|BCLL|9823/3
C0023434|T191|SY|C3163|NCI|Chronic B-Cell Lymphocytic Leukemia|9823/3
C0023434|T191|SY|C3163|NCI|Chronic Lymphatic Leukemia|9823/3
C0023434|T191|PT|C3163|NCI|Chronic Lymphocytic Leukemia|9823/3
C1302547|T191|PT|C27911|NCI|Chronic Lymphocytic Leukemia/Small Lymphocytic Lymphoma|9823/3
C1302547|T191|SY|TCGA|NCI|Chronic Lymphocytic Leukemia/Small Lymphocytic Lymphoma|9823/3
C0023434|T191|SY|C3163|NCI|Chronic Lymphogenous Leukemia|9823/3
C0023434|T191|AB|C3163|NCI|CLL|9823/3
C1302547|T191|AB|C27911|NCI|CLL/SLL|9823/3
C0023434|T191|PT|C3163|NCI_CPTAC|Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|PT|10008960|NCI_CTEP-SDC|Chronic lymphocytic leukemia, NOS|9823/3
C0023434|T191|SY|C3163|NCI_CTRP|Chronic Lymphocytic Leukemia|9823/3
C0023434|T191|PT|CDR0000044846|NCI_NCI-GLOSS|chronic lymphocytic leukemia|9823/3
C1302547|T191|PT|CDR0000641290|NCI_NCI-GLOSS|chronic lymphocytic leukemia/small lymphocytic lymphoma|9823/3
C0023434|T191|PT|CDR0000346545|NCI_NCI-GLOSS|CLL|9823/3
C1302547|T191|PT|CDR0000641291|NCI_NCI-GLOSS|CLL/SLL|9823/3
C0023434|T191|SY|CDR0000039824|PDQ|B cell chronic lymphocytic leukemia|9823/3
C0023434|T191|PT|CDR0000039824|PDQ|B-cell chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|CDR0000039824|PDQ|B-cell CLL|9823/3
C0023434|T191|PT|CDR0000037765|PDQ|chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|CDR0000039824|PDQ|chronic lymphocytic leukemia, B-cell|9823/3
C0023434|T191|AB|CDR0000037765|PDQ|CLL|9823/3
C0023434|T191|SY|CDR0000039824|PDQ|CLL, B-cell|9823/3
C0023434|T191|SY|CDR0000039824|PDQ|leukemia, B-cell chronic lymphocytic|9823/3
C0023434|T191|SY|CDR0000037765|PDQ|leukemia, chronic lymphocytic|9823/3
C0023434|T191|SY|CDR0000039824|PDQ|lymphocytic leukemia, B-cell chronic|9823/3
C0023434|T191|SY|CDR0000037765|PDQ|lymphocytic leukemia, chronic|9823/3
C0023434|T191|PT|R0121662|QMR|LEUKEMIA CHRONIC LYMPHOCYTIC|9823/3
C0023434|T191|AB|Xa0QP|RCD|B-cell chron lymphocyt leukaem|9823/3
C0023434|T191|PT|Xa0QP|RCD|B-cell chronic lymphocytic leukaemia|9823/3
C0023434|T191|AB|Xa0QP|RCD|B-CLL - B-cell chron lymp leuk|9823/3
C0023434|T191|SY|Xa0QP|RCD|B-CLL - B-cell chronic lymphocytic leukaemia|9823/3
C0023434|T191|SY|B641.|RCD|Chronic lymphatic leukaemia|9823/3
C0023434|T191|SY|B641.|RCD|Chronic lymphocytic leukaemia|9823/3
C0023434|T191|PT|B641.|RCD|Chronic lymphoid leukaemia|9823/3
C0023434|T191|SY|B641.|RCD|CLL - Chronic lymphocytic leukaemia|9823/3
C0023434|T191|AB|B641.|RCD|CLL-Chron lymphocyt leukaemia|9823/3
C0023434|T191|PT|Xa0QP|RCDAE|B-cell chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|Xa0QP|RCDAE|B-CLL - B-cell chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|B641.|RCDAE|Chronic lymphatic leukemia|9823/3
C0023434|T191|SY|B641.|RCDAE|Chronic lymphocytic leukemia|9823/3
C0023434|T191|PT|B641.|RCDAE|Chronic lymphoid leukemia|9823/3
C0023434|T191|SY|B641.|RCDAE|CLL - Chronic lymphocytic leukemia|9823/3
C0023434|T191|AB|B641.|RCDAE|CLL-Chron lymphocyt leukemia|9823/3
C0023434|T191|PT|BBr23|RCDSA|Chronic lymphoid leukemia|9823/3
C0023434|T191|PT|BBr23|RCDSY|Chronic lymphoid leukaemia|9823/3
C0023434|T191|PTGB|277473004|SNOMEDCT_US|B-cell chronic lymphocytic leukaemia|9823/3
C0023434|T191|SYGB|51092000|SNOMEDCT_US|B-cell chronic lymphocytic leukaemia/small lymphocytic lymphoma|9823/3
C0023434|T191|PT|277473004|SNOMEDCT_US|B-cell chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|51092000|SNOMEDCT_US|B-cell chronic lymphocytic leukemia/small lymphocytic lymphoma|9823/3
C0023434|T191|SYGB|277473004|SNOMEDCT_US|B-CLL - B-cell chronic lymphocytic leukaemia|9823/3
C0023434|T191|SY|277473004|SNOMEDCT_US|B-CLL - B-cell chronic lymphocytic leukemia|9823/3
C0023434|T191|SYGB|51092000|SNOMEDCT_US|Chronic lymphatic leukaemia|9823/3
C0023434|T191|SY|51092000|SNOMEDCT_US|Chronic lymphatic leukemia|9823/3
C0023434|T191|PTGB|51092000|SNOMEDCT_US|Chronic lymphocytic leukaemia|9823/3
C0023434|T191|SYGB|51092000|SNOMEDCT_US|Chronic lymphocytic leukaemia, B-cell type|9823/3
C1302547|T191|OAP|399607007|SNOMEDCT_US|Chronic lymphocytic leukaemia/small lymphocytic lymphoma|9823/3
C0023434|T191|PT|51092000|SNOMEDCT_US|Chronic lymphocytic leukemia|9823/3
C0023434|T191|SY|51092000|SNOMEDCT_US|Chronic lymphocytic leukemia, B-cell type|9823/3
C1302547|T191|OAP|399607007|SNOMEDCT_US|Chronic lymphocytic leukemia/small lymphocytic lymphoma|9823/3
C0023434|T191|SYGB|92814006|SNOMEDCT_US|Chronic lymphoid leukaemia|9823/3
C0023434|T191|SYGB|51092000|SNOMEDCT_US|Chronic lymphoid leukaemia|9823/3
C1531666|T191|PTGB|413840004|SNOMEDCT_US|Chronic lymphoid leukaemia - category|9823/3
C0023434|T191|PTGB|92814006|SNOMEDCT_US|Chronic lymphoid leukaemia, disease|9823/3
C0023434|T191|SY|92814006|SNOMEDCT_US|Chronic lymphoid leukemia|9823/3
C0023434|T191|SY|51092000|SNOMEDCT_US|Chronic lymphoid leukemia|9823/3
C1531666|T191|PT|413840004|SNOMEDCT_US|Chronic lymphoid leukemia - category|9823/3
C0023434|T191|PT|92814006|SNOMEDCT_US|Chronic lymphoid leukemia, disease|9823/3
C0023434|T191|SYGB|92814006|SNOMEDCT_US|CLL - Chronic lymphocytic leukaemia|9823/3
C0023434|T191|SY|92814006|SNOMEDCT_US|CLL - Chronic lymphocytic leukemia|9823/3
C4721444|T191|SY|0000007332|CHV|b all|9826/3
C4721444|T191|SY|0000007332|CHV|b-all|9826/3
C4721444|T191|SY|0000007332|CHV|burkitt leukemia|9826/3
C4721444|T191|SY|0000007332|CHV|burkitt's leukemia|9826/3
C4721444|T191|PT|0000007332|CHV|burkitts leukemia|9826/3
C4721444|T191|PT|MTHU013215|ICPC2ICD10ENG|Burkitt; cell leukemia|9826/3
C4721444|T191|PT|MTHU015333|ICPC2ICD10ENG|cell leukemia; Burkitt|9826/3
C4721444|T191|LLT|10067184|MDR|Burkitt's leukaemia|9826/3
C4721444|T191|PT|10067184|MDR|Burkitt's leukaemia|9826/3
C4721444|T191|LLT|10067194|MDR|Burkitt's leukemia|9826/3
C4721444|T191|MTH_PT|10067184|MDR|Burkitt's leukemia|9826/3
C4721444|T191|PT|230906|MEDCIN|Burkitt cell leukemia|9826/3
C4721444|T191|SY|230906|MEDCIN|leukemia Burkitt cell|9826/3
C4721444|T191|ET|D002051|MSH|Burkitt Cell Leukemia|9826/3
C4721444|T191|PEP|D002051|MSH|Burkitt Leukemia|9826/3
C4721444|T191|ET|D002051|MSH|Burkitt's Leukemia|9826/3
C4721444|T191|PM|D002051|MSH|Burkitts Leukemia|9826/3
C4721444|T191|PM|D002051|MSH|L3 Lymphocytic Leukemia|9826/3
C4721444|T191|PM|D002051|MSH|L3 Lymphocytic Leukemias|9826/3
C4721444|T191|PM|D002051|MSH|Leukemia, Burkitt|9826/3
C4721444|T191|PM|D002051|MSH|Leukemia, Burkitt Cell|9826/3
C4721444|T191|PM|D002051|MSH|Leukemia, Burkitt's|9826/3
C4721444|T191|PM|D002051|MSH|Leukemia, L3 Lymphocytic|9826/3
C4721444|T191|ET|D002051|MSH|Leukemia, Lymphoblastic, Burkitt-Type|9826/3
C4721444|T191|ET|D002051|MSH|Leukemia, Lymphocytic, L3|9826/3
C4721444|T191|ET|D002051|MSH|Lymphocytic Leukemia, L3|9826/3
C4721444|T191|PN|NOCODE|MTH|Burkitt Leukemia|9826/3
C4721444|T191|PT|C7400|NCI|Burkitt Leukemia|9826/3
C4721444|T191|SY|TCGA|NCI|Burkitt Leukemia|9826/3
C4721444|T191|SY|C7400|NCI|Burkitt's Cell Leukemia|9826/3
C4721444|T191|SY|C7400|NCI|Burkitt's Leukemia|9826/3
C4721444|T191|OP|C7400|NCI|FAB L3|9826/3
C4721444|T191|OP|C7400|NCI|L3 Acute Lymphoblastic Leukemia|9826/3
C4721444|T191|OP|C7400|NCI|L3 Acute Lymphocytic Leukemia|9826/3
C4721444|T191|OP|C7400|NCI|L3 Acute Lymphogenous Leukemia|9826/3
C4721444|T191|OP|C7400|NCI|L3 Acute Lymphoid Leukemia|9826/3
C4721444|T191|PT|C7400|NCI_CPTAC|Burkitt Leukemia|9826/3
C4721444|T191|PT|10006597|NCI_CTEP-SDC|Burkitt lymphoma/leukemia|9826/3
C4721444|T191|DN|C7400|NCI_CTRP|Burkitt Leukemia|9826/3
C4721444|T191|PT|CDR0000256548|NCI_NCI-GLOSS|Burkitt's leukemia|9826/3
C4721444|T191|OP|BBr26|RCD|Burkitt's cell leukaemia|9826/3
C4721444|T191|OP|BBr26|RCDAE|Burkitt's cell leukemia|9826/3
C4721444|T191|SYGB|22197008|SNOMEDCT_US|Acute lymphoblastic leukaemia, Burkitt's type|9826/3
C4721444|T191|SYGB|22197008|SNOMEDCT_US|Acute lymphoblastic leukaemia, mature B-cell type|9826/3
C4721444|T191|SY|22197008|SNOMEDCT_US|Acute lymphoblastic leukemia, Burkitt's type|9826/3
C4721444|T191|SY|22197008|SNOMEDCT_US|Acute lymphoblastic leukemia, mature B-cell type|9826/3
C4721444|T191|PTGB|277571004|SNOMEDCT_US|B-cell acute lymphoblastic leukaemia|9826/3
C4721444|T191|PTGB|22197008|SNOMEDCT_US|Burkitt cell leukaemia|9826/3
C4721444|T191|PT|22197008|SNOMEDCT_US|Burkitt cell leukemia|9826/3
C4721444|T191|SYGB|22197008|SNOMEDCT_US|Burkitt's cell leukaemia|9826/3
C4721444|T191|SY|22197008|SNOMEDCT_US|Burkitt's cell leukemia|9826/3
C4721444|T191|SYGB|277571004|SNOMEDCT_US|Burkitt's leukaemia|9826/3
C4721444|T191|SY|277571004|SNOMEDCT_US|Burkitt's leukemia|9826/3
C4721444|T191|IS|22197008|SNOMEDCT_US|FAB L3|9826/3
C0023493|T191|PT|0000007355|CHV|adult t-cell leukemia|9827/3
C0023493|T191|SY|0000007355|CHV|adult t-cell leukemias|9827/3
C0023493|T191|SY|0000007355|CHV|adult t-cell lymphoma|9827/3
C0023493|T191|SY|0000007355|CHV|atll|9827/3
C0023493|T191|SY|0000007355|CHV|human t cell leukemia|9827/3
C0023493|T191|SY|0000007354|CHV|t cell acute leukemia|9827/3
C0023493|T191|PT|0000007354|CHV|t-all|9827/3
C0023493|T191|ET|2004-1803|CSP|adult T cell leukemia|9827/3
C0023493|T191|PT|2004-1803|CSP|human T cell leukemia|9827/3
C0023493|T191|PT|C91.5|ICD10|Adult T-cell leukaemia|9827/3
C0023493|T191|PT|C91.5|ICD10AE|Adult T-cell leukemia|9827/3
C0023493|T191|PT|MTHU003786|ICPC2ICD10ENG|adult T-cell; leukemia|9827/3
C0023493|T191|PT|MTHU003787|ICPC2ICD10ENG|adult T-cell; lymphoma|9827/3
C0023493|T191|PT|MTHU044739|ICPC2ICD10ENG|leukemia; adult T-cell|9827/3
C0023493|T191|PT|MTHU046734|ICPC2ICD10ENG|lymphoma; adult T-cell|9827/3
C0023493|T191|PT|MTHU046857|ICPC2ICD10ENG|lymphoma; T-cell, adult|9827/3
C0023493|T191|PT|MTHU073540|ICPC2ICD10ENG|T-cell; lymphoma, adult|9827/3
C0023493|T191|PT|sh94002377|LCH_NW|Adult T-cell leukemia|9827/3
C0023493|T191|LLT|10001412|MDR|Adult T-cell leukemia-lymphoma|9827/3
C0023493|T191|LLT|10001413|MDR|Adult T-cell lymphoma/leukaemia|9827/3
C0023493|T191|PT|10001413|MDR|Adult T-cell lymphoma/leukaemia|9827/3
C0023493|T191|LLT|10001415|MDR|Adult T-cell lymphoma/leukaemia NOS|9827/3
C0023493|T191|LLT|10054298|MDR|Adult T-cell lymphoma/leukemia|9827/3
C0023493|T191|MTH_PT|10001413|MDR|Adult T-cell lymphoma/leukemia|9827/3
C0023493|T191|MTH_LLT|10001415|MDR|Adult T-cell lymphoma/leukemia NOS|9827/3
C0023493|T191|HT|10001414|MDR|Adult T-cell lymphomas/leukaemias|9827/3
C0023493|T191|MTH_HT|10001414|MDR|Adult T-cell lymphomas/leukemias|9827/3
C0023493|T191|OL|10003622|MDR|ATLL|9827/3
C0023493|T191|PT|31474|MEDCIN|adult T-cell leukemia|9827/3
C0023493|T191|PT|338557|MEDCIN|Adult T-cell leukemia/lymphoma|9827/3
C0023493|T191|SY|31474|MEDCIN|leukemia adult T-cell|9827/3
C0023493|T191|SY|338557|MEDCIN|leukemia/lymphoma adult t-cell|9827/3
C0023493|T191|PM|D015459|MSH|Adult T-Cell Leukemia|9827/3
C0023493|T191|PM|D015459|MSH|Adult T-Cell Leukemia-Lymphoma|9827/3
C0023493|T191|PM|D015459|MSH|Adult T-Cell Leukemia-Lymphomas|9827/3
C0023493|T191|PM|D015459|MSH|Adult T-Cell Leukemias|9827/3
C0023493|T191|ET|D015459|MSH|ATLL|9827/3
C0023493|T191|DEV|D015459|MSH|HTLV ALL|9827/3
C0023493|T191|PM|D015459|MSH|HTLV Associated Leukemia Lymphoma|9827/3
C0023493|T191|ET|D015459|MSH|HTLV I Associated T Cell Leukemia Lymphoma|9827/3
C0023493|T191|ET|D015459|MSH|HTLV-Associated Leukemia-Lymphoma|9827/3
C0023493|T191|PM|D015459|MSH|HTLV-Associated Leukemia-Lymphomas|9827/3
C0023493|T191|ET|D015459|MSH|HTLV-I-Associated T-Cell Leukemia-Lymphoma|9827/3
C0023493|T191|PM|D015459|MSH|HTLV-I-Associated T-Cell Leukemia-Lymphomas|9827/3
C0023493|T191|PM|D015459|MSH|Human T Cell Leukemia Lymphoma|9827/3
C0023493|T191|ET|D015459|MSH|Human T Lymphotropic Virus Associated Leukemia Lymphoma|9827/3
C0023493|T191|ET|D015459|MSH|Human T Lymphotropic Virus-Associated Leukemia-Lymphoma|9827/3
C0023493|T191|ET|D015459|MSH|Human T-Cell Leukemia-Lymphoma|9827/3
C0023493|T191|PM|D015459|MSH|Human T-Cell Leukemia-Lymphomas|9827/3
C0023493|T191|ET|D015459|MSH|Leukemia Lymphoma, Adult T Cell|9827/3
C0023493|T191|ET|D015459|MSH|Leukemia Lymphoma, T Cell, Acute, HTLV I Associated|9827/3
C0023493|T191|MH|D015459|MSH|Leukemia-Lymphoma, Adult T-Cell|9827/3
C0023493|T191|PM|D015459|MSH|Leukemia-Lymphoma, HTLV-Associated|9827/3
C0023493|T191|PM|D015459|MSH|Leukemia-Lymphoma, HTLV-I-Associated T-Cell|9827/3
C0023493|T191|PM|D015459|MSH|Leukemia-Lymphoma, Human T-Cell|9827/3
C0023493|T191|ET|D015459|MSH|Leukemia-Lymphoma, T-Cell, Acute, HTLV-I-Associated|9827/3
C0023493|T191|PM|D015459|MSH|Leukemia-Lymphomas, Adult T-Cell|9827/3
C0023493|T191|PM|D015459|MSH|Leukemia-Lymphomas, HTLV-Associated|9827/3
C0023493|T191|PM|D015459|MSH|Leukemia-Lymphomas, HTLV-I-Associated T-Cell|9827/3
C0023493|T191|PM|D015459|MSH|Leukemia-Lymphomas, Human T-Cell|9827/3
C0023493|T191|PM|D015459|MSH|Leukemia, Adult T Cell|9827/3
C0023493|T191|ET|D015459|MSH|Leukemia, Adult T-Cell|9827/3
C0023493|T191|PM|D015459|MSH|Leukemias, Adult T-Cell|9827/3
C0023493|T191|PM|D015459|MSH|T Cell Leukemia Lymphoma, Adult|9827/3
C0023493|T191|ET|D015459|MSH|T Cell Leukemia Lymphoma, HTLV I Associated|9827/3
C0023493|T191|ET|D015459|MSH|T Cell Leukemia, Adult|9827/3
C0023493|T191|ET|D015459|MSH|T-Cell Leukemia-Lymphoma, Adult|9827/3
C0023493|T191|ET|D015459|MSH|T-Cell Leukemia-Lymphoma, HTLV-I-Associated|9827/3
C0023493|T191|PM|D015459|MSH|T-Cell Leukemia-Lymphoma, Human|9827/3
C0023493|T191|PM|D015459|MSH|T-Cell Leukemia-Lymphomas, Adult|9827/3
C0023493|T191|PM|D015459|MSH|T-Cell Leukemia-Lymphomas, HTLV-I-Associated|9827/3
C0023493|T191|PM|D015459|MSH|T-Cell Leukemia-Lymphomas, Human|9827/3
C0023493|T191|ET|D015459|MSH|T-Cell Leukemia, Adult|9827/3
C0023493|T191|PM|D015459|MSH|T-Cell Leukemias, Adult|9827/3
C0023493|T191|PT|U000477|MTH|Adult T-cell leukemia|9827/3
C0023493|T191|PN|NOCODE|MTH|Adult T-Cell Lymphoma/Leukemia|9827/3
C0023493|T191|SY|C3184|NCI|Adult T Cell Lymphoma/Leukemia|9827/3
C0023493|T191|PT|C3184|NCI|Adult T-Cell Leukemia/Lymphoma|9827/3
C0023493|T191|SY|TCGA|NCI|Adult T-Cell Leukemia/Lymphoma|9827/3
C0023493|T191|SY|C3184|NCI|Adult T-Cell Lymphoma/Leukemia|9827/3
C0023493|T191|SY|C3184|NCI|ATLL|9827/3
C0023493|T191|SY|C3184|NCI|HTLV-1 Associated Adult T-Cell Lymphoma/Leukemia|9827/3
C0023493|T191|SY|C3184|NCI|HTLV-I Associated Adult T-Cell Leukemia/Lymphoma|9827/3
C0023493|T191|PT|10001415|NCI_CTEP-SDC|Adult T-cell leukemia/lymphoma|9827/3
C0023493|T191|DN|C3184|NCI_CTRP|Adult T-Cell Leukemia/Lymphoma|9827/3
C0023493|T191|PT|CDR0000269410|NCI_NCI-GLOSS|adult T-cell leukemia/lymphoma|9827/3
C0023493|T191|PT|CDR0000269411|NCI_NCI-GLOSS|ATLL|9827/3
C0023493|T191|SY|CDR0000040694|PDQ|Adult T Cell Lymphoma/Leukemia|9827/3
C0023493|T191|PT|CDR0000040694|PDQ|adult T-cell leukemia/lymphoma|9827/3
C0023493|T191|SY|CDR0000040694|PDQ|Adult T-Cell Lymphoma/Leukemia|9827/3
C0023493|T191|SY|CDR0000040694|PDQ|ATLL|9827/3
C0023493|T191|SY|CDR0000040694|PDQ|HTLV-1 Associated Adult T-Cell Lymphoma/Leukemia|9827/3
C0023493|T191|SY|CDR0000040694|PDQ|HTLV-I associated adult T-cell leukemia/lymphoma|9827/3
C0023493|T191|SY|CDR0000040694|PDQ|leukemia/lymphoma, adult T-cell|9827/3
C0023493|T191|ET|CDR0000040694|PDQ|T-cell leukemia/lymphoma, adult|9827/3
C0023493|T191|OP|B64y2|RCD|Adult T-cell leukaemia|9827/3
C0023493|T191|OP|B64y2|RCDAE|Adult T-cell leukemia|9827/3
C0023493|T191|OP|BBr27|RCDSA|Adult T-cell leukemia/lymphoma|9827/3
C0023493|T191|OA|BBr27|RCDSY|Adul T-cell leukem/lymphoma|9827/3
C0023493|T191|OP|BBr27|RCDSY|Adult T-cell leukaemia/lymphoma|9827/3
C0023493|T191|PTGB|188729005|SNOMEDCT_US|Adult T-cell leukaemia|9827/3
C0023493|T191|SYGB|77430005|SNOMEDCT_US|Adult T-cell leukaemia|9827/3
C0023493|T191|IS|110007008|SNOMEDCT_US|Adult T-cell leukaemia|9827/3
C0023493|T191|PTGB|110007008|SNOMEDCT_US|Adult T-cell leukaemia/lymphoma|9827/3
C0023493|T191|PTGB|77430005|SNOMEDCT_US|Adult T-cell leukaemia/lymphoma|9827/3
C0023493|T191|PT|188729005|SNOMEDCT_US|Adult T-cell leukemia|9827/3
C0023493|T191|IS|110007008|SNOMEDCT_US|Adult T-cell leukemia|9827/3
C0023493|T191|SY|77430005|SNOMEDCT_US|Adult T-cell leukemia|9827/3
C0023493|T191|PT|77430005|SNOMEDCT_US|Adult T-cell leukemia/lymphoma|9827/3
C0023493|T191|PT|110007008|SNOMEDCT_US|Adult T-cell leukemia/lymphoma|9827/3
C0023493|T191|SY|77430005|SNOMEDCT_US|Adult T-cell lymphoma|9827/3
C0023493|T191|SYGB|77430005|SNOMEDCT_US|Adult T-cell lymphoma/leukaemia|9827/3
C0023493|T191|SY|77430005|SNOMEDCT_US|Adult T-cell lymphoma/leukemia|9827/3
C1955861|T191|PT|MTHU046872|ICPC2ICD10ENG|lymphoproliferative; disease, T-gamma|9831/1
C1955861|T191|LLT|10065862|MDR|T-cell large granular lymphocytic leukemia|9831/1
C1955861|T191|SY|392217|MEDCIN|leukemia lymphocytic chronic T-cell large granular|9831/1
C1955861|T191|PT|392217|MEDCIN|T-cell large granular lymphocytic leukemia|9831/1
C1955861|T191|PM|D054066|MSH|Granular Lymphocytoses, Large|9831/1
C1955861|T191|PM|D054066|MSH|Granular Lymphocytosis, Large|9831/1
C1955861|T191|PM|D054066|MSH|Large Granular Lymphocytoses|9831/1
C1955861|T191|ET|D054066|MSH|Large Granular Lymphocytosis|9831/1
C1955861|T191|PM|D054066|MSH|Leukemia, T Cell Large Granular Lymphocytic|9831/1
C1955861|T191|PM|D054066|MSH|Leukemia, T LGL|9831/1
C1955861|T191|PEP|D054066|MSH|Leukemia, T-Cell Large Granular Lymphocytic|9831/1
C1955861|T191|ET|D054066|MSH|Leukemia, T-LGL|9831/1
C1955861|T191|PM|D054066|MSH|Leukemias, T-LGL|9831/1
C1955861|T191|PM|D054066|MSH|Lymphocytoses, Large Granular|9831/1
C1955861|T191|PM|D054066|MSH|Lymphocytosis, Large Granular|9831/1
C1955861|T191|PM|D054066|MSH|T Cell Large Granular Lymphocyte Leukemia|9831/1
C1955861|T191|PM|D054066|MSH|T Cell Large Granular Lymphocytic Leukemia|9831/1
C1955861|T191|PM|D054066|MSH|T LGL Leukemia|9831/1
C1955861|T191|ET|D054066|MSH|T-Cell Large Granular Lymphocyte Leukemia|9831/1
C1955861|T191|ET|D054066|MSH|T-Cell Large Granular Lymphocytic Leukemia|9831/1
C1955861|T191|ET|D054066|MSH|T-LGL Leukemia|9831/1
C1955861|T191|PM|D054066|MSH|T-LGL Leukemias|9831/1
C1955861|T191|PN|NOCODE|MTH|T-Cell Large Granular Lymphocyte Leukemia|9831/1
C1955861|T191|SY|C4664|NCI|Large Cell Granular Lymphogenous Leukemia|9831/1
C1955861|T191|SY|C4664|NCI|Large Cell Granular Lymphoid Leukemia|9831/1
C1955861|T191|SY|C4664|NCI|Large Granular Lymphocytic Leukemia|9831/1
C1955861|T191|SY|C4664|NCI|Large Granular Lymphocytosis|9831/1
C1955861|T191|AB|C4664|NCI|LGLL|9831/1
C1955861|T191|SY|C4664|NCI|T Gamma Lymphoproliferative Disorder|9831/1
C1955861|T191|SY|TCGA|NCI|T-Cell Large Granular Lymphocyte Leukemia|9831/1
C1955861|T191|PT|C4664|NCI|T-Cell Large Granular Lymphocyte Leukemia|9831/1
C1955861|T191|SY|C4664|NCI|T-Cell Large Granular Lymphocytic Leukemia|9831/1
C1955861|T191|SY|C4664|NCI|T-Gamma Lymphoproliferative Disorder|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|Large Cell Granular Lymphogenous Leukemia|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|Large Cell Granular Lymphoid Leukemia|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|Large Granular Lymphocytic Leukemia|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|Large Granular Lymphocytosis|9831/1
C1955861|T191|PT|C4664|NCI_CDISC|LEUKEMIA, LARGE GRANULAR LYMPHOCYTIC, MALIGNANT|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|LGLL|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|T Gamma Lymphoproliferative Disorder|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|T-Cell Large Granular Lymphocytic Leukemia|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|T-Gamma Lymphoproliferative Disorder|9831/1
C1955861|T191|SY|C4664|NCI_CDISC|Tgamma Large Granular Lymphocyte Leukemia|9831/1
C1955861|T191|SY|10065862|NCI_CTEP-SDC|T-cell large gran. lymph. leuk.|9831/1
C1955861|T191|PT|10065862|NCI_CTEP-SDC|T-cell large granular lymphocytic leukemia|9831/1
C1955861|T191|DN|C4664|NCI_CTRP|T-Cell Large Granular Lymphocyte Leukemia|9831/1
C1955861|T191|PT|CDR0000633892|NCI_NCI-GLOSS|T-cell large granular lymphocyte leukemia|9831/1
C1955861|T191|PT|CDR0000633893|NCI_NCI-GLOSS|T-LGL leukemia|9831/1
C1955861|T191|PT|CDR0000039823|PDQ|T-cell large granular lymphocyte leukemia|9831/1
C1955861|T191|OP|CDR0000040442|PDQ|T-gamma lymphoproliferative disorder|9831/1
C1955861|T191|SY|CDR0000039823|PDQ|T-gamma lymphoproliferative disorder|9831/1
C1955861|T191|OA|BBmC.|RCDSY|T-gam lymphoprolif disease|9831/1
C1955861|T191|OP|BBmC.|RCDSY|T-gamma lymphoproliferative disease|9831/1
C1955861|T191|PTGB|699818003|SNOMEDCT_US|T-cell large granular lymphocytic leukaemia|9831/1
C1955861|T191|PTGB|128819001|SNOMEDCT_US|T-cell large granular lymphocytic leukaemia|9831/1
C1955861|T191|PT|128819001|SNOMEDCT_US|T-cell large granular lymphocytic leukemia|9831/1
C1955861|T191|PT|699818003|SNOMEDCT_US|T-cell large granular lymphocytic leukemia|9831/1
C1955861|T191|SY|128819001|SNOMEDCT_US|T-cell large granular lymphocytosis|9831/1
C1955861|T191|PT|55081009|SNOMEDCT_US|T-gamma lymphoproliferative disease|9831/1
C1955861|T191|PT|MTHU046872|ICPC2ICD10ENG|lymphoproliferative; disease, T-gamma|9831/3
C1955861|T191|LLT|10065862|MDR|T-cell large granular lymphocytic leukemia|9831/3
C1512709|T191|PT|366687|MEDCIN|Chronic lymphoproliferative disorder of natural killer cells|9831/3
C1955861|T191|SY|392217|MEDCIN|leukemia lymphocytic chronic T-cell large granular|9831/3
C1512709|T191|SY|366687|MEDCIN|lymphoma mature nk/t-cell chronic lymphoproliferative of natural killer cells|9831/3
C1955861|T191|PT|392217|MEDCIN|T-cell large granular lymphocytic leukemia|9831/3
C1955861|T191|PM|D054066|MSH|Granular Lymphocytoses, Large|9831/3
C1955861|T191|PM|D054066|MSH|Granular Lymphocytosis, Large|9831/3
C1955861|T191|PM|D054066|MSH|Large Granular Lymphocytoses|9831/3
C1955861|T191|ET|D054066|MSH|Large Granular Lymphocytosis|9831/3
C1955861|T191|PM|D054066|MSH|Leukemia, T Cell Large Granular Lymphocytic|9831/3
C1955861|T191|PM|D054066|MSH|Leukemia, T LGL|9831/3
C1955861|T191|PEP|D054066|MSH|Leukemia, T-Cell Large Granular Lymphocytic|9831/3
C1955861|T191|ET|D054066|MSH|Leukemia, T-LGL|9831/3
C1955861|T191|PM|D054066|MSH|Leukemias, T-LGL|9831/3
C1955861|T191|PM|D054066|MSH|Lymphocytoses, Large Granular|9831/3
C1955861|T191|PM|D054066|MSH|Lymphocytosis, Large Granular|9831/3
C1955861|T191|PM|D054066|MSH|T Cell Large Granular Lymphocyte Leukemia|9831/3
C1955861|T191|PM|D054066|MSH|T Cell Large Granular Lymphocytic Leukemia|9831/3
C1955861|T191|PM|D054066|MSH|T LGL Leukemia|9831/3
C1955861|T191|ET|D054066|MSH|T-Cell Large Granular Lymphocyte Leukemia|9831/3
C1955861|T191|ET|D054066|MSH|T-Cell Large Granular Lymphocytic Leukemia|9831/3
C1955861|T191|ET|D054066|MSH|T-LGL Leukemia|9831/3
C1955861|T191|PM|D054066|MSH|T-LGL Leukemias|9831/3
C1512709|T191|PN|NOCODE|MTH|Chronic Lymphoproliferative Disorder of NK-Cells|9831/3
C1955861|T191|PN|NOCODE|MTH|T-Cell Large Granular Lymphocyte Leukemia|9831/3
C1512709|T191|PT|C39591|NCI|Chronic Lymphoproliferative Disorder of NK-Cells|9831/3
C1512709|T191|SY|C39591|NCI|Chronic NK-Cell Lymphocytosis|9831/3
C1512709|T191|SY|C39591|NCI|Chronic NK-Large Granular Lymphocyte Lymphoproliferative Disorder|9831/3
C1512709|T191|SY|C39591|NCI|Chronic NK-LGL Lymphoproliferative Disorder|9831/3
C1512709|T191|AB|C39591|NCI|CLPD-NK|9831/3
C1512709|T191|SY|C39591|NCI|Indolent Large Granular NK-Cell Lymphoproliferative Disorder|9831/3
C1512709|T191|SY|C39591|NCI|Indolent NK-Cell Lymphoproliferative Disorder|9831/3
C1955861|T191|SY|C4664|NCI|Large Cell Granular Lymphogenous Leukemia|9831/3
C1955861|T191|SY|C4664|NCI|Large Cell Granular Lymphoid Leukemia|9831/3
C1955861|T191|SY|C4664|NCI|Large Granular Lymphocytic Leukemia|9831/3
C1955861|T191|SY|C4664|NCI|Large Granular Lymphocytosis|9831/3
C1955861|T191|AB|C4664|NCI|LGLL|9831/3
C1512709|T191|SY|C39591|NCI|NK-Cell Large Granular Lymphocyte Lymphocytosis|9831/3
C1512709|T191|SY|C39591|NCI|NK-Type Lymphoproliferative Disorder of Granular Lymphocytes|9831/3
C1955861|T191|SY|C4664|NCI|T Gamma Lymphoproliferative Disorder|9831/3
C1955861|T191|PT|C4664|NCI|T-Cell Large Granular Lymphocyte Leukemia|9831/3
C1955861|T191|SY|TCGA|NCI|T-Cell Large Granular Lymphocyte Leukemia|9831/3
C1955861|T191|SY|C4664|NCI|T-Cell Large Granular Lymphocytic Leukemia|9831/3
C1955861|T191|SY|C4664|NCI|T-Gamma Lymphoproliferative Disorder|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|Large Cell Granular Lymphogenous Leukemia|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|Large Cell Granular Lymphoid Leukemia|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|Large Granular Lymphocytic Leukemia|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|Large Granular Lymphocytosis|9831/3
C1955861|T191|PT|C4664|NCI_CDISC|LEUKEMIA, LARGE GRANULAR LYMPHOCYTIC, MALIGNANT|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|LGLL|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|T Gamma Lymphoproliferative Disorder|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|T-Cell Large Granular Lymphocytic Leukemia|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|T-Gamma Lymphoproliferative Disorder|9831/3
C1955861|T191|SY|C4664|NCI_CDISC|Tgamma Large Granular Lymphocyte Leukemia|9831/3
C1955861|T191|SY|10065862|NCI_CTEP-SDC|T-cell large gran. lymph. leuk.|9831/3
C1955861|T191|PT|10065862|NCI_CTEP-SDC|T-cell large granular lymphocytic leukemia|9831/3
C1512709|T191|DN|C39591|NCI_CTRP|Chronic Lymphoproliferative Disorder of NK-Cells|9831/3
C1955861|T191|DN|C4664|NCI_CTRP|T-Cell Large Granular Lymphocyte Leukemia|9831/3
C1512709|T191|PT|CDR0000644322|NCI_NCI-GLOSS|natural killer-cell large granular lymphocyte leukemia|9831/3
C1512709|T191|PT|CDR0000659612|NCI_NCI-GLOSS|NK-LGL leukemia|9831/3
C1512709|T191|PT|CDR0000644323|NCI_NCI-GLOSS|NK-LGLL|9831/3
C1955861|T191|PT|CDR0000633892|NCI_NCI-GLOSS|T-cell large granular lymphocyte leukemia|9831/3
C1955861|T191|PT|CDR0000633893|NCI_NCI-GLOSS|T-LGL leukemia|9831/3
C1512709|T191|PT|CDR0000754723|PDQ|chronic lymphoproliferative disorder of NK cells|9831/3
C1512709|T191|LV|CDR0000754723|PDQ|Chronic Lymphoproliferative Disorder of NK-Cells|9831/3
C1512709|T191|SY|CDR0000754723|PDQ|chronic NK-cell lymphocytosis|9831/3
C1512709|T191|SY|CDR0000754723|PDQ|chronic NK-large granular lymphocyte lymphoproliferative disorder|9831/3
C1512709|T191|SY|CDR0000754723|PDQ|chronic NK-LGL lymphoproliferative disorder|9831/3
C1512709|T191|AB|CDR0000754723|PDQ|CLPD-NK|9831/3
C1512709|T191|SY|CDR0000754723|PDQ|indolent large granular NK-cell lymphoproliferative disorder|9831/3
C1512709|T191|SY|CDR0000754723|PDQ|indolent NK-cell lymphoproliferative disorder|9831/3
C1512709|T191|SY|CDR0000754723|PDQ|NK-cell large granular lymphocyte lymphocytosis|9831/3
C1955861|T191|PT|CDR0000039823|PDQ|T-cell large granular lymphocyte leukemia|9831/3
C1955861|T191|SY|CDR0000039823|PDQ|T-gamma lymphoproliferative disorder|9831/3
C1955861|T191|OP|CDR0000040442|PDQ|T-gamma lymphoproliferative disorder|9831/3
C1955861|T191|OA|BBmC.|RCDSY|T-gam lymphoprolif disease|9831/3
C1955861|T191|OP|BBmC.|RCDSY|T-gamma lymphoproliferative disease|9831/3
C1512709|T191|PT|722955006|SNOMEDCT_US|Chronic lymphoproliferative disorder of natural killer cells|9831/3
C1512709|T191|SY|722955006|SNOMEDCT_US|Chronic lymphoproliferative disorder of NK-cells|9831/3
C1955861|T191|PTGB|699818003|SNOMEDCT_US|T-cell large granular lymphocytic leukaemia|9831/3
C1955861|T191|PTGB|128819001|SNOMEDCT_US|T-cell large granular lymphocytic leukaemia|9831/3
C1955861|T191|PT|699818003|SNOMEDCT_US|T-cell large granular lymphocytic leukemia|9831/3
C1955861|T191|PT|128819001|SNOMEDCT_US|T-cell large granular lymphocytic leukemia|9831/3
C1955861|T191|SY|128819001|SNOMEDCT_US|T-cell large granular lymphocytosis|9831/3
C1955861|T191|PT|55081009|SNOMEDCT_US|T-gamma lymphoproliferative disease|9831/3
C0023486|T191|SY|0000007350|CHV|pll prolymphocytic leukemia|9832/3
C0023486|T191|SY|0000007350|CHV|pro-lymphocytic leukemia|9832/3
C0023486|T191|PT|0000007350|CHV|prolymphocytic leukemia|9832/3
C0023486|T191|PT|C91.3|ICD10|Prolymphocytic leukaemia|9832/3
C0023486|T191|PT|C91.3|ICD10AE|Prolymphocytic leukemia|9832/3
C0023486|T191|PT|MTHU044795|ICPC2ICD10ENG|leukemia; prolymphocytic|9832/3
C0023486|T191|PT|MTHU062033|ICPC2ICD10ENG|prolymphocytic; leukemia|9832/3
C0023486|T191|LLT|10036763|MDR|Pro-lymphocytic leukaemia|9832/3
C0023486|T191|LLT|10054582|MDR|Pro-lymphocytic leukemia|9832/3
C0023486|T191|LLT|10036888|MDR|Prolymphocytic leukaemia|9832/3
C0023486|T191|PT|10036888|MDR|Prolymphocytic leukaemia|9832/3
C0023486|T191|LLT|10036889|MDR|Prolymphocytic leukemia|9832/3
C0023486|T191|MTH_PT|10036888|MDR|Prolymphocytic leukemia|9832/3
C0023486|T191|SY|230907|MEDCIN|leukemia prolymphocytic|9832/3
C0023486|T191|PT|230907|MEDCIN|prolymphocytic leukemia|9832/3
C0023486|T191|MH|D015463|MSH|Leukemia, Prolymphocytic|9832/3
C0023486|T191|PM|D015463|MSH|Leukemias, Prolymphocytic|9832/3
C0023486|T191|ET|D015463|MSH|Prolymphocytic Leukemia|9832/3
C0023486|T191|PM|D015463|MSH|Prolymphocytic Leukemias|9832/3
C0023486|T191|PN|NOCODE|MTH|Prolymphocytic Leukemia|9832/3
C0023486|T191|PT|C3181|NCI|Prolymphocytic Leukemia|9832/3
C0023486|T191|DN|C3181|NCI_CTRP|Prolymphocytic Leukemia|9832/3
C0023486|T191|PT|CDR0000403143|NCI_NCI-GLOSS|PLL|9832/3
C0023486|T191|PT|CDR0000045380|NCI_NCI-GLOSS|prolymphocytic leukemia|9832/3
C0023486|T191|SY|CDR0000041618|PDQ|leukemia, prolymphocytic|9832/3
C0023486|T191|PT|CDR0000041618|PDQ|prolymphocytic leukemia|9832/3
C0023486|T191|ET|CDR0000041618|PDQ|Prolymphocytic leukemia|9832/3
C0023486|T191|SY|B64y1|RCD|PLL - Prolymphocytic leukaemia|9832/3
C0023486|T191|PT|B64y1|RCD|Prolymphocytic leukaemia|9832/3
C0023486|T191|SY|B64y1|RCDAE|PLL - Prolymphocytic leukemia|9832/3
C0023486|T191|PT|B64y1|RCDAE|Prolymphocytic leukemia|9832/3
C0023486|T191|PT|BBr25|RCDSA|Prolymphocytic leukemia|9832/3
C0023486|T191|PT|BBr25|RCDSY|Prolymphocytic leukaemia|9832/3
C0023486|T191|SYGB|110006004|SNOMEDCT_US|PLL - Prolymphocytic leukaemia|9832/3
C0023486|T191|SY|110006004|SNOMEDCT_US|PLL - Prolymphocytic leukemia|9832/3
C0023486|T191|OAP|10300002|SNOMEDCT_US|Prolymphocytic leukaemia|9832/3
C0023486|T191|PTGB|128923008|SNOMEDCT_US|Prolymphocytic leukaemia|9832/3
C0023486|T191|SYGB|110006004|SNOMEDCT_US|Prolymphocytic leukaemia|9832/3
C0023486|T191|IS|10300002|SNOMEDCT_US|Prolymphocytic leukaemia -RETIRED-|9832/3
C0023486|T191|OAP|10300002|SNOMEDCT_US|Prolymphocytic leukemia|9832/3
C0023486|T191|SY|110006004|SNOMEDCT_US|Prolymphocytic leukemia|9832/3
C0023486|T191|PT|128923008|SNOMEDCT_US|Prolymphocytic leukemia|9832/3
C0023486|T191|IS|10300002|SNOMEDCT_US|Prolymphocytic leukemia -RETIRED-|9832/3
C0023486|T191|OF|10300002|SNOMEDCT_US|Prolymphocytic leukemia -RETIRED-|9832/3
C0475801|T191|AB|C91.3|ICD10CM|Prolymphocytic leukemia of B-cell type|9833/3
C0475801|T191|HT|C91.3|ICD10CM|Prolymphocytic leukemia of B-cell type|9833/3
C0475801|T191|ET|C91.30|ICD10CM|Prolymphocytic leukemia of B-cell type NOS|9833/3
C0475801|T191|LLT|10073480|MDR|B-cell prolymphocytic leukaemia|9833/3
C0475801|T191|PT|10073480|MDR|B-cell prolymphocytic leukaemia|9833/3
C0475801|T191|LLT|10073483|MDR|B-cell prolymphocytic leukemia|9833/3
C0475801|T191|MTH_PT|10073480|MDR|B-cell prolymphocytic leukemia|9833/3
C0475801|T191|PT|230908|MEDCIN|B-cell prolymphocytic leukemia|9833/3
C0475801|T191|SY|230908|MEDCIN|B-cell type prolymphocytic leukemia|9833/3
C0475801|T191|SY|230908|MEDCIN|leukemia prolymphocytic B-cell type|9833/3
C0475801|T191|PM|D054403|MSH|B Cell Prolymphocytic Leukemia|9833/3
C0475801|T191|ET|D054403|MSH|B-Cell Prolymphocytic Leukemia|9833/3
C0475801|T191|PM|D054403|MSH|B-Cell Prolymphocytic Leukemias|9833/3
C0475801|T191|PM|D054403|MSH|Leukemia, B-Cell Prolymphocytic|9833/3
C0475801|T191|MH|D054403|MSH|Leukemia, Prolymphocytic, B-Cell|9833/3
C0475801|T191|PM|D054403|MSH|Leukemias, B-Cell Prolymphocytic|9833/3
C0475801|T191|PM|D054403|MSH|Prolymphocytic Leukemia, B-Cell|9833/3
C0475801|T191|PM|D054403|MSH|Prolymphocytic Leukemias, B-Cell|9833/3
C0475801|T191|SY|C4753|NCI|B Prolymphocytic Leukemia|9833/3
C0475801|T191|PT|C4753|NCI|B-Cell Prolymphocytic Leukemia|9833/3
C0475801|T191|SY|TCGA|NCI|B-Cell Prolymphocytic Leukemia|9833/3
C0475801|T191|AB|Xa0T5|RCD|B-cell prolymphocyt leukaemia|9833/3
C0475801|T191|PT|Xa0T5|RCD|B-cell prolymphocytic leukaemia|9833/3
C0475801|T191|AB|Xa0T5|RCDAE|B-cell prolymphocyt leukemia|9833/3
C0475801|T191|PT|Xa0T5|RCDAE|B-cell prolymphocytic leukemia|9833/3
C0475801|T191|PTGB|277619001|SNOMEDCT_US|B-cell prolymphocytic leukaemia|9833/3
C0475801|T191|PT|277619001|SNOMEDCT_US|B-cell prolymphocytic leukemia|9833/3
C0475801|T191|PTGB|128820007|SNOMEDCT_US|Prolymphocytic leukaemia, B-cell type|9833/3
C0475801|T191|SY|277619001|SNOMEDCT_US|Prolymphocytic leukemia of B-cell type|9833/3
C0475801|T191|PT|128820007|SNOMEDCT_US|Prolymphocytic leukemia, B-cell type|9833/3
C2363142|T191|AB|C91.6|ICD10CM|Prolymphocytic leukemia of T-cell type|9834/3
C2363142|T191|HT|C91.6|ICD10CM|Prolymphocytic leukemia of T-cell type|9834/3
C2363142|T191|ET|C91.60|ICD10CM|Prolymphocytic leukemia of T-cell type NOS|9834/3
C2363142|T191|LLT|10042985|MDR|T-cell prolymphocytic leukaemia|9834/3
C2363142|T191|PT|10042985|MDR|T-cell prolymphocytic leukaemia|9834/3
C2363142|T191|LLT|10042986|MDR|T-cell prolymphocytic leukemia|9834/3
C2363142|T191|MTH_PT|10042985|MDR|T-cell prolymphocytic leukemia|9834/3
C2363142|T191|SY|230909|MEDCIN|leukemia prolymphocytic T-cell type|9834/3
C2363142|T191|PT|230909|MEDCIN|T-cell prolymphocytic leukemia|9834/3
C2363142|T191|SY|230909|MEDCIN|T-cell type prolymphocytic leukemia|9834/3
C2363142|T191|MH|D015461|MSH|Leukemia, Prolymphocytic, T-Cell|9834/3
C2363142|T191|PM|D015461|MSH|Leukemia, T-Cell Prolymphocytic|9834/3
C2363142|T191|PM|D015461|MSH|Leukemias, T-Cell Prolymphocytic|9834/3
C2363142|T191|PM|D015461|MSH|Prolymphocytic Leukemia, T-Cell|9834/3
C2363142|T191|PM|D015461|MSH|Prolymphocytic Leukemias, T-Cell|9834/3
C2363142|T191|PM|D015461|MSH|T Cell Prolymphocytic Leukemia|9834/3
C2363142|T191|ET|D015461|MSH|T-Cell Prolymphocytic Leukemia|9834/3
C2363142|T191|PM|D015461|MSH|T-Cell Prolymphocytic Leukemias|9834/3
C2363142|T191|PN|NOCODE|MTH|T-Cell Prolymphocytic Leukemia|9834/3
C2363142|T191|SY|C4752|NCI|T Cell Prolymphocytic Leukemia|9834/3
C2363142|T191|SY|C4752|NCI|T Prolymphocytic Leukemia|9834/3
C2363142|T191|SY|TCGA|NCI|T-Cell Prolymphocytic Leukemia|9834/3
C2363142|T191|PT|C4752|NCI|T-Cell Prolymphocytic Leukemia|9834/3
C2363142|T191|AB|Xa0S9|RCD|T-cell prolymphocyt leukaemia|9834/3
C2363142|T191|PT|Xa0S9|RCD|T-cell prolymphocytic leukaemia|9834/3
C2363142|T191|AB|Xa0S9|RCDAE|T-cell prolymphocyt leukemia|9834/3
C2363142|T191|PT|Xa0S9|RCDAE|T-cell prolymphocytic leukemia|9834/3
C2363142|T191|PTGB|128821006|SNOMEDCT_US|Prolymphocytic leukaemia, T-cell type|9834/3
C2363142|T191|SY|277567002|SNOMEDCT_US|Prolymphocytic leukemia of T-cell type|9834/3
C2363142|T191|PT|128821006|SNOMEDCT_US|Prolymphocytic leukemia, T-cell type|9834/3
C2363142|T191|PTGB|277567002|SNOMEDCT_US|T-cell prolymphocytic leukaemia|9834/3
C2363142|T191|SYGB|128821006|SNOMEDCT_US|T-cell prolymphocytic leukaemia|9834/3
C2363142|T191|PT|277567002|SNOMEDCT_US|T-cell prolymphocytic leukemia|9834/3
C2363142|T191|SY|128821006|SNOMEDCT_US|T-cell prolymphocytic leukemia|9834/3
C0023449|T191|PT|BI00288|BI|acute lymphocytic leukemia|9835/3
C0023449|T191|PT|0002315|CCPSS|LEUKEMIA ACUTE LYMPHOBLASTIC|9835/3
C0023449|T191|SY|0000007337|CHV|acute leukaemia lymphoblastic|9835/3
C0023449|T191|SY|0000007337|CHV|acute leukemia lymphoblastic|9835/3
C0023449|T191|SY|0000007337|CHV|acute leukemia lymphocytic|9835/3
C0023449|T191|SY|0000007337|CHV|acute leukemia lymphoid|9835/3
C0023449|T191|SY|0000007337|CHV|acute lymphatic leukaemia|9835/3
C0023449|T191|SY|0000007337|CHV|acute lymphatic leukemia|9835/3
C0023449|T191|SY|0000007337|CHV|acute lymphoblastic leukaemia|9835/3
C0023449|T191|SY|0000007337|CHV|acute lymphoblastic leukemia|9835/3
C0023449|T191|SY|0000007337|CHV|acute lymphoblastic leukemias|9835/3
C0023449|T191|SY|0000007337|CHV|acute lymphocytic leukaemia|9835/3
C0023449|T191|SY|0000007337|CHV|acute lymphocytic leukemia|9835/3
C0023449|T191|SY|0000007337|CHV|acute lymphoid leukemia|9835/3
C0023449|T191|SY|0000007337|CHV|leukemia - acute lymphoblastic|9835/3
C0023449|T191|SY|0000007337|CHV|leukemia acute lymphoblastic|9835/3
C0023449|T191|SY|0000056422|CHV|leukemia lymphoblastic|9835/3
C0023449|T191|SY|0000056422|CHV|lymphoblastic leukaemia|9835/3
C0023449|T191|PT|0000056422|CHV|lymphoblastic leukemia|9835/3
C0023449|T191|SY|0000007337|CHV|lymphocytic leukemia acute|9835/3
C0023449|T191|PT|U000011|COSTAR|ACUTE LYMPHOCYTIC LEUKEMIA|9835/3
C0023449|T191|ET|2004-1620|CSP|acute lymphatic leukemia|9835/3
C0023449|T191|ET|2004-1620|CSP|acute lymphoblastic leukemia|9835/3
C0023449|T191|PT|2004-1620|CSP|acute lymphocytic leukemia|9835/3
C0023449|T191|ET|2004-1620|CSP|acute lymphogenous leukemia|9835/3
C0023449|T191|ET|2004-1620|CSP|ALL|9835/3
C0023449|T191|PT|LEUKEMIA ACUTE LYMPHO|CST|ACUTE LYMPHOBLASTIC LEUKEMIA|9835/3
C0023449|T191|GT|LEUKEMIA ACUTE LYMPHO|CST|LEUKEMIA LYMPHOBLASTIC ACUTE|9835/3
C0023449|T191|SY|NOCODE|DXP|ALL|9835/3
C0023449|T191|DI|U001047|DXP|LEUKEMIA, LYMPHOBLASTIC, ACUTE|9835/3
C0023449|T191|SY|NOCODE|DXP|LEUKEMIA, LYMPHOCYTIC, ACUTE|9835/3
C0023449|T191|SY|HP:0006721|HPO|Acute lymphatic leukemia|9835/3
C0023449|T191|PT|HP:0006721|HPO|Acute lymphoblastic leukemia|9835/3
C0023449|T191|SY|HP:0006721|HPO|Acute lymphocytic leukemia|9835/3
C0023449|T191|SY|HP:0006721|HPO|Acute lymphoid leukemia|9835/3
C0023449|T191|PT|C91.0|ICD10|Acute lymphoblastic leukaemia|9835/3
C0023449|T191|PT|C91.0|ICD10AE|Acute lymphoblastic leukemia|9835/3
C0023449|T191|ET|C91.00|ICD10CM|Acute lymphoblastic leukemia NOS|9835/3
C0023449|T191|HT|204.0|ICD9CM|Lymphoid leukemia, acute|9835/3
C0023449|T191|PT|MTHU044762|ICPC2ICD10ENG|leukemia; lymphatic, acute|9835/3
C0023449|T191|PT|MTHU046612|ICPC2ICD10ENG|lymphatic; leukemia, acute|9835/3
C0023449|T191|PTN|B73003|ICPC2P|acute lymphocytic leukaemia|9835/3
C0023449|T191|MTH_PTN|B73003|ICPC2P|acute lymphocytic leukemia|9835/3
C0023449|T191|PT|B73003|ICPC2P|Leukaemia;acute lymphocytic|9835/3
C0023449|T191|MTH_PT|B73003|ICPC2P|Leukemia;acute lymphocytic|9835/3
C1961102|T191|PT|sh85079143|LCH_NW|Lymphoblastic leukemia|9835/3
C0023449|T191|LLT|10000842|MDR|Acute lymphatic leukaemia|9835/3
C0023449|T191|LLT|10000843|MDR|Acute lymphatic leukemia|9835/3
C0023449|T191|LLT|10000844|MDR|Acute lymphoblastic leukaemia|9835/3
C0023449|T191|LLT|10000845|MDR|Acute lymphoblastic leukemia|9835/3
C0023449|T191|PT|10000846|MDR|Acute lymphocytic leukaemia|9835/3
C0023449|T191|LLT|10000846|MDR|Acute lymphocytic leukaemia|9835/3
C0023449|T191|LLT|10000848|MDR|Acute lymphocytic leukemia|9835/3
C0023449|T191|MTH_PT|10000846|MDR|Acute lymphocytic leukemia|9835/3
C0023449|T191|LLT|10000849|MDR|Acute lymphoid leukaemia|9835/3
C0023449|T191|LLT|10060555|MDR|Acute lymphoid leukemia|9835/3
C0023449|T191|OL|10001690|MDR|ALL|9835/3
C0023449|T191|LLT|10060390|MDR|Leukaemia lymphoblastic acute|9835/3
C0023449|T191|HT|10024290|MDR|Leukaemias acute lymphocytic|9835/3
C0023449|T191|LLT|10024338|MDR|Leukemia lymphoblastic acute|9835/3
C0023449|T191|MTH_HT|10024290|MDR|Leukemias acute lymphocytic|9835/3
C0023449|T191|LLT|10025301|MDR|Lymphoid leukaemia, acute|9835/3
C0023449|T191|LLT|10025305|MDR|Lymphoid leukemia, acute|9835/3
C0023449|T191|PT|31478|MEDCIN|acute lymphocytic leukemia|9835/3
C1961102|T191|SY|230910|MEDCIN|leukemia precursor cell lymphoblastic|9835/3
C1961102|T191|PT|230910|MEDCIN|precursor cell lymphoblastic leukemia|9835/3
C0023449|T191|ET|1437|MEDLINEPLUS|Acute Lymphoblastic Leukemia|9835/3
C0023449|T191|SY|1437|MEDLINEPLUS|Acute lymphoblastic leukemia|9835/3
C0023449|T191|PT|1437|MEDLINEPLUS|Acute Lymphocytic Leukemia|9835/3
C0023449|T191|ET|1437|MEDLINEPLUS|ALL|9835/3
C0023449|T191|SY|1437|MEDLINEPLUS|ALL|9835/3
C1961102|T191|ET|1437|MEDLINEPLUS|Leukemia, Acute Lymphoblastic|9835/3
C0023449|T191|ET|1437|MEDLINEPLUS|Leukemia, Acute Lymphocytic|9835/3
C1961102|T191|PM|D054198|MSH|Acute Lymphoblastic Leukemia|9835/3
C1961102|T191|PM|D054198|MSH|Acute Lymphocytic Leukemia|9835/3
C1961102|T191|ET|D054198|MSH|Acute Lymphoid Leukemia|9835/3
C1961102|T191|ET|D054198|MSH|Leukemia, Acute Lymphoblastic|9835/3
C1961102|T191|PM|D054198|MSH|Leukemia, Acute Lymphocytic|9835/3
C1961102|T191|PM|D054198|MSH|Leukemia, Acute Lymphoid|9835/3
C1961102|T191|ET|D054198|MSH|Leukemia, Lymphoblastic|9835/3
C1961102|T191|ET|D054198|MSH|Leukemia, Lymphoblastic, Acute|9835/3
C1961102|T191|ET|D054198|MSH|Leukemia, Lymphocytic, Acute|9835/3
C1961102|T191|ET|D054198|MSH|Leukemia, Lymphoid, Acute|9835/3
C1961102|T191|ET|D054198|MSH|Lymphoblastic Leukemia|9835/3
C1961102|T191|ET|D054198|MSH|Lymphoblastic Leukemia, Acute|9835/3
C1961102|T191|ET|D054198|MSH|Lymphoblastic Lymphoma|9835/3
C1961102|T191|ET|D054198|MSH|Lymphocytic Leukemia, Acute|9835/3
C1961102|T191|PM|D054198|MSH|Lymphoid Leukemia, Acute|9835/3
C1961102|T191|ET|D054198|MSH|Lymphoma, Lymphoblastic|9835/3
C1961102|T191|PM|D054198|MSH|Precursor Cell Lymphoblastic Leukemia Lymphoma|9835/3
C1961102|T191|MH|D054198|MSH|Precursor Cell Lymphoblastic Leukemia-Lymphoma|9835/3
C0023449|T191|PN|NOCODE|MTH|Acute lymphocytic leukemia|9835/3
C1961102|T191|PN|NOCODE|MTH|Precursor Cell Lymphoblastic Leukemia Lymphoma|9835/3
C0023449|T191|PT|C3167|NCI|Acute Lymphoblastic Leukemia|9835/3
C0023449|T191|OP|C3167|NCI|Acute Lymphocytic Leukaemia|9835/3
C0023449|T191|OP|C3167|NCI|Acute Lymphocytic Leukemia|9835/3
C0023449|T191|OP|C3167|NCI|Acute Lymphocytic Leukemias|9835/3
C0023449|T191|OP|C3167|NCI|Acute Lymphogenous Leukemia|9835/3
C0023449|T191|SY|C3167|NCI|Acute Lymphoid Leukemia|9835/3
C0023449|T191|AB|C3167|NCI|ALL|9835/3
C0023449|T191|SY|C3167|NCI|ALL - Acute Lymphocytic Leukemia|9835/3
C0023449|T191|SY|C3167|NCI|Lymphoblastic Leukemia|9835/3
C0023449|T191|SY|C3167|NCI|Precursor Cell Lymphoblastic Leukemia|9835/3
C0023449|T191|SY|C3167|NCI|Precursor Lymphoblastic Leukemia|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|Acute Lymphocytic Leukaemia|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|Acute Lymphocytic Leukemias|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|Acute Lymphogenous Leukemia|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|Acute Lymphoid Leukemia|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|ALL|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|ALL - Acute Lymphocytic Leukemia|9835/3
C0023449|T191|PT|C3167|NCI_CDISC|LEUKEMIA, LYMPHOBLASTIC, MALIGNANT|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|Lymphoblastic Leukemia|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|Precursor Cell Lymphoblastic Leukemia|9835/3
C0023449|T191|SY|C3167|NCI_CDISC|Precursor Lymphoblasic Leukemia|9835/3
C0023449|T191|PT|C3167|NCI_CPTAC|Acute Lymphoblastic Leukemia|9835/3
C0023449|T191|SY|10000846|NCI_CTEP-SDC|Acute lymphoblastic leukemia|9835/3
C0023449|T191|PT|10000846|NCI_CTEP-SDC|Acute lymphoblastic leukemia, NOS|9835/3
C0023449|T191|SY|C3167|NCI_CTRP|Acute Lymphoblastic Leukemia|9835/3
C0023449|T191|PT|CDR0000045586|NCI_NCI-GLOSS|acute lymphoblastic leukemia|9835/3
C0023449|T191|PT|CDR0000046332|NCI_NCI-GLOSS|acute lymphocytic leukemia|9835/3
C0023449|T191|PT|CDR0000044362|NCI_NCI-GLOSS|ALL|9835/3
C0023449|T191|PT|C3167|NCI_NICHD|Acute Lymphoblastic Leukemia|9835/3
C0023449|T191|SY|C3167|NCI_NICHD|Acute Lymphocytic Leukemia|9835/3
C0023449|T191|SY|CDR0000043423|PDQ|Acute Lymphoblastic Leukemia|9835/3
C0023449|T191|IS|CDR0000043423|PDQ|Acute Lymphocytic Leukaemia|9835/3
C0023449|T191|PT|CDR0000043423|PDQ|acute lymphocytic leukemia|9835/3
C0023449|T191|SY|CDR0000043423|PDQ|Acute Lymphocytic Leukemias|9835/3
C0023449|T191|SY|CDR0000043423|PDQ|Acute Lymphogenous Leukemia|9835/3
C0023449|T191|SY|CDR0000043423|PDQ|Acute Lymphoid Leukemia|9835/3
C0023449|T191|AB|CDR0000043423|PDQ|ALL|9835/3
C0023449|T191|SY|CDR0000043423|PDQ|ALL - Acute Lymphocytic Leukemia|9835/3
C0023449|T191|SY|CDR0000043423|PDQ|leukemia, acute lymphocytic|9835/3
C0023449|T191|SY|CDR0000043423|PDQ|Lymphoblastic Leukemia|9835/3
C1961102|T191|SY|CDR0000043423|PDQ|Precursor Cell Lymphoblastic Leukemia|9835/3
C1961102|T191|SY|CDR0000043423|PDQ|Precursor Lymphoblastic Leukemia|9835/3
C0023449|T191|PT|R0121660|QMR|LEUKEMIA ACUTE LYMPHOBLASTIC|9835/3
C0023449|T191|SY|B640.|RCD|Acute lymphatic leukaemia|9835/3
C0023449|T191|SY|B640.|RCD|Acute lymphoblastic leukaemia|9835/3
C0023449|T191|PT|B640.|RCD|Acute lymphoid leukaemia|9835/3
C0023449|T191|AB|B640.|RCD|ALL - Acute lymphobl leukaemia|9835/3
C0023449|T191|SY|B640.|RCD|ALL - Acute lymphoblastic leukaemia|9835/3
C0023449|T191|SY|B640.|RCDAE|Acute lymphatic leukemia|9835/3
C0023449|T191|SY|B640.|RCDAE|Acute lymphoblastic leukemia|9835/3
C0023449|T191|PT|B640.|RCDAE|Acute lymphoid leukemia|9835/3
C0023449|T191|AB|B640.|RCDAE|ALL - Acute lymphobl leukemia|9835/3
C0023449|T191|SY|B640.|RCDAE|ALL - Acute lymphoblastic leukemia|9835/3
C0023449|T191|PT|BBr21|RCDSA|Acute lymphoid leukemia|9835/3
C0023449|T191|PT|BBr21|RCDSY|Acute lymphoid leukaemia|9835/3
C0023449|T191|SYGB|128822004|SNOMEDCT_US|Acute lymphatic leukaemia|9835/3
C0023449|T191|IS|90151006|SNOMEDCT_US|Acute lymphatic leukemia|9835/3
C0023449|T191|SY|128822004|SNOMEDCT_US|Acute lymphatic leukemia|9835/3
C0023449|T191|SYGB|128822004|SNOMEDCT_US|Acute lymphoblastic leukaemia|9835/3
C1531702|T191|PTGB|413440007|SNOMEDCT_US|Acute lymphoblastic leukaemia - category|9835/3
C0023449|T191|IS|90151006|SNOMEDCT_US|Acute lymphoblastic leukaemia -RETIRED-|9835/3
C0023449|T191|SYGB|128822004|SNOMEDCT_US|Acute lymphoblastic leukaemia-lymphoma|9835/3
C1961102|T191|SYGB|128822004|SNOMEDCT_US|Acute lymphoblastic leukaemia, precursor-cell type|9835/3
C0023449|T191|OAP|90151006|SNOMEDCT_US|Acute lymphoblastic leukemia|9835/3
C0023449|T191|SY|128822004|SNOMEDCT_US|Acute lymphoblastic leukemia|9835/3
C1531702|T191|PT|413440007|SNOMEDCT_US|Acute lymphoblastic leukemia - category|9835/3
C0023449|T191|IS|90151006|SNOMEDCT_US|Acute lymphoblastic leukemia -RETIRED-|9835/3
C0023449|T191|OF|90151006|SNOMEDCT_US|Acute lymphoblastic leukemia -RETIRED-|9835/3
C0023449|T191|SY|128822004|SNOMEDCT_US|Acute lymphoblastic leukemia-lymphoma|9835/3
C0023449|T191|IS|90151006|SNOMEDCT_US|Acute lymphoblastic leukemia, NOS|9835/3
C1961102|T191|SY|128822004|SNOMEDCT_US|Acute lymphoblastic leukemia, precursor-cell type|9835/3
C0023449|T191|SYGB|128822004|SNOMEDCT_US|Acute lymphocytic leukaemia|9835/3
C0023449|T191|SY|128822004|SNOMEDCT_US|Acute lymphocytic leukemia|9835/3
C0023449|T191|IS|90151006|SNOMEDCT_US|Acute lymphocytic leukemia|9835/3
C0023449|T191|PTGB|91857003|SNOMEDCT_US|Acute lymphoid leukaemia|9835/3
C0023449|T191|SYGB|91857003|SNOMEDCT_US|Acute lymphoid leukaemia, disease|9835/3
C0023449|T191|PT|91857003|SNOMEDCT_US|Acute lymphoid leukemia|9835/3
C0023449|T191|SY|91857003|SNOMEDCT_US|Acute lymphoid leukemia, disease|9835/3
C0023449|T191|SYGB|91857003|SNOMEDCT_US|ALL - Acute lymphoblastic leukaemia|9835/3
C0023449|T191|SY|91857003|SNOMEDCT_US|ALL - Acute lymphoblastic leukemia|9835/3
C0023449|T191|SYGB|128822004|SNOMEDCT_US|Lymphoblastic leukaemia|9835/3
C0023449|T191|SY|128822004|SNOMEDCT_US|Lymphoblastic leukemia|9835/3
C0023449|T191|IS|90151006|SNOMEDCT_US|Lymphoblastic leukemia, NOS|9835/3
C1961102|T191|PTGB|128822004|SNOMEDCT_US|Precursor cell lymphoblastic leukaemia|9835/3
C1961102|T191|SYGB|128822004|SNOMEDCT_US|Precursor cell lymphoblastic leukaemia, not phenotyped|9835/3
C1961102|T191|PT|128822004|SNOMEDCT_US|Precursor cell lymphoblastic leukemia|9835/3
C1961102|T191|SY|128822004|SNOMEDCT_US|Precursor cell lymphoblastic leukemia, not phenotyped|9835/3
C1292769|T191|SY|0000057459|CHV|c all|9836/3
C1292769|T191|SY|0000057459|CHV|pre-b|9836/3
C1292769|T191|PT|0000057459|CHV|precursor b-cell lymphoblastic leukemia|9836/3
C1292769|T191|SY|0000057459|CHV|pro b|9836/3
C1292769|T191|LLT|10003917|MDR|B-cell type acute leukaemia|9836/3
C1292769|T191|PT|10003917|MDR|B-cell type acute leukaemia|9836/3
C1292769|T191|LLT|10003918|MDR|B-cell type acute leukaemia NOS|9836/3
C1292769|T191|LLT|10003919|MDR|B-cell type acute leukemia|9836/3
C1292769|T191|MTH_PT|10003917|MDR|B-cell type acute leukemia|9836/3
C1292769|T191|LLT|10003920|MDR|B-cell type acute leukemia NOS|9836/3
C1292769|T191|PT|339623|MEDCIN|B-cell acute lymphocytic leukemia|9836/3
C1292769|T191|SY|230911|MEDCIN|leukemia precursor cell lymphoblastic B-cell|9836/3
C1292769|T191|PT|230911|MEDCIN|precursor B-cell lymphoblastic leukemia|9836/3
C1292769|T191|PN|NOCODE|MTH|Precursor B-cell lymphoblastic leukemia|9836/3
C1292769|T191|OP|C8644|NCI|Acute B Cell Lymphocytic Leukemia|9836/3
C1292769|T191|OP|C8644|NCI|Acute B-Cell Lymphocytic Leukemia|9836/3
C1292769|T191|PT|C8644|NCI|B Acute Lymphoblastic Leukemia|9836/3
C1292769|T191|OP|C8644|NCI|B Cell Acute Lymphocytic Leukemia|9836/3
C1292769|T191|SY|C8644|NCI|B Cell Precursor Type Acute Leukemia|9836/3
C4329382|T191|SY|C129787|NCI|B Lymphoblastic Leukemia/Lymphoma with Translocations Involving Tyrosine Kinases or Cytokine Receptors|9836/3
C4329382|T191|PT|C129787|NCI|B Lymphoblastic Leukemia/Lymphoma, BCR-ABL1-Like|9836/3
C1292769|T191|AB|C8644|NCI|B-ALL|9836/3
C1292769|T191|SY|C8644|NCI|B-Cell Acute Lymphoblastic Leukemia|9836/3
C1292769|T191|OP|C8644|NCI|B-Cell Acute Lymphocytic Leukemia|9836/3
C1292769|T191|SY|C8644|NCI|B-Cell Lymphoblastic Leukemia|9836/3
C1292769|T191|SY|C8644|NCI|B-Cell Precursor Type Acute Leukemia|9836/3
C1292769|T191|SY|C8644|NCI|B-Cell Type Acute Leukemia|9836/3
C1292769|T191|SY|C8644|NCI|Precursor B-Lymphoblastic Leukemia|9836/3
C1292769|T191|SY|10003890|NCI_CTEP-SDC|B-precursor ALL|9836/3
C1292769|T191|SY|CDR0000543504|NCI_NCI-GLOSS|B-cell acute lymphoblastic leukemia|9836/3
C1292769|T191|PT|CDR0000543509|NCI_NCI-GLOSS|B-cell acute lymphocytic leukemia|9836/3
C1292769|T191|SY|CDR0000524192|NCI_NCI-GLOSS|precursor B-lymphoblastic leukemia|9836/3
C1292769|T191|PT|C8644|NCI_NICHD|B Acute Lymphoblastic Leukemia|9836/3
C1292769|T191|SY|C8644|NCI_NICHD|B-ALL|9836/3
C1292769|T191|AB|Xa0SD|RCD|B-cell acute lymphob leukaemia|9836/3
C1292769|T191|PT|Xa0SD|RCD|B-cell acute lymphoblastic leukaemia|9836/3
C1292769|T191|AB|Xa0SD|RCDAE|B-cell acute lymphob leukemia|9836/3
C1292769|T191|PT|Xa0SD|RCDAE|B-cell acute lymphoblastic leukemia|9836/3
C1292769|T191|PT|277571004|SNOMEDCT_US|B-cell acute lymphoblastic leukemia|9836/3
C4329382|T191|PTGB|783744003|SNOMEDCT_US|B-lymphoblastic leukaemia lymphoma BCR-ABL1-like|9836/3
C4329382|T191|PT|783744003|SNOMEDCT_US|B-lymphoblastic leukemia lymphoma BCR-ABL1-like|9836/3
C1292769|T191|SY|128823009|SNOMEDCT_US|c-ALL|9836/3
C1292769|T191|SY|128823009|SNOMEDCT_US|Common ALL|9836/3
C1292769|T191|SY|128823009|SNOMEDCT_US|Common precursor B ALL|9836/3
C1292769|T191|SYGB|277571004|SNOMEDCT_US|Mature B-cell leukaemia Burkitt type|9836/3
C1292769|T191|SY|277571004|SNOMEDCT_US|Mature B-cell leukemia Burkitt type|9836/3
C1292769|T191|SY|128823009|SNOMEDCT_US|Pre-B ALL|9836/3
C1292769|T191|SY|128823009|SNOMEDCT_US|Pre-pre-B ALL|9836/3
C1292769|T191|PTGB|128823009|SNOMEDCT_US|Precursor B-cell lymphoblastic leukaemia|9836/3
C1292769|T191|PT|128823009|SNOMEDCT_US|Precursor B-cell lymphoblastic leukemia|9836/3
C1292769|T191|SY|128823009|SNOMEDCT_US|Pro-B ALL|9836/3
C1961099|T191|ET|2004-1803|CSP|acute T cell leukemia|9837/3
C1961099|T191|ET|2004-1600|CSP|acute T cell leukemia|9837/3
C1961099|T191|PT|HP:0006727|HPO|T-cell acute lymphoblastic leukemias|9837/3
C1301359|T191|LLT|10036543|MDR|Precursor T-lymphoblastic lymphoma/leukaemia|9837/3
C1301359|T191|PT|10036543|MDR|Precursor T-lymphoblastic lymphoma/leukaemia|9837/3
C1301359|T191|LLT|10036545|MDR|Precursor T-lymphoblastic lymphoma/leukaemia NOS|9837/3
C1301359|T191|LLT|10054569|MDR|Precursor T-lymphoblastic lymphoma/leukemia|9837/3
C1301359|T191|MTH_PT|10036543|MDR|Precursor T-lymphoblastic lymphoma/leukemia|9837/3
C1301359|T191|LLT|10054570|MDR|Precursor T-lymphoblastic lymphoma/leukemia NOS|9837/3
C1301359|T191|HT|10036544|MDR|Precursor T-lymphoblastic lymphomas/leukaemias|9837/3
C1301359|T191|MTH_HT|10036544|MDR|Precursor T-lymphoblastic lymphomas/leukemias|9837/3
C1961099|T191|LLT|10066105|MDR|T-cell lymphoblastic leukaemia acute|9837/3
C1961099|T191|LLT|10066110|MDR|T-cell lymphoblastic leukemia acute|9837/3
C1961099|T191|LLT|10042987|MDR|T-cell type acute leukaemia|9837/3
C1961099|T191|PT|10042987|MDR|T-cell type acute leukaemia|9837/3
C1961099|T191|LLT|10054655|MDR|T-cell type acute leukemia|9837/3
C1961099|T191|MTH_PT|10042987|MDR|T-cell type acute leukemia|9837/3
C1961099|T191|SY|230912|MEDCIN|leukemia precursor cell lymphoblastic T-cell|9837/3
C1301359|T191|PT|355493|MEDCIN|malignant precursor T-cell lymphoblastic leukemia or lymphoma|9837/3
C1961099|T191|PT|230912|MEDCIN|precursor T-cell lymphoblastic leukemia|9837/3
C1301359|T191|SY|355493|MEDCIN|precursor T-cell lymphoblastic leukemia or lymphoma|9837/3
C1961099|T191|PT|339627|MEDCIN|T-cell acute lymphoblastic leukemia|9837/3
C1961099|T191|PM|D054218|MSH|Acute T-Cell Leukemia|9837/3
C1961099|T191|PM|D054218|MSH|Acute T-Cell Leukemias|9837/3
C1961099|T191|PM|D054218|MSH|Acute T-Lymphocytic Leukemia|9837/3
C1961099|T191|PM|D054218|MSH|Acute T-Lymphocytic Leukemias|9837/3
C1961099|T191|PM|D054218|MSH|Leukemia, Acute T-Cell|9837/3
C1961099|T191|PM|D054218|MSH|Leukemia, Acute T-Lymphocytic|9837/3
C1961099|T191|ET|D054218|MSH|Leukemia, Lymphoblastic, Acute, T Cell|9837/3
C1961099|T191|ET|D054218|MSH|Leukemia, Lymphoblastic, Acute, T-Cell|9837/3
C1961099|T191|ET|D054218|MSH|Leukemia, Lymphocytic, Acute T Cell|9837/3
C1961099|T191|ET|D054218|MSH|Leukemia, Lymphocytic, Acute, T-Cell|9837/3
C1961099|T191|ET|D054218|MSH|Leukemia, T-Cell, Acute|9837/3
C1961099|T191|PM|D054218|MSH|Leukemias, Acute T-Cell|9837/3
C1961099|T191|PM|D054218|MSH|Leukemias, Acute T-Lymphocytic|9837/3
C1961099|T191|ET|D054218|MSH|Lymphoblastic Leukemia, Acute, T Cell|9837/3
C1961099|T191|ET|D054218|MSH|Lymphoblastic Leukemia, Acute, T-Cell|9837/3
C1961099|T191|DSV|D054218|MSH|LYMPHOCYTIC LEUKEMIA ACUTE BT|9837/3
C1961099|T191|ET|D054218|MSH|Lymphocytic Leukemia, T Cell, Acute|9837/3
C1961099|T191|ET|D054218|MSH|Lymphocytic Leukemia, T-Cell, Acute|9837/3
C1961099|T191|PM|D054218|MSH|Precursor T Cell Lymphoblastic Leukemia|9837/3
C1961099|T191|PM|D054218|MSH|Precursor T Cell Lymphoblastic Leukemia Lymphoma|9837/3
C1961099|T191|PM|D054218|MSH|Precursor T Cell Lymphoblastic Lymphoma|9837/3
C1961099|T191|ET|D054218|MSH|Precursor T-Cell Lymphoblastic Leukemia|9837/3
C1961099|T191|MH|D054218|MSH|Precursor T-Cell Lymphoblastic Leukemia-Lymphoma|9837/3
C1961099|T191|ET|D054218|MSH|Precursor T-Cell Lymphoblastic Lymphoma|9837/3
C1961099|T191|PM|D054218|MSH|T Cell Leukemia, Acute|9837/3
C1961099|T191|PM|D054218|MSH|T Lymphocytic Leukemia, Acute|9837/3
C1961099|T191|ET|D054218|MSH|T-ALL|9837/3
C1961099|T191|ET|D054218|MSH|T-Cell Acute Lymphocytic Leukemia|9837/3
C1961099|T191|ET|D054218|MSH|T-Cell Leukemia, Acute|9837/3
C1961099|T191|PM|D054218|MSH|T-Cell Leukemias, Acute|9837/3
C1961099|T191|ET|D054218|MSH|T-Lymphocytic Leukemia, Acute|9837/3
C1961099|T191|PM|D054218|MSH|T-Lymphocytic Leukemias, Acute|9837/3
C1961099|T191|PN|NOCODE|MTH|Precursor T-Cell Lymphoblastic Leukemia-Lymphoma|9837/3
C1961099|T191|SY|C3183|NCI|Acute T Cell Leukemia|9837/3
C1961099|T191|SY|C3183|NCI|Acute T Cell Lymphoblastic Leukemia|9837/3
C1961099|T191|OP|C3183|NCI|Acute T Cell Lymphocytic Leukemia|9837/3
C1961099|T191|SY|C3183|NCI|Acute T-Cell Leukemia|9837/3
C1961099|T191|SY|C3183|NCI|Acute T-Cell Lymphoblastic Leukemia|9837/3
C1961099|T191|OP|C3183|NCI|Acute T-Cell Lymphocytic Leukemia|9837/3
C2826059|T191|PT|C82217|NCI|Natural Killer Cell Lymphoblastic Leukemia/Lymphoma|9837/3
C2826059|T191|SY|C82217|NCI|NK Cell Lymphoblastic Leukemia/Lymphoma|9837/3
C2826059|T191|SY|C82217|NCI|NK Lymphoblastic Leukemia/Lymphoma|9837/3
C2826059|T191|AB|C82217|NCI|NK-ALL/LBL|9837/3
C2826059|T191|SY|C82217|NCI|NK-Lymphoblastic Leukemia/Lymphoma|9837/3
C1961099|T191|OP|C27261|NCI|Pre T-ALL|9837/3
C1961099|T191|PT|C27261|NCI|Pre T-ALL|9837/3
C2826059|T191|SY|C82217|NCI|Precursor Natural Killer Cell Lymphoblastic Leukemia/Lymphoma|9837/3
C2826059|T191|SY|C82217|NCI|Precursor NK Cell Lymphoblastic Leukemia/Lymphoma|9837/3
C1301359|T191|SY|C8694|NCI|Precursor T Lymphoblastic Leukemia/Lymphoma|9837/3
C1301359|T191|SY|C8694|NCI|Precursor T Lymphoblastic Lymphoma/Leukemia|9837/3
C1961099|T191|SY|C3183|NCI|Precursor T-Lymphoblastic Leukemia|9837/3
C1301359|T191|SY|C8694|NCI|Precursor T-Lymphoblastic Lymphoma/Leukemia|9837/3
C1961099|T191|PT|C3183|NCI|T Acute Lymphoblastic Leukemia|9837/3
C1301359|T191|PT|C8694|NCI|T Lymphoblastic Leukemia/Lymphoma|9837/3
C1301359|T191|SY|TCGA|NCI|T Lymphoblastic Leukemia/Lymphoma|9837/3
C1961099|T191|AB|C3183|NCI|T-ALL|9837/3
C1961099|T191|SY|C3183|NCI|T-Cell Acute Lymphoblastic Leukemia|9837/3
C1961099|T191|SY|C3183|NCI|T-Cell Type Acute Leukemia|9837/3
C1301359|T191|SY|C8694|NCI|T-Lymphoblastic Leukemia/Lymphoma|9837/3
C1961099|T191|SY|10054569|NCI_CTEP-SDC|T-cell ALL|9837/3
C1301359|T191|DN|C8694|NCI_CTRP|T Lymphoblastic Leukemia/Lymphoma|9837/3
C1961099|T191|SY|CDR0000509729|NCI_NCI-GLOSS|precursor T-lymphoblastic leukemia|9837/3
C1961099|T191|PT|CDR0000509731|NCI_NCI-GLOSS|T-cell acute lymphoblastic leukemia|9837/3
C1961099|T191|SY|CDR0000509747|NCI_NCI-GLOSS|T-cell acute lymphocytic leukemia|9837/3
C1961099|T191|PT|C3183|NCI_NICHD|T Acute Lymphoblastic Leukemia|9837/3
C1961099|T191|SY|C3183|NCI_NICHD|T-ALL|9837/3
C1961099|T191|AB|Xa0SH|RCD|T-cell acute lymphobl leukaem|9837/3
C1961099|T191|PT|Xa0SH|RCD|T-cell acute lymphoblastic leukaemia|9837/3
C1961099|T191|PT|Xa0SH|RCDAE|T-cell acute lymphoblastic leukemia|9837/3
C1961099|T191|SYGB|277575008|SNOMEDCT_US|Acute T-cell lymphoblastic leukaemia|9837/3
C1961099|T191|SY|277575008|SNOMEDCT_US|Acute T-cell lymphoblastic leukemia|9837/3
C1961099|T191|SY|128824003|SNOMEDCT_US|Cortical T ALL|9837/3
C2826059|T191|SYGB|783414002|SNOMEDCT_US|Natural killer-lymphoblastic leukaemia/lymphoma|9837/3
C2826059|T191|SY|783414002|SNOMEDCT_US|Natural killer-lymphoblastic leukemia/lymphoma|9837/3
C2826059|T191|PTGB|783414002|SNOMEDCT_US|NK-lymphoblastic leukaemia/lymphoma|9837/3
C2826059|T191|PT|783414002|SNOMEDCT_US|NK-lymphoblastic leukemia/lymphoma|9837/3
C1961099|T191|SY|128824003|SNOMEDCT_US|Pre-T ALL|9837/3
C1301359|T191|PT|420890002|SNOMEDCT_US|Precursor T cell lymphoblastic leukemia/lymphoblastic lymphoma|9837/3
C1301359|T191|PT|397348006|SNOMEDCT_US|Precursor T cell lymphoblastic leukemia/lymphoblastic lymphoma|9837/3
C1961099|T191|PTGB|128824003|SNOMEDCT_US|Precursor T-cell lymphoblastic leukaemia|9837/3
C1961099|T191|SYGB|277575008|SNOMEDCT_US|Precursor T-cell lymphoblastic leukaemia|9837/3
C1961099|T191|PT|128824003|SNOMEDCT_US|Precursor T-cell lymphoblastic leukemia|9837/3
C1961099|T191|SY|277575008|SNOMEDCT_US|Precursor T-cell lymphoblastic leukemia|9837/3
C1961099|T191|SY|128824003|SNOMEDCT_US|Pro-T ALL|9837/3
C1301359|T191|PTGB|703821009|SNOMEDCT_US|T lymphoblastic leukaemia/lymphoma|9837/3
C1301359|T191|PT|703821009|SNOMEDCT_US|T lymphoblastic leukemia/lymphoma|9837/3
C1961099|T191|PTGB|277575008|SNOMEDCT_US|T-cell acute lymphoblastic leukaemia|9837/3
C1961099|T191|PT|277575008|SNOMEDCT_US|T-cell acute lymphoblastic leukemia|9837/3
C1301359|T191|SYGB|397348006|SNOMEDCT_US|T-lymphoblastic lymphoma/leukaemia|9837/3
C1301359|T191|SY|397348006|SNOMEDCT_US|T-lymphoblastic lymphoma/leukemia|9837/3
C0023440|T191|SY|0000007334|CHV|acute erythroblastic leukemia|9840/3
C0023440|T191|SY|0000007334|CHV|aml m6|9840/3
C0023440|T191|SY|0000007334|CHV|di guglielmo disease|9840/3
C0023440|T191|SY|0000007334|CHV|diguglielmo's syndrome|9840/3
C0023440|T191|SY|0000007334|CHV|erythremic myelosis|9840/3
C0023440|T191|SY|0000007334|CHV|erythroid leukemia acute|9840/3
C0023440|T191|SY|0000007334|CHV|erythroleukaemia|9840/3
C0023440|T191|PT|0000007334|CHV|erythroleukemia|9840/3
C0023440|T191|ET|2004-1746|CSP|DiGugliemo syndrome|9840/3
C0023440|T191|ET|2004-1746|CSP|erythremic myelosis|9840/3
C0023440|T191|PT|2004-1746|CSP|erythroleukemia|9840/3
C0023440|T191|GT|MARROW HYPERPLASIA|CST|DI GUGLIELMO'S SYNDROME|9840/3
C0023440|T191|GT|MARROW HYPERPLASIA|CST|ERYTHREMIC MYELOSIS|9840/3
C0023440|T191|GT|LEUKEMIA|CST|ERYTHROLEUKEMIA|9840/3
C0023440|T191|GT|MARROW HYPERPLASIA|CST|MYELOSIS ERYTHREMIC|9840/3
C0023440|T191|GT|MARROW HYPERPLASIA|CST|SYNDROME DIGUGLIELMO'S|9840/3
C0023440|T191|SY|NOCODE|DXP|DI GUGLIELMO SYNDROME|9840/3
C0023440|T191|SY|NOCODE|DXP|DIGUGLIELMO DISEASE|9840/3
C0023440|T191|DI|U000593|DXP|ERYTHROLEUKEMIA|9840/3
C0023440|T191|AB|C94.0|ICD10CM|Acute erythroid leukemia|9840/3
C0023440|T191|HT|C94.0|ICD10CM|Acute erythroid leukemia|9840/3
C0023440|T191|ET|C94.00|ICD10CM|Acute erythroid leukemia NOS|9840/3
C0023440|T191|ET|C94.0|ICD10CM|Erythroleukemia|9840/3
C0023440|T191|PT|MTHU022754|ICPC2ICD10ENG|Di Guglielmo|9840/3
C0023440|T191|PT|MTHU027041|ICPC2ICD10ENG|erythremic; myelosis|9840/3
C0023440|T191|PT|MTHU027042|ICPC2ICD10ENG|erythremic; myelosis, acute|9840/3
C0023440|T191|PT|MTHU027066|ICPC2ICD10ENG|erythroleukemia|9840/3
C0023440|T191|PT|MTHU050920|ICPC2ICD10ENG|myelosis; erythremic|9840/3
C0023440|T191|PT|MTHU050921|ICPC2ICD10ENG|myelosis; erythremic, acute|9840/3
C0023440|T191|LLT|10000739|MDR|Acute erythroid leukaemia|9840/3
C0023440|T191|LLT|10000740|MDR|Acute erythroid leukemia|9840/3
C0023440|T191|LLT|10012593|MDR|Di Guglielmo's syndrome|9840/3
C0023440|T191|LLT|10015245|MDR|Erythraemic myelosis|9840/3
C0023440|T191|LLT|10015249|MDR|Erythremic myelosis|9840/3
C0023440|T191|LLT|10015281|MDR|Erythroleukaemia|9840/3
C0023440|T191|PT|10015281|MDR|Erythroleukaemia|9840/3
C0023440|T191|LLT|10015282|MDR|Erythroleukemia|9840/3
C0023440|T191|MTH_PT|10015281|MDR|Erythroleukemia|9840/3
C0023440|T191|LLT|10060401|MDR|Myelosis erythraemic|9840/3
C0023440|T191|LLT|10028579|MDR|Myelosis erythremic|9840/3
C0023440|T191|LLT|10042799|MDR|Syndrome DiGuglielmo's|9840/3
C0023440|T191|PT|230913|MEDCIN|acute myelogenous leukemia M6 type|9840/3
C0023440|T191|SY|230913|MEDCIN|AML M6 type|9840/3
C0023440|T191|SY|31472|MEDCIN|di Guglielmo's disease|9840/3
C0023440|T191|PT|31472|MEDCIN|erythroleukemia|9840/3
C0023440|T191|PM|D004915|MSH|Acute Erythroblastic Leukemia|9840/3
C0023440|T191|PM|D004915|MSH|Acute Erythroblastic Leukemias|9840/3
C0023440|T191|DEV|D004915|MSH|DI GUGLIELMO DIS|9840/3
C0023440|T191|ET|D004915|MSH|Di Guglielmo Disease|9840/3
C0023440|T191|ET|D004915|MSH|Di Guglielmo's Disease|9840/3
C0023440|T191|DEV|D004915|MSH|DI GUGLIELMOS DIS|9840/3
C0023440|T191|PM|D004915|MSH|Di Guglielmos Disease|9840/3
C0023440|T191|PM|D004915|MSH|Disease, Di Guglielmo|9840/3
C0023440|T191|PM|D004915|MSH|Disease, Di Guglielmo's|9840/3
C0023440|T191|PM|D004915|MSH|Erythremic Myeloses|9840/3
C0023440|T191|ET|D004915|MSH|Erythremic Myelosis|9840/3
C0023440|T191|ET|D004915|MSH|Erythroblastic Leukemia, Acute|9840/3
C0023440|T191|PM|D004915|MSH|Erythroblastic Leukemias, Acute|9840/3
C0023440|T191|ET|D004915|MSH|Erythroleukemia|9840/3
C0023440|T191|PM|D004915|MSH|Erythroleukemias|9840/3
C0023440|T191|DSV|D004915|MSH|LEUKEMIA MYELOID ACUTE M 06|9840/3
C0023440|T191|PM|D004915|MSH|Leukemia, Acute Erythroblastic|9840/3
C0023440|T191|MH|D004915|MSH|Leukemia, Erythroblastic, Acute|9840/3
C0023440|T191|ET|D004915|MSH|Leukemia, Myeloid, Acute, M6|9840/3
C0023440|T191|PM|D004915|MSH|Leukemias, Acute Erythroblastic|9840/3
C0023440|T191|DSV|D004915|MSH|MYELOID LEUKEMIA ACUTE M 06|9840/3
C0023440|T191|ET|D004915|MSH|Myeloid Leukemia, Acute, M6|9840/3
C0023440|T191|PM|D004915|MSH|Myeloses, Erythremic|9840/3
C0023440|T191|PM|D004915|MSH|Myelosis, Erythremic|9840/3
C0023440|T191|PN|NOCODE|MTH|Acute Erythroblastic Leukemia|9840/3
C0023440|T191|ET|207.0|MTHICD9|Acute erythremic myelosis|9840/3
C0023440|T191|ET|207.0|MTHICD9|Di Guglielmo's disease|9840/3
C0023440|T191|ET|207.0|MTHICD9|Erythremic myelosis|9840/3
C0023440|T191|SY|C8923|NCI|Acute Erythroblastic Leukemia|9840/3
C0023440|T191|PT|C8923|NCI|Acute Erythroid Leukemia|9840/3
C0023440|T191|SY|TCGA|NCI|Acute Erythroid Leukemia|9840/3
C0023440|T191|AB|C8923|NCI|AEL|9840/3
C0023440|T191|PT|C95993|NCI|Di Guglielmo Syndrome|9840/3
C0023440|T191|SY|C8923|NCI|Erythroblastic Leukemia|9840/3
C0023440|T191|AB|C8923|NCI|FAB M6|9840/3
C0023440|T191|SY|C8923|NCI|M6 Acute Myeloid Leukemia|9840/3
C0023440|T191|SY|C8923|NCI_CDISC|Acute Erythroblastic Leukemia|9840/3
C0023440|T191|SY|C8923|NCI_CDISC|Erythroblastic Leukemia|9840/3
C0023440|T191|SY|C8923|NCI_CDISC|Fab M6|9840/3
C0023440|T191|PT|C8923|NCI_CDISC|LEUKEMIA, ERYTHROID, MALIGNANT|9840/3
C0023440|T191|SY|C8923|NCI_CDISC|M6 Acute Myeloid Leukemia|9840/3
C0023440|T191|PT|C8923|NCI_CPTAC|Acute Erythroid Leukemia|9840/3
C0023440|T191|PT|C8923|NCI_NICHD|Acute Erythroid Leukemia|9840/3
C0023440|T191|PT|R0121601|QMR|ERYTHROLEUKEMIA|9840/3
C0023440|T191|SY|XaBAl|RCD|Erythraemic myelosis|9840/3
C0023440|T191|PT|XaBAl|RCD|Erythroleukaemia|9840/3
C0023440|T191|SY|XaBAl|RCD|M6 - Acute erythroleukaemia|9840/3
C0023440|T191|PT|XaBAl|RCDAE|Erythroleukemia|9840/3
C0023440|T191|SY|XaBAl|RCDAE|M6 - Acute erythroleukemia|9840/3
C0023440|T191|PT|BBr40|RCDSA|Erythroleukemia|9840/3
C0023440|T191|OP|BBr4z|RCDSA|Erythroleukemia NOS|9840/3
C0023440|T191|PT|BBr40|RCDSY|Erythroleukaemia|9840/3
C0023440|T191|OP|BBr4z|RCDSY|Erythroleukaemia NOS|9840/3
C0023440|T191|OP|BBr4.|RCDSY|Erythroleukaemias|9840/3
C0023440|T191|IS|36449005|SNOMEDCT_US|Acute erythremic myelosis|9840/3
C0023440|T191|SYGB|14317002|SNOMEDCT_US|Acute erythroid leukaemia|9840/3
C0023440|T191|SY|14317002|SNOMEDCT_US|Acute erythroid leukemia|9840/3
C0023440|T191|PTGB|14317002|SNOMEDCT_US|Acute myeloid leukaemia, M6 type|9840/3
C0023440|T191|PT|14317002|SNOMEDCT_US|Acute myeloid leukemia, M6 type|9840/3
C0023440|T191|IS|14317002|SNOMEDCT_US|AML M6|9840/3
C0023440|T191|SY|93451002|SNOMEDCT_US|Di Guglielmo's disease|9840/3
C0023440|T191|IS|36449005|SNOMEDCT_US|Di Guglielmo's disease|9840/3
C0023440|T191|OAS|188752009|SNOMEDCT_US|Di Guglielmo's disease|9840/3
C0023440|T191|SYGB|93451002|SNOMEDCT_US|Erythraemic myelosis|9840/3
C0023440|T191|SYGB|14317002|SNOMEDCT_US|Erythraemic myelosis|9840/3
C0023440|T191|SY|93451002|SNOMEDCT_US|Erythremic myelosis|9840/3
C0023440|T191|SY|14317002|SNOMEDCT_US|Erythremic myelosis|9840/3
C0023440|T191|IS|14317002|SNOMEDCT_US|Erythremic myelosis, NOS|9840/3
C0023440|T191|SYGB|93451002|SNOMEDCT_US|Erythroleukaemia|9840/3
C0023440|T191|SYGB|14317002|SNOMEDCT_US|Erythroleukaemia|9840/3
C0023440|T191|PTGB|93451002|SNOMEDCT_US|Erythroleukaemia, FAB M6|9840/3
C0023440|T191|SY|93451002|SNOMEDCT_US|Erythroleukemia|9840/3
C0023440|T191|SY|14317002|SNOMEDCT_US|Erythroleukemia|9840/3
C0023440|T191|IS|93451002|SNOMEDCT_US|Erythroleukemia without mention of remission|9840/3
C0023440|T191|PT|93451002|SNOMEDCT_US|Erythroleukemia, FAB M6|9840/3
C0023440|T191|IS|14317002|SNOMEDCT_US|FAB M6|9840/3
C0023440|T191|SYGB|93451002|SNOMEDCT_US|M6 - Acute erythroleukaemia|9840/3
C0023440|T191|SY|93451002|SNOMEDCT_US|M6 - Acute erythroleukemia|9840/3
C0023440|T191|IS|14317002|SNOMEDCT_US|M6B|9840/3
C0023440|T191|IT|0565|WHO|DI GUGLIELMO'S SYNDROME|9840/3
C0023440|T191|IT|0565|WHO|ERYTHRAEMIC MYELOSIS|9840/3
C0023440|T191|PT|1132|WHO|ERYTHROLEUKEMIA|9840/3
C0023470|T191|NP|0000023091|AOD|myeloid leukemia|9860/3
C0206142|T191|SY|0000020820|CHV|eosinophil leukemia|9860/3
C0206142|T191|SY|0000020820|CHV|eosinophilic leukaemia|9860/3
C0206142|T191|PT|0000020820|CHV|eosinophilic leukemia|9860/3
C0206142|T191|SY|0000020820|CHV|eosinophils leukemia|9860/3
C0023470|T191|SY|0000007344|CHV|granulocytic leukaemia|9860/3
C0023470|T191|SY|0000007344|CHV|granulocytic leukemia|9860/3
C0023470|T191|SY|0000007344|CHV|leukaemia myelogenous|9860/3
C0023470|T191|SY|0000007344|CHV|leukemia myelocytic|9860/3
C0023470|T191|SY|0000007344|CHV|leukemia myelogenous|9860/3
C0023470|T191|SY|0000007344|CHV|leukemia myeloid|9860/3
C0023470|T191|SY|0000007344|CHV|myelocytic leukaemia|9860/3
C0023470|T191|SY|0000007344|CHV|myelocytic leukemia|9860/3
C0023470|T191|SY|0000007344|CHV|myelogenous leukaemia|9860/3
C0023470|T191|SY|0000007344|CHV|myelogenous leukemia|9860/3
C0023470|T191|SY|0000007344|CHV|myeloid leukaemia|9860/3
C0023470|T191|SY|0000007344|CHV|myeloid leukemia|9860/3
C0023470|T191|SY|0000007344|CHV|myelosis|9860/3
C0023470|T191|PT|NOCODE|COSTAR|Granulocytic Leukemia|9860/3
C0023470|T191|PT|NOCODE|COSTAR|Myelocytic Leukemia|9860/3
C0023470|T191|ET|2004-4431|CSP|granulocytic leukemia|9860/3
C0023470|T191|ET|2004-4431|CSP|myelocytic leukemia|9860/3
C0023470|T191|PT|2004-4431|CSP|myelogenous leukemia|9860/3
C0023470|T191|ET|2004-4431|CSP|myeloid granulocytic leukemia|9860/3
C0023470|T191|ET|2004-4431|CSP|myeloid leukemia|9860/3
C0023470|T191|ET|2004-4431|CSP|myelosis|9860/3
C0023470|T191|GT|LEUKEMIA CHRON MYELO|CST|LEUKAEMIA GRANULOCYTIC|9860/3
C0206142|T191|GT|LEUKEMIA CHRON MYELO|CST|LEUKEMIA EOSINOPHILIC|9860/3
C0023470|T191|GT|LEUKEMIA CHRON MYELO|CST|LEUKEMIA GRANULOCYTIC|9860/3
C0023470|T191|GT|LEUKEMIA CHRON MYELO|CST|LEUKEMIA MYELOGENOUS|9860/3
C0023470|T191|GT|LEUKEMIA CHRON MYELO|CST|LEUKEMIA MYELOID|9860/3
C0206142|T191|DI|U001046|DXP|LEUKEMIA, EOSINOPHILIC|9860/3
C0023470|T191|PT|HP:0012324|HPO|Myeloid leukemia|9860/3
C0023470|T191|HT|C92|ICD10|Myeloid leukaemia|9860/3
C0023470|T191|PT|C92.9|ICD10|Myeloid leukaemia, unspecified|9860/3
C0023470|T191|HT|C92|ICD10AE|Myeloid leukemia|9860/3
C0023470|T191|PT|C92.9|ICD10AE|Myeloid leukemia, unspecified|9860/3
C0023470|T191|ET|C92|ICD10CM|granulocytic leukemia|9860/3
C0023470|T191|ET|C92|ICD10CM|myelogenous leukemia|9860/3
C0023470|T191|AB|C92|ICD10CM|Myeloid leukemia|9860/3
C0023470|T191|HT|C92|ICD10CM|Myeloid leukemia|9860/3
C0023470|T191|AB|C92.9|ICD10CM|Myeloid leukemia, unspecified|9860/3
C0023470|T191|HT|C92.9|ICD10CM|Myeloid leukemia, unspecified|9860/3
C0023470|T191|ET|C92.90|ICD10CM|Myeloid leukemia, unspecified NOS|9860/3
C0023470|T191|HT|205|ICD9CM|Myeloid leukemia|9860/3
C0023470|T191|HT|205.9|ICD9CM|Unspecified myeloid leukemia|9860/3
C0206142|T191|PT|MTHU026442|ICPC2ICD10ENG|eosinophilic; leukemia|9860/3
C0023470|T191|PT|MTHU032693|ICPC2ICD10ENG|granulocytic; leukemia|9860/3
C0206142|T191|PT|MTHU044751|ICPC2ICD10ENG|leukemia; eosinophilic|9860/3
C0023470|T191|PT|MTHU044753|ICPC2ICD10ENG|leukemia; granulocytic|9860/3
C0023470|T191|PT|MTHU044780|ICPC2ICD10ENG|leukemia; myelocytic|9860/3
C0023470|T191|PT|MTHU044783|ICPC2ICD10ENG|leukemia; myeloid|9860/3
C0023470|T191|PT|MTHU050841|ICPC2ICD10ENG|myelocytic; leukemia|9860/3
C0023470|T191|PT|MTHU050854|ICPC2ICD10ENG|myeloid; leukemia|9860/3
C0023470|T191|PT|sh85089219|LCH_NW|Myeloid leukemia|9860/3
C0206142|T191|LLT|10014947|MDR|Eosinophil leukaemia|9860/3
C0206142|T191|LLT|10054374|MDR|Eosinophil leukemia|9860/3
C0206142|T191|PT|10014958|MDR|Eosinophilic leukaemia|9860/3
C0206142|T191|LLT|10014958|MDR|Eosinophilic leukaemia|9860/3
C0206142|T191|LLT|10014959|MDR|Eosinophilic leukemia|9860/3
C0206142|T191|MTH_PT|10014958|MDR|Eosinophilic leukemia|9860/3
C0206142|T191|LLT|10060389|MDR|Leukaemia eosinophilic|9860/3
C0023470|T191|LLT|10024299|MDR|Leukaemia granulocytic|9860/3
C0023470|T191|PT|10024299|MDR|Leukaemia granulocytic|9860/3
C0023470|T191|LLT|10024300|MDR|Leukaemia granulocytic NOS|9860/3
C0023470|T191|LLT|10024307|MDR|Leukaemia myelogenous|9860/3
C0023470|T191|LLT|10024308|MDR|Leukaemia myeloid|9860/3
C0206142|T191|LLT|10024334|MDR|Leukemia eosinophilic|9860/3
C0023470|T191|LLT|10024335|MDR|Leukemia granulocytic|9860/3
C0023470|T191|MTH_PT|10024299|MDR|Leukemia granulocytic|9860/3
C0023470|T191|LLT|10024336|MDR|Leukemia granulocytic NOS|9860/3
C0023470|T191|LLT|10024348|MDR|Leukemia myelogenous|9860/3
C0023470|T191|LLT|10024349|MDR|Leukemia myeloid|9860/3
C0023470|T191|OL|10024360|MDR|Leukemic granulocytic|9860/3
C0023470|T191|LLT|10028530|MDR|Myelocytic leukaemia|9860/3
C0023470|T191|LLT|10028531|MDR|Myelocytic leukemia|9860/3
C0023470|T191|PT|10028549|MDR|Myeloid leukaemia|9860/3
C0023470|T191|LLT|10028549|MDR|Myeloid leukaemia|9860/3
C0023470|T191|LLT|10028550|MDR|Myeloid leukaemia NOS|9860/3
C0023470|T191|MTH_PT|10028549|MDR|Myeloid leukemia|9860/3
C0023470|T191|LLT|10028555|MDR|Myeloid leukemia|9860/3
C0023470|T191|LLT|10028556|MDR|Myeloid leukemia NOS|9860/3
C0023470|T191|LLT|10029550|MDR|Non-lymphoblastic leukaemia NOS|9860/3
C0023470|T191|LLT|10029552|MDR|Non-lymphoblastic leukemia NOS|9860/3
C0023470|T191|LLT|10046039|MDR|Unspecified myeloid leukaemia|9860/3
C0023470|T191|LLT|10046040|MDR|Unspecified myeloid leukemia|9860/3
C0206142|T191|PT|31482|MEDCIN|eosinophilic leukemia|9860/3
C0206142|T191|SY|31482|MEDCIN|leukemia eosinophilic|9860/3
C0023470|T191|SY|99751|MEDCIN|leukemia myelogenous|9860/3
C0023470|T191|PT|99751|MEDCIN|myelogenous leukemia|9860/3
C0206142|T191|PM|D017681|MSH|Eosinophilic Leukemia|9860/3
C0206142|T191|PM|D017681|MSH|Eosinophilic Leukemias|9860/3
C0023470|T191|ET|D007951|MSH|Granulocytic Leukemia|9860/3
C0023470|T191|PM|D007951|MSH|Granulocytic Leukemias|9860/3
C0206142|T191|PEP|D017681|MSH|Leukemia, Eosinophilic|9860/3
C0023470|T191|ET|D007951|MSH|Leukemia, Granulocytic|9860/3
C0023470|T191|ET|D007951|MSH|Leukemia, Myelocytic|9860/3
C0023470|T191|ET|D007951|MSH|Leukemia, Myelogenous|9860/3
C0023470|T191|MH|D007951|MSH|Leukemia, Myeloid|9860/3
C0206142|T191|PM|D017681|MSH|Leukemias, Eosinophilic|9860/3
C0023470|T191|PM|D007951|MSH|Leukemias, Granulocytic|9860/3
C0023470|T191|PM|D007951|MSH|Leukemias, Myelocytic|9860/3
C0023470|T191|PM|D007951|MSH|Leukemias, Myelogenous|9860/3
C0023470|T191|PM|D007951|MSH|Leukemias, Myeloid|9860/3
C0023470|T191|ET|D007951|MSH|Myelocytic Leukemia|9860/3
C0023470|T191|PM|D007951|MSH|Myelocytic Leukemias|9860/3
C0023470|T191|ET|D007951|MSH|Myelogenous Leukemia|9860/3
C0023470|T191|PM|D007951|MSH|Myelogenous Leukemias|9860/3
C0023470|T191|ET|D007951|MSH|Myeloid Leukemia|9860/3
C0023470|T191|PM|D007951|MSH|Myeloid Leukemias|9860/3
C0206142|T191|PN|NOCODE|MTH|Eosinophilic leukemia|9860/3
C0023470|T191|SY|NOCODE|MTH|LEUKEMIA GRANULOCYTIC|9860/3
C0023470|T191|SY|NOCODE|MTH|LEUKEMIA MYELOGENOUS|9860/3
C0023470|T191|SY|NOCODE|MTH|LEUKEMIA MYELOID|9860/3
C0023470|T191|PN|NOCODE|MTH|Myeloid Leukemia|9860/3
C0206142|T191|ET|205.1|MTHICD9|Eosinophilic leukemia|9860/3
C0023470|T191|SY|C3172|NCI|Myelocytic Leukemia|9860/3
C0023470|T191|SY|C3172|NCI|Myelogenous Leukemia|9860/3
C0023470|T191|PT|C3172|NCI|Myeloid Leukemia|9860/3
C0023470|T191|OP|C3172|NCI|Non-Lymphoblastic Leukemia|9860/3
C0023470|T191|OP|C3172|NCI|Non-Lymphocytic Leukemia|9860/3
C0023470|T191|SY|C3172|NCI_CDISC|Leukemia Granulocytic|9860/3
C0023470|T191|SY|C3172|NCI_CDISC|Leukemia Myeloid|9860/3
C0023470|T191|PT|C3172|NCI_CDISC|LEUKEMIA, GRANULOCYTIC, MALIGNANT|9860/3
C0023470|T191|SY|C3172|NCI_CDISC|Myelocytic Leukemia|9860/3
C0023470|T191|SY|C3172|NCI_CDISC|Myelogenous Leukemia|9860/3
C0023470|T191|SY|C3172|NCI_CDISC|Non-lymphoblastic Leukemia|9860/3
C0023470|T191|SY|C3172|NCI_CDISC|Non-lymphocytic Leukemia|9860/3
C0023470|T191|PT|C3172|NCI_CPTAC|Myeloid Leukemia|9860/3
C0023470|T191|DN|C3172|NCI_CTRP|Myeloid Leukemia|9860/3
C0023470|T191|PT|C3172|NCI_CTRP|Myeloid Leukemia|9860/3
C0206142|T191|SY|CDR0000276487|PDQ|Eosinophilic Leukemia|9860/3
C0206142|T191|PT|BBr80|RCD|Eosinophilic leukaemia|9860/3
C0023470|T191|SY|B65..|RCD|Granulocytic leukaemia|9860/3
C0023470|T191|PT|B65..|RCD|Myeloid leukaemia|9860/3
C0023470|T191|OP|B65z.|RCD|Myeloid leukaemia NOS|9860/3
C0206142|T191|PT|BBr80|RCDAE|Eosinophilic leukemia|9860/3
C0023470|T191|SY|B65..|RCDAE|Granulocytic leukemia|9860/3
C0023470|T191|PT|B65..|RCDAE|Myeloid leukemia|9860/3
C0023470|T191|OP|B65z.|RCDAE|Myeloid leukemia NOS|9860/3
C0206142|T191|OP|BBr8z|RCDSA|Eosinophilic leukemia NOS|9860/3
C0206142|T191|OP|BBr8.|RCDSA|Eosinophilic leukemias|9860/3
C0023470|T191|OP|BBr60|RCDSA|Myeloid leukemia NOS|9860/3
C0023470|T191|PT|BBr6.|RCDSA|Myeloid leukemias|9860/3
C0206142|T191|OP|BBr8z|RCDSY|Eosinophilic leukaemia NOS|9860/3
C0206142|T191|OP|BBr8.|RCDSY|Eosinophilic leukaemias|9860/3
C0023470|T191|OP|BBr60|RCDSY|Myeloid leukaemia NOS|9860/3
C0023470|T191|PT|BBr6.|RCDSY|Myeloid leukaemias|9860/3
C0206142|T191|OAP|57147001|SNOMEDCT_US|Eosinophilic leukaemia|9860/3
C0206142|T191|PTGB|190055003|SNOMEDCT_US|Eosinophilic leukaemia|9860/3
C0206142|T191|SYGB|37810007|SNOMEDCT_US|Eosinophilic leukaemia|9860/3
C0206142|T191|IS|57147001|SNOMEDCT_US|Eosinophilic leukaemia -RETIRED-|9860/3
C0206142|T191|PT|190055003|SNOMEDCT_US|Eosinophilic leukemia|9860/3
C0206142|T191|SY|37810007|SNOMEDCT_US|Eosinophilic leukemia|9860/3
C0206142|T191|OAP|57147001|SNOMEDCT_US|Eosinophilic leukemia|9860/3
C0206142|T191|IS|57147001|SNOMEDCT_US|Eosinophilic leukemia -RETIRED-|9860/3
C0206142|T191|OF|57147001|SNOMEDCT_US|Eosinophilic leukemia -RETIRED-|9860/3
C0023470|T191|SYGB|37810007|SNOMEDCT_US|Granulocytic leukaemia|9860/3
C0023470|T191|SYGB|188732008|SNOMEDCT_US|Granulocytic leukaemia|9860/3
C0023470|T191|SY|37810007|SNOMEDCT_US|Granulocytic leukemia|9860/3
C0023470|T191|SY|188732008|SNOMEDCT_US|Granulocytic leukemia|9860/3
C0023470|T191|IS|37810007|SNOMEDCT_US|Granulocytic leukemia, NOS|9860/3
C0023470|T191|SYGB|37810007|SNOMEDCT_US|Myelocytic leukaemia|9860/3
C0023470|T191|SY|37810007|SNOMEDCT_US|Myelocytic leukemia|9860/3
C0023470|T191|IS|37810007|SNOMEDCT_US|Myelocytic leukemia, NOS|9860/3
C0023470|T191|SYGB|37810007|SNOMEDCT_US|Myelogenous leukaemia|9860/3
C0023470|T191|SY|37810007|SNOMEDCT_US|Myelogenous leukemia|9860/3
C0023470|T191|IS|37810007|SNOMEDCT_US|Myelogenous leukemia, NOS|9860/3
C0023470|T191|OAS|154587007|SNOMEDCT_US|Myeloid leukaemia|9860/3
C0023470|T191|OAS|269631008|SNOMEDCT_US|Myeloid leukaemia|9860/3
C0023470|T191|PTGB|37810007|SNOMEDCT_US|Myeloid leukaemia|9860/3
C0023470|T191|PTGB|188732008|SNOMEDCT_US|Myeloid leukaemia|9860/3
C0023470|T191|OAP|94717009|SNOMEDCT_US|Myeloid leukaemia|9860/3
C0023470|T191|OAP|324170002|SNOMEDCT_US|Myeloid leukaemia|9860/3
C0023470|T191|SYGB|128934006|SNOMEDCT_US|Myeloid leukaemia - category|9860/3
C0023470|T191|OAP|188743000|SNOMEDCT_US|Myeloid leukaemia NOS|9860/3
C0023470|T191|IS|37810007|SNOMEDCT_US|Myeloid leukaemia, NOS|9860/3
C0023470|T191|OAP|94717009|SNOMEDCT_US|Myeloid leukemia|9860/3
C0023470|T191|OAP|324170002|SNOMEDCT_US|Myeloid leukemia|9860/3
C0023470|T191|OAS|269631008|SNOMEDCT_US|Myeloid leukemia|9860/3
C0023470|T191|OAS|154587007|SNOMEDCT_US|Myeloid leukemia|9860/3
C0023470|T191|PT|37810007|SNOMEDCT_US|Myeloid leukemia|9860/3
C0023470|T191|PT|188732008|SNOMEDCT_US|Myeloid leukemia|9860/3
C0023470|T191|SY|128934006|SNOMEDCT_US|Myeloid leukemia - category|9860/3
C0023470|T191|OAP|188743000|SNOMEDCT_US|Myeloid leukemia NOS|9860/3
C0023470|T191|SY|37810007|SNOMEDCT_US|Myeloid leukemia, no International Classification of Diseases for Oncology subtype|9860/3
C0023470|T191|IS|37810007|SNOMEDCT_US|Myeloid leukemia, NOS|9860/3
C0023470|T191|SYGB|37810007|SNOMEDCT_US|Non-lymphocytic leukaemia|9860/3
C0023470|T191|SY|37810007|SNOMEDCT_US|Non-lymphocytic leukemia|9860/3
C0023470|T191|PT|0575|WHO|LEUKAEMIA GRANULOCYTIC|9860/3
C0023470|T191|IT|0575|WHO|LEUKAEMIA MYELOGENOUS|9860/3
C0023470|T191|IT|0575|WHO|LEUKAEMIA MYELOID|9860/3
C0023467|T191|PT|BI00289|BI|acute myelogenous leukemia|9861/3
C0023467|T191|AB|BI00289|BI|aml|9861/3
C0023467|T191|PT|0062086|CCPSS|LEUKEMIA ACUTE MYELOGENOUS|9861/3
C0023467|T191|SY|0000007343|CHV|acute granulocytic leukemia|9861/3
C0023467|T191|SY|0000050375|CHV|acute leukemias non lymphoblastic|9861/3
C0023467|T191|SY|0000007343|CHV|acute myeloblastic leukemia|9861/3
C0023467|T191|SY|0000007343|CHV|acute myelocytic leukaemia|9861/3
C0023467|T191|SY|0000007343|CHV|acute myelocytic leukemia|9861/3
C0023467|T191|SY|0000007343|CHV|acute myelogenous leukaemia|9861/3
C0023467|T191|SY|0000007343|CHV|acute myelogenous leukemia|9861/3
C0023467|T191|SY|0000007343|CHV|acute myeloid leukaemia|9861/3
C0023467|T191|SY|0000007343|CHV|acute myeloid leukemia|9861/3
C0023467|T191|SY|0000007343|CHV|acute myeloid leukemias|9861/3
C0023467|T191|SY|0000050375|CHV|acute non-lymphoblastic leukemia|9861/3
C0023467|T191|SY|0000007343|CHV|acute non-lymphocytic leukemia|9861/3
C0023467|T191|SY|0000007348|CHV|acute nonlymphoblastic leukemia|9861/3
C0023467|T191|SY|0000007348|CHV|acute nonlymphocytic leukemia|9861/3
C0023467|T191|SY|0000007343|CHV|aml|9861/3
C0023467|T191|SY|0000007348|CHV|anll|9861/3
C0023467|T191|PT|0000050375|CHV|non-lymphoblastic leukemia acute|9861/3
C0023467|T191|PT|025|COSTAR|ACUTE MYELOGENOUS LEUKEMIA|9861/3
C0023467|T191|ET|4000-0108|CSP|acute granulocytic leukemia|9861/3
C0023467|T191|ET|4000-0108|CSP|acute myeloblastic leukemia|9861/3
C0023467|T191|ET|4000-0108|CSP|acute myelocytic leukemia|9861/3
C0023467|T191|PT|4000-0108|CSP|acute myelogenous leukemia|9861/3
C0023467|T191|ET|4000-0108|CSP|acute myeloid leukemia|9861/3
C0023467|T191|PT|4001-0002|CSP|acute nonlymphocytic leukemia|9861/3
C0023467|T191|ET|4000-0108|CSP|AML|9861/3
C0023467|T191|ET|4001-0002|CSP|ANLL|9861/3
C0023467|T191|PT|LEUKEMIA ACUTE MYELO|CST|ACUTE MYELOBLASTIC LEUKEMIA|9861/3
C0023467|T191|GT|LEUKEMIA ACUTE MYELO|CST|LEUKEMIA MYELOBLASTIC ACUTE|9861/3
C0023467|T191|SY|NOCODE|DXP|AML|9861/3
C0023467|T191|SY|NOCODE|DXP|LEUKEMIA, GRANULOCYTIC, ACUTE|9861/3
C0023467|T191|DI|U001051|DXP|LEUKEMIA, MYELOBLASTIC, ACUTE|9861/3
C0023467|T191|SY|NOCODE|DXP|LEUKEMIA, MYELOCYTIC, ACUTE|9861/3
C0023467|T191|SY|NOCODE|DXP|LEUKEMIA, MYELOGENOUS, ACUTE|9861/3
C0023467|T191|SY|NOCODE|DXP|LEUKEMIA, MYELOID, ACUTE|9861/3
C0023467|T191|SY|HP:0004808|HPO|Acute myeloblastic leukemia|9861/3
C0023467|T191|SY|HP:0004808|HPO|Acute myelocytic leukemia|9861/3
C0023467|T191|SY|HP:0004808|HPO|Acute myelogenous leukemia|9861/3
C0023467|T191|PT|HP:0004808|HPO|Acute myeloid leukemia|9861/3
C0023467|T191|SY|HP:0004808|HPO|AML|9861/3
C0023467|T191|PT|C92.0|ICD10|Acute myeloid leukaemia|9861/3
C0023467|T191|PT|C92.0|ICD10AE|Acute myeloid leukemia|9861/3
C0023467|T191|AB|C92.0|ICD10CM|Acute myeloblastic leukemia|9861/3
C0023467|T191|HT|C92.0|ICD10CM|Acute myeloblastic leukemia|9861/3
C0023467|T191|ET|C92.00|ICD10CM|Acute myeloblastic leukemia NOS|9861/3
C0023467|T191|HT|205.0|ICD9CM|Myeloid leukemia, acute|9861/3
C0023467|T191|PT|MTHU032694|ICPC2ICD10ENG|granulocytic; leukemia, acute|9861/3
C0023467|T191|PT|MTHU044754|ICPC2ICD10ENG|leukemia; granulocytic, acute|9861/3
C0023467|T191|PT|MTHU044781|ICPC2ICD10ENG|leukemia; myelocytic, acute|9861/3
C0023467|T191|PT|MTHU044784|ICPC2ICD10ENG|leukemia; myeloid, acute|9861/3
C0023467|T191|PT|MTHU050842|ICPC2ICD10ENG|myelocytic; leukemia, acute|9861/3
C0023467|T191|PT|MTHU050855|ICPC2ICD10ENG|myeloid; leukemia, acute|9861/3
C0023467|T191|PTN|B73002|ICPC2P|acute myeloid leukaemia|9861/3
C0023467|T191|MTH_PTN|B73002|ICPC2P|acute myeloid leukemia|9861/3
C0023467|T191|PT|B73002|ICPC2P|Leukaemia;acute myeloid|9861/3
C0023467|T191|MTH_PT|B73002|ICPC2P|Leukemia;acute myeloid|9861/3
C0023467|T191|PT|sh90001715|LCH_NW|Acute myeloid leukemia|9861/3
C0023467|T191|LA|LA26787-4|LNC|Acute myeloid leukemia|9861/3
C0023467|T191|LLT|10000801|MDR|Acute granulocytic leukaemia|9861/3
C0023467|T191|LLT|10060553|MDR|Acute granulocytic leukemia|9861/3
C0023467|T191|LLT|10060354|MDR|Acute myeloblastic leukaemia|9861/3
C0023467|T191|LLT|10000878|MDR|Acute myeloblastic leukemia|9861/3
C0023467|T191|LLT|10051003|MDR|Acute myelocytic leukaemia|9861/3
C0023467|T191|LLT|10060557|MDR|Acute myelocytic leukemia|9861/3
C0023467|T191|LLT|10000880|MDR|Acute myeloid leukaemia|9861/3
C0023467|T191|PT|10000880|MDR|Acute myeloid leukaemia|9861/3
C0023467|T191|LLT|10000884|MDR|Acute myeloid leukaemia NOS|9861/3
C0023467|T191|LLT|10000886|MDR|Acute myeloid leukemia|9861/3
C0023467|T191|MTH_PT|10000880|MDR|Acute myeloid leukemia|9861/3
C0023467|T191|LLT|10054296|MDR|Acute myeloid leukemia NOS|9861/3
C0023467|T191|OL|10001941|MDR|AML|9861/3
C0023467|T191|LLT|10060394|MDR|Leukaemia myeloblastic acute|9861/3
C0023467|T191|HT|10024291|MDR|Leukaemias acute myeloid|9861/3
C0023467|T191|LLT|10024346|MDR|Leukemia myeloblastic acute|9861/3
C0023467|T191|MTH_HT|10024291|MDR|Leukemias acute myeloid|9861/3
C0023467|T191|LLT|10028552|MDR|Myeloid leukaemia, acute|9861/3
C0023467|T191|LLT|10028557|MDR|Myeloid leukemia, acute|9861/3
C0023467|T191|LLT|10029549|MDR|Non-lymphoblastic leukaemia acute|9861/3
C0023467|T191|LLT|10029551|MDR|Non-lymphoblastic leukemia acute|9861/3
C0023467|T191|PT|338565|MEDCIN|acute myeloblastic leukemia|9861/3
C0023467|T191|PT|31476|MEDCIN|acute myelogenous leukemia|9861/3
C0023467|T191|SY|338565|MEDCIN|leukemia acute myeloblastic|9861/3
C0023467|T191|ET|5622|MEDLINEPLUS|Acute Myeloblastic Leukemia|9861/3
C0023467|T191|SY|5622|MEDLINEPLUS|Acute myelogenous leukemia|9861/3
C0023467|T191|PT|5622|MEDLINEPLUS|Acute Myeloid Leukemia|9861/3
C0023467|T191|SY|5622|MEDLINEPLUS|AML|9861/3
C0023467|T191|ET|5622|MEDLINEPLUS|AML|9861/3
C0023467|T191|SY|5622|MEDLINEPLUS|ANLL|9861/3
C0023467|T191|ET|5622|MEDLINEPLUS|Leukemia, Myeloblastic, Acute|9861/3
C0023467|T191|ET|5622|MEDLINEPLUS|Leukemia, Myelogenous, Acute|9861/3
C0023467|T191|ET|5622|MEDLINEPLUS|Leukemia, Myeloid, Acute|9861/3
C0023467|T191|PM|D015470|MSH|Acute Myeloblastic Leukemia|9861/3
C0023467|T191|PM|D015470|MSH|Acute Myeloblastic Leukemias|9861/3
C0023467|T191|PM|D015470|MSH|Acute Myelocytic Leukemia|9861/3
C0023467|T191|PM|D015470|MSH|Acute Myelocytic Leukemias|9861/3
C0023467|T191|ET|D015470|MSH|Acute Myelogenous Leukemia|9861/3
C0023467|T191|PM|D015470|MSH|Acute Myelogenous Leukemias|9861/3
C0023467|T191|ET|D015470|MSH|Acute Myeloid Leukemia|9861/3
C0023467|T191|PM|D015470|MSH|Acute Myeloid Leukemias|9861/3
C0023467|T191|PM|D015470|MSH|Acute Nonlymphoblastic Leukemia|9861/3
C0023467|T191|PM|D015470|MSH|Acute Nonlymphoblastic Leukemias|9861/3
C0023467|T191|PM|D015470|MSH|Acute Nonlymphocytic Leukemia|9861/3
C0023467|T191|PM|D015470|MSH|Acute Nonlymphocytic Leukemias|9861/3
C0023467|T191|ET|D015470|MSH|ANLL|9861/3
C0023467|T191|PM|D015470|MSH|Leukemia, Acute Myeloblastic|9861/3
C0023467|T191|PM|D015470|MSH|Leukemia, Acute Myelocytic|9861/3
C0023467|T191|ET|D015470|MSH|Leukemia, Acute Myelogenous|9861/3
C0023467|T191|ET|D015470|MSH|Leukemia, Acute Myeloid|9861/3
C0023467|T191|PM|D015470|MSH|Leukemia, Acute Nonlymphoblastic|9861/3
C0023467|T191|PM|D015470|MSH|Leukemia, Acute Nonlymphocytic|9861/3
C0023467|T191|ET|D015470|MSH|Leukemia, Myeloblastic, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Leukemia, Myelocytic, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Leukemia, Myelogenous, Acute|9861/3
C0023467|T191|MH|D015470|MSH|Leukemia, Myeloid, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Leukemia, Nonlymphoblastic, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Leukemia, Nonlymphocytic, Acute|9861/3
C0023467|T191|PM|D015470|MSH|Leukemias, Acute Myeloblastic|9861/3
C0023467|T191|PM|D015470|MSH|Leukemias, Acute Myelocytic|9861/3
C0023467|T191|PM|D015470|MSH|Leukemias, Acute Myelogenous|9861/3
C0023467|T191|PM|D015470|MSH|Leukemias, Acute Myeloid|9861/3
C0023467|T191|PM|D015470|MSH|Leukemias, Acute Nonlymphoblastic|9861/3
C0023467|T191|PM|D015470|MSH|Leukemias, Acute Nonlymphocytic|9861/3
C0023467|T191|ET|D015470|MSH|Myeloblastic Leukemia, Acute|9861/3
C0023467|T191|PM|D015470|MSH|Myeloblastic Leukemias, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Myelocytic Leukemia, Acute|9861/3
C0023467|T191|PM|D015470|MSH|Myelocytic Leukemias, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Myelogenous Leukemia, Acute|9861/3
C0023467|T191|PM|D015470|MSH|Myelogenous Leukemias, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Myeloid Leukemia, Acute|9861/3
C0023467|T191|PM|D015470|MSH|Myeloid Leukemias, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Nonlymphoblastic Leukemia, Acute|9861/3
C0023467|T191|PM|D015470|MSH|Nonlymphoblastic Leukemias, Acute|9861/3
C0023467|T191|ET|D015470|MSH|Nonlymphocytic Leukemia, Acute|9861/3
C0023467|T191|PM|D015470|MSH|Nonlymphocytic Leukemias, Acute|9861/3
C0023467|T191|PN|NOCODE|MTH|Leukemia, Myelocytic, Acute|9861/3
C0023467|T191|SY|C3171|NCI|Acute Myeloblastic Leukemia|9861/3
C0023467|T191|OP|C3171|NCI|Acute Myelocytic Leukemia|9861/3
C0023467|T191|SY|C3171|NCI|Acute Myelogenous Leukemia|9861/3
C0023467|T191|SY|C3171|NCI|Acute Myelogenous Leukemias|9861/3
C0023467|T191|PT|C3171|NCI|Acute Myeloid Leukemia|9861/3
C0023467|T191|SY|TCGA|NCI|Acute Myeloid Leukemia|9861/3
C0023467|T191|SY|C27753|NCI|Acute Myeloid Leukemia NOS|9861/3
C0023467|T191|SY|C27753|NCI|Acute Myeloid Leukemia Not Otherwise Categorized|9861/3
C0023467|T191|PT|C27753|NCI|Acute Myeloid Leukemia Not Otherwise Specified|9861/3
C0023467|T191|SY|TCGA|NCI|Acute Myeloid Leukemia Not Otherwise Specified|9861/3
C1275661|T191|SY|C7175|NCI|Acute Myeloid Leukemia with Balanced Translocations/Inversions|9861/3
C4329268|T191|PT|C129785|NCI|Acute Myeloid Leukemia with BCR-ABL1|9861/3
C2826177|T191|SY|C82431|NCI|Acute Myeloid Leukemia with Cytoplasmic Nucleophosmin|9861/3
C2826178|T191|PT|C82433|NCI|Acute Myeloid Leukemia with Mutated CEBPA|9861/3
C2826178|T191|SY|TCGA|NCI|Acute Myeloid Leukemia with Mutated CEBPA|9861/3
C2826177|T191|PT|C82431|NCI|Acute Myeloid Leukemia with Mutated NPM1|9861/3
C2826177|T191|SY|TCGA|NCI|Acute Myeloid Leukemia with Mutated NPM1|9861/3
C4329271|T191|PT|C129786|NCI|Acute Myeloid Leukemia with Mutated RUNX1|9861/3
C2826178|T191|SY|C82433|NCI|Acute Myeloid Leukemia with Non-Germline Mutated CEBPA|9861/3
C4329271|T191|SY|C129786|NCI|Acute Myeloid Leukemia with Non-Germline Mutated RUNX1|9861/3
C1275661|T191|PT|C7175|NCI|Acute Myeloid Leukemia with Recurrent Genetic Abnormalities|9861/3
C1275661|T191|SY|TCGA|NCI|Acute Myeloid Leukemia with Recurrent Genetic Abnormalities|9861/3
C0023467|T191|SY|C27753|NCI|Acute Myeloid Leukemia, NOS|9861/3
C0023467|T191|OP|C3171|NCI|Acute Nonlymphocytic Leukemia|9861/3
C0023467|T191|AB|C3171|NCI|AML|9861/3
C0023467|T191|SY|C3171|NCI|AML - Acute Myeloid Leukemia|9861/3
C2826178|T191|SY|C82433|NCI|AML with Mutated CEBPA|9861/3
C2826177|T191|SY|C82431|NCI|AML with Mutated NPM1|9861/3
C0023467|T191|AB|C27753|NCI|AML, NOS|9861/3
C0023467|T191|AB|C3171|NCI|ANLL|9861/3
C2826178|T191|SY|C82433|NCI|Non-Familial Acute Myeloid Leukemia with Mutated CEBPA|9861/3
C2826177|T191|AB|C82431|NCI|NPMc+ AML|9861/3
C0023467|T191|PT|C3171|NCI_CPTAC|Acute Myeloid Leukemia|9861/3
C0023467|T191|SY|10000884|NCI_CTEP-SDC|Acute myeloid leukemia|9861/3
C0023467|T191|PT|10000884|NCI_CTEP-SDC|Acute myeloid leukemia, NOS|9861/3
C0023467|T191|SY|C3171|NCI_CTRP|Acute Myeloid Leukemia|9861/3
C0023467|T191|SY|CDR0000575435|NCI_NCI-GLOSS|acute myeloblastic leukemia|9861/3
C0023467|T191|PT|CDR0000046757|NCI_NCI-GLOSS|acute myelogenous leukemia|9861/3
C0023467|T191|PT|CDR0000046347|NCI_NCI-GLOSS|acute myeloid leukemia|9861/3
C0023467|T191|PT|CDR0000046215|NCI_NCI-GLOSS|acute nonlymphocytic leukemia|9861/3
C0023467|T191|PT|CDR0000044363|NCI_NCI-GLOSS|AML|9861/3
C0023467|T191|SY|CDR0000575436|NCI_NCI-GLOSS|ANLL|9861/3
C0023467|T191|SY|C3171|NCI_NICHD|Acute Granulocytic Leukemia|9861/3
C0023467|T191|SY|C3171|NCI_NICHD|Acute Myelocytic Leukemia|9861/3
C0023467|T191|SY|C3171|NCI_NICHD|Acute Myelogenous Leukemia|9861/3
C0023467|T191|PT|C3171|NCI_NICHD|Acute Myeloid Leukemia|9861/3
C2826178|T191|PT|C82433|NCI_NICHD|Acute Myeloid Leukemia with Mutated CEBPA|9861/3
C2826177|T191|PT|C82431|NCI_NICHD|Acute Myeloid Leukemia with Mutated NPM1|9861/3
C1275661|T191|PT|C7175|NCI_NICHD|Acute Myeloid Leukemia with Recurrent Genetic Abnormalities|9861/3
C0023467|T191|SY|C3171|NCI_NICHD|AML|9861/3
C2826178|T191|SY|C82433|NCI_NICHD|AML with Mutated CEBPA|9861/3
C2826177|T191|SY|C82431|NCI_NICHD|AML with Mutated NPM1|9861/3
C1275661|T191|SY|C7175|NCI_NICHD|AML with Recurrent Genetic Abnormalities|9861/3
C0023467|T191|SY|CDR0000043424|PDQ|acute myeloblastic leukemia|9861/3
C0023467|T191|IS|CDR0000043424|PDQ|acute myelocytic leukemia|9861/3
C0023467|T191|SY|CDR0000043424|PDQ|acute myelogenous leukemia|9861/3
C0023467|T191|SY|CDR0000043424|PDQ|acute myelogenous leukemias|9861/3
C0023467|T191|PT|CDR0000043424|PDQ|acute myeloid leukemia|9861/3
C0023467|T191|IS|CDR0000043424|PDQ|acute nonlymphocytic leukemia|9861/3
C0023467|T191|AB|CDR0000043424|PDQ|AML|9861/3
C0023467|T191|SY|CDR0000043424|PDQ|AML - Acute Myeloid Leukemia|9861/3
C0023467|T191|AB|CDR0000043424|PDQ|ANLL|9861/3
C0023467|T191|SY|CDR0000043424|PDQ|leukemia, acute myeloid|9861/3
C0023467|T191|SY|CDR0000043424|PDQ|leukemia, acute nonlymphocytic|9861/3
C0023467|T191|PT|R0121661|QMR|LEUKEMIA ACUTE MYELOBLASTIC|9861/3
C0023467|T191|PT|Xa0Sk|RCD|Acute myeloblastic leukaemia|9861/3
C0023467|T191|PT|B650.|RCD|Acute myeloid leukaemia|9861/3
C0023467|T191|AB|Xa0Sk|RCD|AML - Acute myelobl leukaemia|9861/3
C0023467|T191|SY|Xa0Sk|RCD|AML - Acute myeloblastic leukaemia|9861/3
C0023467|T191|SY|B650.|RCD|AML - Acute myeloid leukaemia|9861/3
C0023467|T191|PT|Xa0Sk|RCDAE|Acute myeloblastic leukemia|9861/3
C0023467|T191|PT|B650.|RCDAE|Acute myeloid leukemia|9861/3
C0023467|T191|AB|Xa0Sk|RCDAE|AML - Acute myelobl leukemia|9861/3
C0023467|T191|SY|Xa0Sk|RCDAE|AML - Acute myeloblastic leukemia|9861/3
C0023467|T191|SY|B650.|RCDAE|AML - Acute myeloid leukemia|9861/3
C0023467|T191|PT|BBr61|RCDSA|Acute myeloid leukemia|9861/3
C0023467|T191|PT|BBr61|RCDSY|Acute myeloid leukaemia|9861/3
C0023467|T191|SYGB|17788007|SNOMEDCT_US|Acute granulocytic leukaemia|9861/3
C0023467|T191|SY|17788007|SNOMEDCT_US|Acute granulocytic leukemia|9861/3
C0023467|T191|OAP|277600006|SNOMEDCT_US|Acute myeloblastic leukaemia|9861/3
C0023467|T191|SYGB|17788007|SNOMEDCT_US|Acute myeloblastic leukaemia|9861/3
C0023467|T191|OAP|277600006|SNOMEDCT_US|Acute myeloblastic leukemia|9861/3
C0023467|T191|SY|17788007|SNOMEDCT_US|Acute myeloblastic leukemia|9861/3
C0023467|T191|SYGB|91861009|SNOMEDCT_US|Acute myelocytic leukaemia|9861/3
C0023467|T191|SYGB|17788007|SNOMEDCT_US|Acute myelocytic leukaemia|9861/3
C0023467|T191|SY|91861009|SNOMEDCT_US|Acute myelocytic leukemia|9861/3
C0023467|T191|SY|17788007|SNOMEDCT_US|Acute myelocytic leukemia|9861/3
C0023467|T191|SYGB|17788007|SNOMEDCT_US|Acute myelogenous leukaemia|9861/3
C0023467|T191|SY|17788007|SNOMEDCT_US|Acute myelogenous leukemia|9861/3
C0023467|T191|PTGB|413443009|SNOMEDCT_US|Acute myeloid leukaemia|9861/3
C0023467|T191|OP|17788007|SNOMEDCT_US|Acute myeloid leukaemia|9861/3
C0023467|T191|SYGB|91861009|SNOMEDCT_US|Acute myeloid leukaemia|9861/3
C0023467|T191|SYGB|413443009|SNOMEDCT_US|Acute myeloid leukaemia - category|9861/3
C4329268|T191|PTGB|783017000|SNOMEDCT_US|Acute myeloid leukaemia with BCR-ABL1|9861/3
C4543165|T191|PTGB|734524001|SNOMEDCT_US|Acute myeloid leukaemia with FMS-like tyrosine kinase-3 mutation|9861/3
C4543165|T191|PTGB|734522002|SNOMEDCT_US|Acute myeloid leukaemia with FMS-like tyrosine kinase-3 mutation|9861/3
C4543165|T191|SYGB|734522002|SNOMEDCT_US|Acute myeloid leukaemia with FTL3 mutation|9861/3
C4543165|T191|SYGB|734524001|SNOMEDCT_US|Acute myeloid leukaemia with FTL3 mutation|9861/3
C2826178|T191|OP|703819004|SNOMEDCT_US|Acute myeloid leukaemia with mutated CEBPA|9861/3
C2826177|T191|PTGB|703820005|SNOMEDCT_US|Acute myeloid leukaemia with mutated NPM1|9861/3
C4329271|T191|PTGB|783263001|SNOMEDCT_US|Acute myeloid leukaemia with mutated RUNX1|9861/3
C2826178|T191|SYGB|703819004|SNOMEDCT_US|Acute myeloid leukaemia with mutation of CCAAT enhancer binding protein alpha gene|9861/3
C1275661|T191|PTGB|397340004|SNOMEDCT_US|Acute myeloid leukaemia with recurrent genetic abnormality|9861/3
C0023467|T191|PTGB|91861009|SNOMEDCT_US|Acute myeloid leukaemia, disease|9861/3
C0023467|T191|PTGB|17788007|SNOMEDCT_US|Acute myeloid leukaemia, no ICD-O subtype|9861/3
C0023467|T191|PT|413443009|SNOMEDCT_US|Acute myeloid leukemia|9861/3
C0023467|T191|SY|91861009|SNOMEDCT_US|Acute myeloid leukemia|9861/3
C0023467|T191|OP|17788007|SNOMEDCT_US|Acute myeloid leukemia|9861/3
C0023467|T191|SY|413443009|SNOMEDCT_US|Acute myeloid leukemia - category|9861/3
C4329268|T191|PT|783017000|SNOMEDCT_US|Acute myeloid leukemia with BCR-ABL1|9861/3
C4543165|T191|PT|734524001|SNOMEDCT_US|Acute myeloid leukemia with FMS-like tyrosine kinase-3 mutation|9861/3
C4543165|T191|PT|734522002|SNOMEDCT_US|Acute myeloid leukemia with FMS-like tyrosine kinase-3 mutation|9861/3
C4543165|T191|SY|734524001|SNOMEDCT_US|Acute myeloid leukemia with FTL3 mutation|9861/3
C4543165|T191|SY|734522002|SNOMEDCT_US|Acute myeloid leukemia with FTL3 mutation|9861/3
C2826178|T191|OP|703819004|SNOMEDCT_US|Acute myeloid leukemia with mutated CEBPA|9861/3
C2826177|T191|PT|703820005|SNOMEDCT_US|Acute myeloid leukemia with mutated NPM1|9861/3
C4329271|T191|PT|783263001|SNOMEDCT_US|Acute myeloid leukemia with mutated RUNX1|9861/3
C2826178|T191|SY|703819004|SNOMEDCT_US|Acute myeloid leukemia with mutation of CCAAT enhancer binding protein alpha gene|9861/3
C1275661|T191|PT|397340004|SNOMEDCT_US|Acute myeloid leukemia with recurrent genetic abnormality|9861/3
C0023467|T191|PT|91861009|SNOMEDCT_US|Acute myeloid leukemia, disease|9861/3
C0023467|T191|PT|17788007|SNOMEDCT_US|Acute myeloid leukemia, no ICD-O subtype|9861/3
C0023467|T191|SY|17788007|SNOMEDCT_US|Acute myeloid leukemia, no International Classification of Diseases for Oncology subtype|9861/3
C0023467|T191|SYGB|17788007|SNOMEDCT_US|Acute non-lymphocytic leukaemia|9861/3
C0023467|T191|SY|17788007|SNOMEDCT_US|Acute non-lymphocytic leukemia|9861/3
C0023467|T191|OAS|277600006|SNOMEDCT_US|AML - Acute myeloblastic leukaemia|9861/3
C0023467|T191|SYGB|91861009|SNOMEDCT_US|AML - Acute myeloblastic leukaemia|9861/3
C0023467|T191|OAS|277600006|SNOMEDCT_US|AML - Acute myeloblastic leukemia|9861/3
C0023467|T191|SY|91861009|SNOMEDCT_US|AML - Acute myeloblastic leukemia|9861/3
C0023467|T191|SYGB|91861009|SNOMEDCT_US|AML - Acute myeloid leukaemia|9861/3
C0023467|T191|SY|91861009|SNOMEDCT_US|AML - Acute myeloid leukemia|9861/3
C1275661|T191|SY|397340004|SNOMEDCT_US|AML with recurrent genetic abnormality|9861/3
C0023473|T191|PT|BI00304|BI|chronic myelogenous leukemia|9863/3
C0023473|T191|AB|BI00304|BI|cml|9863/3
C0023473|T191|PT|0003456|CCPSS|LEUKEMIA CHRONIC MYELOGENOUS|9863/3
C0023473|T191|SY|0000007345|CHV|chronic granulocytic leukaemia|9863/3
C0023473|T191|SY|0000007345|CHV|chronic granulocytic leukemia|9863/3
C0023473|T191|SY|0000007345|CHV|chronic myelocytic leukemia|9863/3
C0023473|T191|SY|0000007345|CHV|chronic myelogenous leukaemia|9863/3
C0023473|T191|SY|0000007345|CHV|chronic myelogenous leukemia|9863/3
C0023473|T191|SY|0000007345|CHV|chronic myeloid leukaemia|9863/3
C0023473|T191|SY|0000007345|CHV|chronic myeloid leukemia|9863/3
C0023473|T191|SY|0000007345|CHV|chronic myeloid leukemias|9863/3
C0023473|T191|SY|0000007345|CHV|cml|9863/3
C0023473|T191|PT|U000138|COSTAR|CHRONIC GRANULOCYTIC LEUKEMIA|9863/3
C0023473|T191|ET|2004-1700|CSP|chronic granulocytic leukemia|9863/3
C0023473|T191|ET|2004-1700|CSP|chronic myelocytic leukemia|9863/3
C0023473|T191|PT|2004-1700|CSP|chronic myelogenous leukemia|9863/3
C0023473|T191|ET|2004-1700|CSP|chronic myeloid leukemia|9863/3
C0023473|T191|ET|2004-1700|CSP|CML|9863/3
C0023473|T191|PT|LEUKEMIA CHRON MYELO|CST|CHRONIC MYELOCYTIC LEUKEMIA|9863/3
C0023473|T191|GT|LEUKEMIA CHRON MYELO|CST|LEUKEMIA MYELOCYTIC CHRONIC|9863/3
C0023473|T191|SY|NOCODE|DXP|CML|9863/3
C0023473|T191|SY|NOCODE|DXP|LEUKEMIA, GRANULOCYTIC, CHRONIC|9863/3
C0023473|T191|DI|U001052|DXP|LEUKEMIA, MYELOCYTIC, CHRONIC|9863/3
C0023473|T191|SY|NOCODE|DXP|LEUKEMIA, MYELOGENOUS, CHRONIC|9863/3
C0023473|T191|SY|NOCODE|DXP|LEUKEMIA, MYELOID, CHRONIC|9863/3
C0023473|T191|SY|HP:0005506|HPO|Chronic myelocytic leukemia|9863/3
C0023473|T191|PT|HP:0005506|HPO|Chronic myelogenous leukemia|9863/3
C0023473|T191|SY|HP:0005506|HPO|Chronic myeloid leukemia|9863/3
C0023473|T191|PT|C92.1|ICD10|Chronic myeloid leukaemia|9863/3
C0023473|T191|PT|C92.1|ICD10AE|Chronic myeloid leukemia|9863/3
C0023473|T191|HT|205.1|ICD9CM|Myeloid leukemia, chronic|9863/3
C0023473|T191|PT|MTHU016669|ICPC2ICD10ENG|chronic; myelosis|9863/3
C0023473|T191|PT|MTHU032697|ICPC2ICD10ENG|granulocytic; leukemia, chronic|9863/3
C0023473|T191|PT|MTHU044757|ICPC2ICD10ENG|leukemia; granulocytic, chronic|9863/3
C0023473|T191|PT|MTHU044782|ICPC2ICD10ENG|leukemia; myelocytic, chronic|9863/3
C0023473|T191|PT|MTHU044786|ICPC2ICD10ENG|leukemia; myeloid, chronic|9863/3
C0023473|T191|PT|MTHU050843|ICPC2ICD10ENG|myelocytic; leukemia, chronic|9863/3
C0023473|T191|PT|MTHU050857|ICPC2ICD10ENG|myeloid; leukemia, chronic|9863/3
C0023473|T191|PT|MTHU050919|ICPC2ICD10ENG|myelosis; chronic|9863/3
C0023473|T191|PTN|B73005|ICPC2P|chronic myeloid leukaemia|9863/3
C0023473|T191|MTH_PTN|B73005|ICPC2P|chronic myeloid leukemia|9863/3
C0023473|T191|PT|B73005|ICPC2P|Leukaemia;chronic myeloid|9863/3
C0023473|T191|MTH_PT|B73005|ICPC2P|Leukemia;chronic myeloid|9863/3
C0023473|T191|PT|sh2004008307|LCH_NW|Chronic myeloid leukemia|9863/3
C0023473|T191|LA|LA26791-6|LNC|Chronic myelogenous leukemia|9863/3
C0023473|T191|LLT|10008904|MDR|Chronic granulocytic leukaemia|9863/3
C0023473|T191|LLT|10008905|MDR|Chronic granulocytic leukemia|9863/3
C0023473|T191|LLT|10058245|MDR|Chronic myelocytic leukaemia|9863/3
C0023473|T191|LLT|10009011|MDR|Chronic myelocytic leukemia|9863/3
C0023473|T191|LLT|10058246|MDR|Chronic myelogenous leukaemia|9863/3
C0023473|T191|LLT|10009012|MDR|Chronic myelogenous leukemia|9863/3
C0023473|T191|LLT|10009013|MDR|Chronic myeloid leukaemia|9863/3
C0023473|T191|PT|10009013|MDR|Chronic myeloid leukaemia|9863/3
C0023473|T191|LLT|10009015|MDR|Chronic myeloid leukemia|9863/3
C0023473|T191|MTH_PT|10009013|MDR|Chronic myeloid leukemia|9863/3
C0023473|T191|LLT|10009700|MDR|CML|9863/3
C0023473|T191|LLT|10058247|MDR|Leukaemia myelocytic chronic|9863/3
C0023473|T191|HT|10024296|MDR|Leukaemias chronic myeloid|9863/3
C0023473|T191|LLT|10024347|MDR|Leukemia myelocytic chronic|9863/3
C0023473|T191|MTH_HT|10024296|MDR|Leukemias chronic myeloid|9863/3
C0023473|T191|LLT|10028553|MDR|Myeloid leukaemia, chronic|9863/3
C0023473|T191|LLT|10028558|MDR|Myeloid leukemia, chronic|9863/3
C0023473|T191|PT|31475|MEDCIN|chronic myelogenous leukemia|9863/3
C0023473|T191|SY|5624|MEDLINEPLUS|Chronic granulocytic leukemia|9863/3
C0023473|T191|ET|5624|MEDLINEPLUS|Chronic Granulocytic Leukemia|9863/3
C0023473|T191|ET|5624|MEDLINEPLUS|Chronic Myelogenous Leukemia|9863/3
C0023473|T191|SY|5624|MEDLINEPLUS|Chronic myelogenous leukemia|9863/3
C0023473|T191|PT|5624|MEDLINEPLUS|Chronic Myeloid Leukemia|9863/3
C0023473|T191|SY|5624|MEDLINEPLUS|CML|9863/3
C0023473|T191|ET|5624|MEDLINEPLUS|CML|9863/3
C0023473|T191|ET|5624|MEDLINEPLUS|Leukemia, Myeloid, Chronic|9863/3
C0023473|T191|PM|D015464|MSH|Chronic Granulocytic Leukemia|9863/3
C0023473|T191|PM|D015464|MSH|Chronic Granulocytic Leukemias|9863/3
C0023473|T191|PM|D015464|MSH|Chronic Myelocytic Leukemia|9863/3
C0023473|T191|PM|D015464|MSH|Chronic Myelocytic Leukemias|9863/3
C0023473|T191|PM|D015464|MSH|Chronic Myelogenous Leukemia|9863/3
C0023473|T191|PM|D015464|MSH|Chronic Myelogenous Leukemias|9863/3
C0023473|T191|PM|D015464|MSH|Chronic Myeloid Leukemia|9863/3
C0023473|T191|PM|D015464|MSH|Chronic Myeloid Leukemias|9863/3
C0023473|T191|ET|D015464|MSH|Granulocytic Leukemia, Chronic|9863/3
C0023473|T191|PM|D015464|MSH|Granulocytic Leukemias, Chronic|9863/3
C0023473|T191|DEV|D015464|MSH|LEUKEMIA PHILA POS|9863/3
C0023473|T191|PM|D015464|MSH|Leukemia, Chronic Granulocytic|9863/3
C0023473|T191|PM|D015464|MSH|Leukemia, Chronic Myelocytic|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Chronic Myelogenous|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Chronic Myeloid|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Granulocytic, Chronic|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myelocytic, Chronic|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myelogenous, Chronic|9863/3
C0023473|T191|MH|D015464|MSH|Leukemia, Myelogenous, Chronic, BCR-ABL Positive|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myelogenous, Ph1 Positive|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myelogenous, Ph1-Positive|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Chronic|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Ph1 Positive|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Ph1-Positive|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Philadelphia Positive|9863/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Philadelphia-Positive|9863/3
C0023473|T191|PM|D015464|MSH|Leukemia, Ph1-Positive Myelogenous|9863/3
C0023473|T191|PM|D015464|MSH|Leukemia, Ph1-Positive Myeloid|9863/3
C0023473|T191|PM|D015464|MSH|Leukemia, Philadelphia-Positive Myeloid|9863/3
C0023473|T191|PM|D015464|MSH|Leukemias, Chronic Granulocytic|9863/3
C0023473|T191|PM|D015464|MSH|Leukemias, Chronic Myelocytic|9863/3
C0023473|T191|PM|D015464|MSH|Leukemias, Chronic Myelogenous|9863/3
C0023473|T191|PM|D015464|MSH|Leukemias, Chronic Myeloid|9863/3
C0023473|T191|PM|D015464|MSH|Leukemias, Ph1-Positive Myelogenous|9863/3
C0023473|T191|PM|D015464|MSH|Leukemias, Ph1-Positive Myeloid|9863/3
C0023473|T191|PM|D015464|MSH|Leukemias, Philadelphia-Positive Myeloid|9863/3
C0023473|T191|ET|D015464|MSH|Myelocytic Leukemia, Chronic|9863/3
C0023473|T191|PM|D015464|MSH|Myelocytic Leukemias, Chronic|9863/3
C0023473|T191|ET|D015464|MSH|Myelogenous Leukemia, Chronic|9863/3
C0023473|T191|PM|D015464|MSH|Myelogenous Leukemia, Ph1 Positive|9863/3
C0023473|T191|ET|D015464|MSH|Myelogenous Leukemia, Ph1-Positive|9863/3
C0023473|T191|PM|D015464|MSH|Myelogenous Leukemias, Chronic|9863/3
C0023473|T191|PM|D015464|MSH|Myelogenous Leukemias, Ph1-Positive|9863/3
C0023473|T191|ET|D015464|MSH|Myeloid Leukemia, Chronic|9863/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemia, Ph1 Positive|9863/3
C0023473|T191|ET|D015464|MSH|Myeloid Leukemia, Ph1-Positive|9863/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemia, Philadelphia Positive|9863/3
C0023473|T191|ET|D015464|MSH|Myeloid Leukemia, Philadelphia-Positive|9863/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemias, Chronic|9863/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemias, Ph1-Positive|9863/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemias, Philadelphia-Positive|9863/3
C0023473|T191|PM|D015464|MSH|Ph1-Positive Myelogenous Leukemia|9863/3
C0023473|T191|PM|D015464|MSH|Ph1-Positive Myelogenous Leukemias|9863/3
C0023473|T191|PM|D015464|MSH|Ph1-Positive Myeloid Leukemia|9863/3
C0023473|T191|PM|D015464|MSH|Ph1-Positive Myeloid Leukemias|9863/3
C0023473|T191|PM|D015464|MSH|Philadelphia-Positive Myeloid Leukemia|9863/3
C0023473|T191|PM|D015464|MSH|Philadelphia-Positive Myeloid Leukemias|9863/3
C0023473|T191|PN|NOCODE|MTH|Myeloid Leukemia, Chronic|9863/3
C0023473|T191|SY|C3174|NCI|BCR-ABL Positive Chronic Myelogenous Leukemia|9863/3
C0023473|T191|SY|C3174|NCI|Chronic Granulocytic Leukemia|9863/3
C0023473|T191|SY|C3174|NCI|Chronic Myelocytic Leukemia|9863/3
C0023473|T191|SY|C3174|NCI|Chronic Myelogenous Leukemia|9863/3
C0023473|T191|PT|C3174|NCI|Chronic Myelogenous Leukemia, BCR-ABL1 Positive|9863/3
C0023473|T191|SY|TCGA|NCI|Chronic Myelogenous Leukemia, BCR-ABL1 Positive|9863/3
C0023473|T191|SY|C3174|NCI|Chronic Myelogenous Leukemias|9863/3
C0023473|T191|SY|C3174|NCI|Chronic Myeloid Leukemia|9863/3
C0023473|T191|AB|C3174|NCI|CML|9863/3
C0023473|T191|SY|C3174|NCI|CML - Chronic Myelogenous Leukemia|9863/3
C0023473|T191|PT|C3174|NCI_CPTAC|Chronic Myelogenous Leukemia, BCR-ABL1 Positive|9863/3
C0023473|T191|SY|C3174|NCI_CTRP|Chronic Myelogenous Leukemia, BCR-ABL1 Positive|9863/3
C0023473|T191|PT|CDR0000046754|NCI_NCI-GLOSS|chronic granulocytic leukemia|9863/3
C0023473|T191|PT|CDR0000044901|NCI_NCI-GLOSS|chronic myelogenous leukemia|9863/3
C0023473|T191|PT|CDR0000046755|NCI_NCI-GLOSS|chronic myeloid leukemia|9863/3
C0023473|T191|PT|CDR0000044382|NCI_NCI-GLOSS|CML|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|CGL|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|chronic granulocytic leukemia|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|chronic myelocytic leukemia|9863/3
C0023473|T191|PT|CDR0000037900|PDQ|chronic myelogenous leukemia|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|Chronic Myelogenous Leukemias|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|Chronic Myeloid Leukemia|9863/3
C0023473|T191|AB|CDR0000037900|PDQ|CML|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|CML - Chronic Myelogenous Leukemia|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|granulocytic leukemia, chronic|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|leukemia, chronic myelogenous|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|myelocytic leukemia, chronic|9863/3
C0023473|T191|SY|CDR0000037900|PDQ|myelogenous leukemia, chronic|9863/3
C0023473|T191|PT|R0121663|QMR|LEUKEMIA CHRONIC MYELOCYTIC|9863/3
C0023473|T191|AB|B651.|RCD|CGL - Chronic granul leukaemia|9863/3
C0023473|T191|SY|B651.|RCD|CGL - Chronic granulocytic leukaemia|9863/3
C0023473|T191|SY|B651.|RCD|Chronic granulocytic leukaemia|9863/3
C0023473|T191|PT|B651.|RCD|Chronic myeloid leukaemia|9863/3
C0023473|T191|OP|B651z|RCD|Chronic myeloid leukaemia NOS|9863/3
C0023473|T191|AB|B651.|RCD|CML - Chronic myeloid leukaem|9863/3
C0023473|T191|SY|B651.|RCD|CML - Chronic myeloid leukaemia|9863/3
C0023473|T191|AB|B651.|RCDAE|CGL - Chronic granul leukemia|9863/3
C0023473|T191|SY|B651.|RCDAE|CGL - Chronic granulocytic leukemia|9863/3
C0023473|T191|SY|B651.|RCDAE|Chronic granulocytic leukemia|9863/3
C0023473|T191|PT|B651.|RCDAE|Chronic myeloid leukemia|9863/3
C0023473|T191|OP|B651z|RCDAE|Chronic myeloid leukemia NOS|9863/3
C0023473|T191|SY|B651.|RCDAE|CML - Chronic myeloid leukemia|9863/3
C0023473|T191|OP|BBr63|RCDSA|Chronic myeloid leukemia|9863/3
C0023473|T191|OP|BBr63|RCDSY|Chronic myeloid leukaemia|9863/3
C0023473|T191|SYGB|92818009|SNOMEDCT_US|CGL - Chronic granulocytic leukaemia|9863/3
C0023473|T191|SY|92818009|SNOMEDCT_US|CGL - Chronic granulocytic leukemia|9863/3
C0023473|T191|SYGB|63364005|SNOMEDCT_US|Chronic granulocytic leukaemia|9863/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic granulocytic leukemia|9863/3
C0023473|T191|SYGB|92818009|SNOMEDCT_US|Chronic myelocytic leukaemia|9863/3
C0023473|T191|SYGB|63364005|SNOMEDCT_US|Chronic myelocytic leukaemia|9863/3
C0023473|T191|SY|92818009|SNOMEDCT_US|Chronic myelocytic leukemia|9863/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic myelocytic leukemia|9863/3
C0023473|T191|SYGB|63364005|SNOMEDCT_US|Chronic myelogenous leukaemia|9863/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic myelogenous leukemia|9863/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic myelogenous leukemia, no ICD-O subtype|9863/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic myelogenous leukemia, no International Classification of Diseases for Oncology subtype|9863/3
C0023473|T191|PTGB|92818009|SNOMEDCT_US|Chronic myeloid leukaemia|9863/3
C0023473|T191|PTGB|63364005|SNOMEDCT_US|Chronic myeloid leukaemia|9863/3
C0023473|T191|OAP|154592009|SNOMEDCT_US|Chronic myeloid leukaemia|9863/3
C0023473|T191|OF|154592009|SNOMEDCT_US|Chronic myeloid leukaemia|9863/3
C1531667|T191|PTGB|413841000|SNOMEDCT_US|Chronic myeloid leukaemia - category|9863/3
C0023473|T191|OAP|188735005|SNOMEDCT_US|Chronic myeloid leukaemia NOS|9863/3
C0023473|T191|SYGB|92818009|SNOMEDCT_US|Chronic myeloid leukaemia, disease|9863/3
C0023473|T191|PT|92818009|SNOMEDCT_US|Chronic myeloid leukemia|9863/3
C0023473|T191|PT|63364005|SNOMEDCT_US|Chronic myeloid leukemia|9863/3
C0023473|T191|OAP|154592009|SNOMEDCT_US|Chronic myeloid leukemia|9863/3
C1531667|T191|PT|413841000|SNOMEDCT_US|Chronic myeloid leukemia - category|9863/3
C0023473|T191|OAP|188735005|SNOMEDCT_US|Chronic myeloid leukemia NOS|9863/3
C0023473|T191|SY|92818009|SNOMEDCT_US|Chronic myeloid leukemia, disease|9863/3
C0023473|T191|SYGB|92818009|SNOMEDCT_US|CML - Chronic myeloid leukaemia|9863/3
C0023473|T191|SY|92818009|SNOMEDCT_US|CML - Chronic myeloid leukemia|9863/3
C0023487|T191|PT|0018064|CCPSS|LEUKEMIA ACUTE PROMYELOCYTIC|9866/3
C0023487|T191|SY|0000007351|CHV|acute promyelocytic leukaemia|9866/3
C0023487|T191|SY|0000057922|CHV|acute promyelocytic leukaemia|9866/3
C0023487|T191|SY|0000057922|CHV|acute promyelocytic leukemia|9866/3
C0023487|T191|PT|0000007351|CHV|acute promyelocytic leukemia|9866/3
C0023487|T191|SY|0000007351|CHV|acute promyelocytic leukemia apl|9866/3
C0023487|T191|SY|0000057922|CHV|fab m3|9866/3
C0023487|T191|SY|0000007351|CHV|fab m3|9866/3
C0023487|T191|PT|0000057922|CHV|M3 acute promyelocytic leukemia|9866/3
C0023487|T191|SY|0000007351|CHV|progranulocytic leukemia|9866/3
C0023487|T191|ET|4000-0108|CSP|acute promyelocytic leukemia|9866/3
C0023487|T191|ET|2004-4431|CSP|promyelocytic leukemia|9866/3
C0023487|T191|DI|U001054|DXP|LEUKEMIA, PROMYELOCYTIC|9866/3
C0023487|T191|PT|HP:0004836|HPO|Acute promyelocytic leukemia|9866/3
C0023487|T191|PT|C92.4|ICD10|Acute promyelocytic leukaemia|9866/3
C0023487|T191|PT|C92.4|ICD10AE|Acute promyelocytic leukemia|9866/3
C0023487|T191|HT|C92.4|ICD10CM|Acute promyelocytic leukemia|9866/3
C0023487|T191|AB|C92.4|ICD10CM|Acute promyelocytic leukemia|9866/3
C0023487|T191|ET|C92.40|ICD10CM|Acute promyelocytic leukemia NOS|9866/3
C0023487|T191|ET|C92.4|ICD10CM|AML M3|9866/3
C0023487|T191|PT|MTHU044796|ICPC2ICD10ENG|leukemia; promyelocytic|9866/3
C0023487|T191|PT|MTHU062048|ICPC2ICD10ENG|promyelocytic; leukemia|9866/3
C0023487|T191|LA|LA26788-2|LNC|Acute promyelocytic leukemia|9866/3
C0023487|T191|LLT|10001019|MDR|Acute promyelocytic leukaemia|9866/3
C0023487|T191|PT|10001019|MDR|Acute promyelocytic leukaemia|9866/3
C0023487|T191|LLT|10001020|MDR|Acute promyelocytic leukemia|9866/3
C0023487|T191|MTH_PT|10001019|MDR|Acute promyelocytic leukemia|9866/3
C0023487|T191|PT|31481|MEDCIN|acute promyelocytic leukemia|9866/3
C0023487|T191|SY|31481|MEDCIN|leukemia acute promyelocytic|9866/3
C0023487|T191|ET|D015473|MSH|Acute Promyelocytic Leukemia|9866/3
C0023487|T191|PM|D015473|MSH|Acute Promyelocytic Leukemias|9866/3
C0023487|T191|ET|D015473|MSH|AML M3|9866/3
C0023487|T191|PM|D015473|MSH|ANLL, M3|9866/3
C0023487|T191|DSV|D015473|MSH|LEUKEMIA MYELOID ACUTE M 03|9866/3
C0023487|T191|ET|D015473|MSH|Leukemia, Acute Promyelocytic|9866/3
C0023487|T191|ET|D015473|MSH|Leukemia, Myeloid, Acute, M3|9866/3
C0023487|T191|ET|D015473|MSH|Leukemia, Progranulocytic|9866/3
C0023487|T191|MH|D015473|MSH|Leukemia, Promyelocytic, Acute|9866/3
C0023487|T191|ET|D015473|MSH|M3 ANLL|9866/3
C0023487|T191|DSV|D015473|MSH|MYELOID LEUKEMIA ACUTE M 03|9866/3
C0023487|T191|ET|D015473|MSH|Myeloid Leukemia, Acute, M3|9866/3
C0023487|T191|ET|D015473|MSH|Progranulocytic Leukemia|9866/3
C0023487|T191|ET|D015473|MSH|Promyelocytic Leukemia, Acute|9866/3
C0023487|T191|PN|NOCODE|MTH|Acute Promyelocytic Leukemia|9866/3
C0023487|T191|ET|205.0|MTHICD9|Acute promyelocytic leukemia|9866/3
C0023487|T191|SY|C3182|NCI|Acute Promyelocytic Leukemia|9866/3
C0023487|T191|PT|C3182|NCI|Acute Promyelocytic Leukemia with PML-RARA|9866/3
C0023487|T191|AB|C3182|NCI|APL|9866/3
C0023487|T191|AB|C3182|NCI|APML|9866/3
C0023487|T191|SY|C3182|NCI|APML - Acute promyelocytic leukemia|9866/3
C0023487|T191|SY|C3182|NCI|FAB M3|9866/3
C0023487|T191|SY|C3182|NCI|Promyelocytic Leukemia|9866/3
C0023487|T191|PT|C3182|NCI_CPTAC|Acute Promyelocytic Leukemia with PML-RARA|9866/3
C0023487|T191|PT|10001019|NCI_CTEP-SDC|Acute promyelocytic leukemia|9866/3
C0023487|T191|SY|CDR0000444957|NCI_NCI-GLOSS|acute promyelocytic leukemia|9866/3
C0023487|T191|PT|CDR0000522912|NCI_NCI-GLOSS|APL|9866/3
C0023487|T191|PT|CDR0000046159|NCI_NCI-GLOSS|promyelocytic leukemia|9866/3
C0023487|T191|SY|C3182|NCI_NICHD|Acute Promyelocytic Leukemia|9866/3
C0023487|T191|SY|C3182|NCI_NICHD|APL|9866/3
C0023487|T191|SY|C3182|NCI_NICHD|APML|9866/3
C0023487|T191|PT|B65y1|RCD|Acute promyelocytic leukaemia|9866/3
C0023487|T191|AB|B65y1|RCD|APL - Acute promyelocytic leuk|9866/3
C0023487|T191|SY|B65y1|RCD|APL - Acute promyelocytic leukaemia|9866/3
C0023487|T191|AB|B65y1|RCD|APML - Acute promyel leukaemia|9866/3
C0023487|T191|SY|B65y1|RCD|APML - Acute promyelocytic leukaemia|9866/3
C0023487|T191|AB|B65y1|RCD|M3 - Acute promyelocyt leukaem|9866/3
C0023487|T191|SY|B65y1|RCD|M3 - Acute promyelocytic leukaemia|9866/3
C0023487|T191|PT|B65y1|RCDAE|Acute promyelocytic leukemia|9866/3
C0023487|T191|SY|B65y1|RCDAE|APL - Acute promyelocytic leukemia|9866/3
C0023487|T191|AB|B65y1|RCDAE|APML - Acute promyel leukemia|9866/3
C0023487|T191|SY|B65y1|RCDAE|APML - Acute promyelocytic leukemia|9866/3
C0023487|T191|SY|B65y1|RCDAE|M3 - Acute promyelocytic leukemia|9866/3
C0023487|T191|PT|BBr66|RCDSA|Acute promyelocytic leukemia|9866/3
C0023487|T191|AB|BBr66|RCDSY|Acute promyelocytic leukaem|9866/3
C0023487|T191|PT|BBr66|RCDSY|Acute promyelocytic leukaemia|9866/3
C0023487|T191|SYGB|28950004|SNOMEDCT_US|Acute myeloid leukaemia, PML/RAR-alpha|9866/3
C0023487|T191|SY|28950004|SNOMEDCT_US|Acute myeloid leukemia, PML/RAR-alpha|9866/3
C0023487|T191|PTGB|28950004|SNOMEDCT_US|Acute promyelocytic leukaemia|9866/3
C0023487|T191|PTGB|110004001|SNOMEDCT_US|Acute promyelocytic leukaemia, FAB M3|9866/3
C0023487|T191|SYGB|28950004|SNOMEDCT_US|Acute promyelocytic leukaemia, PML/RAR-alpha|9866/3
C0023487|T191|PT|28950004|SNOMEDCT_US|Acute promyelocytic leukemia|9866/3
C0023487|T191|PT|110004001|SNOMEDCT_US|Acute promyelocytic leukemia, FAB M3|9866/3
C0023487|T191|SY|28950004|SNOMEDCT_US|Acute promyelocytic leukemia, PML/RAR-alpha|9866/3
C0023487|T191|SYGB|110004001|SNOMEDCT_US|APL - Acute promyelocytic leukaemia|9866/3
C0023487|T191|SY|110004001|SNOMEDCT_US|APL - Acute promyelocytic leukemia|9866/3
C0023487|T191|SYGB|110004001|SNOMEDCT_US|APML - Acute promyelocytic leukaemia|9866/3
C0023487|T191|SY|110004001|SNOMEDCT_US|APML - Acute promyelocytic leukemia|9866/3
C0023487|T191|SY|28950004|SNOMEDCT_US|FAB M3|9866/3
C0023487|T191|SYGB|110004001|SNOMEDCT_US|M3 - Acute promyelocytic leukaemia|9866/3
C0023487|T191|SY|110004001|SNOMEDCT_US|M3 - Acute promyelocytic leukemia|9866/3
C0023479|T191|SY|0000007346|CHV|acute myelomonocytic leukaemia|9867/3
C0023479|T191|PT|0000007346|CHV|acute myelomonocytic leukemia|9867/3
C0023479|T191|SY|0000007346|CHV|m4 acute myeloid leukemia|9867/3
C0023479|T191|SY|0000007346|CHV|myeloblastic leukemia|9867/3
C0023479|T191|PT|HP:0004820|HPO|Acute myelomonocytic leukemia|9867/3
C0023479|T191|PT|C92.5|ICD10|Acute myelomonocytic leukaemia|9867/3
C0023479|T191|PT|C92.5|ICD10AE|Acute myelomonocytic leukemia|9867/3
C0023479|T191|AB|C92.5|ICD10CM|Acute myelomonocytic leukemia|9867/3
C0023479|T191|HT|C92.5|ICD10CM|Acute myelomonocytic leukemia|9867/3
C0023479|T191|ET|C92.50|ICD10CM|Acute myelomonocytic leukemia NOS|9867/3
C0023479|T191|ET|C92.5|ICD10CM|AML M4|9867/3
C0023479|T191|PT|MTHU003166|ICPC2ICD10ENG|acute; myelosis|9867/3
C0023479|T191|PT|MTHU011166|ICPC2ICD10ENG|blastic; leukemia, granulocytic|9867/3
C0023479|T191|PT|MTHU032696|ICPC2ICD10ENG|granulocytic; leukemia, blastic|9867/3
C0023479|T191|PT|MTHU044749|ICPC2ICD10ENG|leukemia; blastic, granulocytic|9867/3
C0023479|T191|PT|MTHU044756|ICPC2ICD10ENG|leukemia; granulocytic, blastic|9867/3
C0023479|T191|PT|MTHU044779|ICPC2ICD10ENG|leukemia; myeloblastic|9867/3
C0023479|T191|PT|MTHU044789|ICPC2ICD10ENG|leukemia; myelomonocytic, acute|9867/3
C0023479|T191|PT|MTHU044792|ICPC2ICD10ENG|leukemia; Naegeli-type monocytic|9867/3
C0023479|T191|PT|MTHU050295|ICPC2ICD10ENG|monocytic; leukemia, Naegeli-type|9867/3
C0023479|T191|PT|MTHU050838|ICPC2ICD10ENG|myeloblastic; leukemia|9867/3
C0023479|T191|PT|MTHU050873|ICPC2ICD10ENG|myelomonocytic; leukemia, acute|9867/3
C0023479|T191|PT|MTHU050917|ICPC2ICD10ENG|myelosis; acute|9867/3
C0023479|T191|PT|MTHU051490|ICPC2ICD10ENG|Naegeli-type monocytic; leukemia|9867/3
C0023479|T191|LLT|10000890|MDR|Acute myelomonocytic leukaemia|9867/3
C0023479|T191|PT|10000890|MDR|Acute myelomonocytic leukaemia|9867/3
C0023479|T191|LLT|10054297|MDR|Acute myelomonocytic leukemia|9867/3
C0023479|T191|MTH_PT|10000890|MDR|Acute myelomonocytic leukemia|9867/3
C0023479|T191|PT|230916|MEDCIN|acute myelomonocytic leukemia|9867/3
C0023479|T191|SY|230916|MEDCIN|leukemia acute myelomonocytic|9867/3
C0023479|T191|PM|D015479|MSH|Acute Myelomonocytic Leukemia|9867/3
C0023479|T191|PM|D015479|MSH|Acute Myelomonocytic Leukemias|9867/3
C0023479|T191|DSV|D015479|MSH|LEUKEMIA MYELOID ACUTE M 04|9867/3
C0023479|T191|PM|D015479|MSH|Leukemia, Acute Myelomonocytic|9867/3
C0023479|T191|ET|D015479|MSH|Leukemia, Myeloid, Acute, M4|9867/3
C0023479|T191|ET|D015479|MSH|Leukemia, Myeloid, Naegeli-Type|9867/3
C0023479|T191|MH|D015479|MSH|Leukemia, Myelomonocytic, Acute|9867/3
C0023479|T191|PM|D015479|MSH|Leukemia, Naegeli-Type Myeloid|9867/3
C0023479|T191|PM|D015479|MSH|Leukemias, Acute Myelomonocytic|9867/3
C0023479|T191|DSV|D015479|MSH|MYELOID LEUKEMIA ACUTE M 04|9867/3
C0023479|T191|ET|D015479|MSH|Myeloid Leukemia, Acute, M4|9867/3
C0023479|T191|PM|D015479|MSH|Myeloid Leukemia, Naegeli Type|9867/3
C0023479|T191|ET|D015479|MSH|Myeloid Leukemia, Naegeli-Type|9867/3
C0023479|T191|ET|D015479|MSH|Myelomonocytic Leukemia, Acute|9867/3
C0023479|T191|PM|D015479|MSH|Myelomonocytic Leukemias, Acute|9867/3
C0023479|T191|PM|D015479|MSH|Naegeli-Type Myeloid Leukemia|9867/3
C0023479|T191|PN|NOCODE|MTH|Acute myelomonocytic leukemia|9867/3
C0023479|T191|SY|C7463|NCI|Acute M4 Myeloid Leukemia|9867/3
C0023479|T191|PT|C7463|NCI|Acute Myelomonocytic Leukemia|9867/3
C0023479|T191|SY|TCGA|NCI|Acute Myelomonocytic Leukemia|9867/3
C0023479|T191|AB|C7463|NCI|AMML|9867/3
C0023479|T191|PT|C7463|NCI_CPTAC|Acute Myelomonocytic Leukemia|9867/3
C0023479|T191|PT|C7463|NCI_NICHD|Acute Myelomonocytic Leukemia|9867/3
C0023479|T191|PT|B690.|RCD|Acute myelomonocytic leukaemia|9867/3
C0023479|T191|AB|B690.|RCD|AMML - Acut myelomon leukaemia|9867/3
C0023479|T191|SY|B690.|RCD|AMML - Acute myelomonocytic leukaemia|9867/3
C0023479|T191|AB|B690.|RCD|M4 - Acute myelomonocy leukaem|9867/3
C0023479|T191|SY|B690.|RCD|M4 - Acute myelomonocytic leukaemia|9867/3
C0023479|T191|AB|Xa0Sl|RCD|Naegeli-type monocyt leukaemia|9867/3
C0023479|T191|SY|Xa0Sl|RCD|Naegeli-type monocytic leukaemia|9867/3
C0023479|T191|PT|B690.|RCDAE|Acute myelomonocytic leukemia|9867/3
C0023479|T191|AB|B690.|RCDAE|AMML - Acut myelomon leukemia|9867/3
C0023479|T191|SY|B690.|RCDAE|AMML - Acute myelomonocytic leukemia|9867/3
C0023479|T191|SY|B690.|RCDAE|M4 - Acute myelomonocytic leukemia|9867/3
C0023479|T191|AB|Xa0Sl|RCDAE|Naegeli-type monocyt leukemia|9867/3
C0023479|T191|SY|Xa0Sl|RCDAE|Naegeli-type monocytic leukemia|9867/3
C0023479|T191|OP|BBr67|RCDSA|Acute myelomonocytic leukemia|9867/3
C0023479|T191|OA|BBr67|RCDSY|Acte myelomonocytic leukaem|9867/3
C0023479|T191|OP|BBr67|RCDSY|Acute myelomonocytic leukaemia|9867/3
C0023479|T191|PTGB|30962008|SNOMEDCT_US|Acute myelomonocytic leukaemia|9867/3
C0023479|T191|PTGB|110005000|SNOMEDCT_US|Acute myelomonocytic leukaemia, FAB M4|9867/3
C0023479|T191|PT|30962008|SNOMEDCT_US|Acute myelomonocytic leukemia|9867/3
C0023479|T191|PT|110005000|SNOMEDCT_US|Acute myelomonocytic leukemia, FAB M4|9867/3
C0023479|T191|SYGB|110005000|SNOMEDCT_US|AMML - Acute myelomonocytic leukaemia|9867/3
C0023479|T191|SY|110005000|SNOMEDCT_US|AMML - Acute myelomonocytic leukemia|9867/3
C0023479|T191|SY|30962008|SNOMEDCT_US|FAB M4|9867/3
C0023479|T191|SYGB|110005000|SNOMEDCT_US|M4 - Acute myelomonocytic leukaemia|9867/3
C0023479|T191|SY|110005000|SNOMEDCT_US|M4 - Acute myelomonocytic leukemia|9867/3
C0023479|T191|SYGB|277601005|SNOMEDCT_US|Naegeli-type monocytic leukaemia|9867/3
C0023479|T191|SY|277601005|SNOMEDCT_US|Naegeli-type monocytic leukemia|9867/3
C0023437|T191|ET|C94.8|ICD10CM|Acute basophilic leukemia|9870/3
C0023437|T191|PT|230919|MEDCIN|acute basophilic leukemia|9870/3
C0023437|T191|SY|230919|MEDCIN|leukemia acute basophilic|9870/3
C0023437|T191|PM|D015471|MSH|Acute Basophilic Leukemia|9870/3
C0023437|T191|PM|D015471|MSH|Acute Basophilic Leukemias|9870/3
C0023437|T191|ET|D015471|MSH|Basophilic Leukemia, Acute|9870/3
C0023437|T191|PM|D015471|MSH|Basophilic Leukemias, Acute|9870/3
C0023437|T191|PM|D015471|MSH|Leukemia, Acute Basophilic|9870/3
C0023437|T191|MH|D015471|MSH|Leukemia, Basophilic, Acute|9870/3
C0023437|T191|PM|D015471|MSH|Leukemias, Acute Basophilic|9870/3
C0023437|T191|PN|NOCODE|MTH|Acute Basophilic Leukemia|9870/3
C0023437|T191|SY|TCGA|NCI|Acute Basophilic Leukemia|9870/3
C0023437|T191|PT|C3164|NCI|Acute Basophilic Leukemia|9870/3
C0023437|T191|SY|C3164|NCI|Basophilic Leukemia|9870/3
C0023437|T191|SY|C3164|NCI|Leukemia Basophilic|9870/3
C0023437|T191|PT|C3164|NCI_NICHD|Acute Basophilic Leukemia|9870/3
C0023437|T191|PTGB|69077002|SNOMEDCT_US|Acute basophilic leukaemia|9870/3
C0023437|T191|PT|69077002|SNOMEDCT_US|Acute basophilic leukemia|9870/3
C0522630|T191|SY|C9287|NCI|Acute Myeloid Leukemia with Abnormal Marrow Eosinophils|9871/3
C0522630|T191|SY|C9287|NCI|Acute Myeloid Leukemia, CBF-beta/MYH11|9871/3
C0522630|T191|SY|C9287|NCI|Acute Myeloid Leukemia, CBFB-MYH11|9871/3
C0522630|T191|SYGB|103688009|SNOMEDCT_US|Acute myeloid leukaemia, CBF-beta/MYH11|9871/3
C0522630|T191|PT|103688009|SNOMEDCT_US|Acute myeloid leukemia with abnormal marrow eosinophils|9871/3
C0522630|T191|SY|103688009|SNOMEDCT_US|Acute myeloid leukemia, CBF-beta/MYH11|9871/3
C0522631|T191|ET|C92.0|ICD10CM|Acute myeloblastic leukemia M0|9872/3
C0522631|T191|ET|C92.0|ICD10CM|Acute myeloblastic leukemia, minimal differentiation|9872/3
C0522631|T191|LLT|10000885|MDR|Acute myeloid leukaemia with minimal differentiation|9872/3
C0522631|T191|LLT|10000888|MDR|Acute myeloid leukemia with minimal differentiation|9872/3
C0522631|T191|SY|C8460|NCI|Acute Myeloblastic Leukemia with Minimal Differentiation|9872/3
C0522631|T191|SY|C8460|NCI|Acute Myeloblastic Leukemia, Minimally Differentiated|9872/3
C0522631|T191|SY|C8460|NCI|Acute Myelocytic Leukemia with Minimal Differentiation|9872/3
C0522631|T191|SY|C8460|NCI|Acute Myelogenous Leukemia with Minimal Differentiation|9872/3
C0522631|T191|PT|C8460|NCI|Acute Myeloid Leukemia with Minimal Differentiation|9872/3
C0522631|T191|SY|TCGA|NCI|Acute Myeloid Leukemia with Minimal Differentiation|9872/3
C0522631|T191|SY|C8460|NCI|Acute Myeloid Leukemia, Minimally Differentiated|9872/3
C0522631|T191|SY|C8460|NCI|AML with Minimal Differentiation|9872/3
C0522631|T191|SY|C8460|NCI|M0 Acute Granulocytic Leukemia|9872/3
C0522631|T191|SY|C8460|NCI|M0 Acute Granulocytic Leukemia with Minimal Differentiation|9872/3
C0522631|T191|SY|C8460|NCI|M0 Acute Myeloblastic Leukemia|9872/3
C0522631|T191|SY|C8460|NCI|M0 Acute Myelocytic Leukemia|9872/3
C0522631|T191|SY|C8460|NCI|M0 Acute Myelogenous Leukemia|9872/3
C0522631|T191|SY|C8460|NCI|M0 Acute Myelogenous Leukemia with Minimal Differentiation|9872/3
C0522631|T191|SY|C8460|NCI|M0 Myeloid Leukemia|9872/3
C0522631|T191|SY|C8460|NCI|M0 Myeloid Leukemia with Minimal Differentiation|9872/3
C0522631|T191|PT|C8460|NCI_NICHD|Acute Myeloid Leukemia with Minimal Differentiation|9872/3
C0522631|T191|SYGB|103689001|SNOMEDCT_US|Acute granulocytic leukaemia, minimal differentiation|9872/3
C0522631|T191|SY|103689001|SNOMEDCT_US|Acute granulocytic leukemia, minimal differentiation|9872/3
C0522631|T191|SYGB|103689001|SNOMEDCT_US|Acute myeloblastic leukaemia, minimal differentiation|9872/3
C0522631|T191|SY|103689001|SNOMEDCT_US|Acute myeloblastic leukemia, minimal differentiation|9872/3
C0522631|T191|SYGB|103689001|SNOMEDCT_US|Acute myelocytic leukaemia, minimal differentiation|9872/3
C0522631|T191|SY|103689001|SNOMEDCT_US|Acute myelocytic leukemia, minimal differentiation|9872/3
C0522631|T191|SYGB|103689001|SNOMEDCT_US|Acute myelogenous leukaemia, minimal differentiation|9872/3
C0522631|T191|SY|103689001|SNOMEDCT_US|Acute myelogenous leukemia, minimal differentiation|9872/3
C0522631|T191|PTGB|103689001|SNOMEDCT_US|Acute myeloid leukaemia, minimal differentiation|9872/3
C0522631|T191|PT|103689001|SNOMEDCT_US|Acute myeloid leukemia, minimal differentiation|9872/3
C0522631|T191|SY|103689001|SNOMEDCT_US|FAB M0|9872/3
C0026998|T191|ET|C92.0|ICD10CM|Acute myeloblastic leukemia M1|9873/3
C0026998|T191|PT|230920|MEDCIN|acute myelogenous leukemia without maturation|9873/3
C0026998|T191|SY|230920|MEDCIN|AML FAB-M1|9873/3
C0026998|T191|SY|230920|MEDCIN|AML without maturation|9873/3
C0026998|T191|ET|D015470|MSH|Acute Myeloid Leukemia without Maturation|9873/3
C0026998|T191|ET|D015470|MSH|Leukemia, Myeloid, Acute, M1|9873/3
C0026998|T191|PEP|D015470|MSH|Myeloid Leukemia, Acute, M1|9873/3
C0026998|T191|PN|NOCODE|MTH|Acute Myeloid Leukemia, M1|9873/3
C0026998|T191|SY|C3249|NCI|Acute Granulocytic Leukemia without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|Acute M1 Myeloid Leukemia|9873/3
C0026998|T191|SY|C3249|NCI|Acute Myeloblastic Leukemia without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|Acute Myelocytic Leukemia without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|Acute Myelogenous Leukemia without Maturation|9873/3
C0026998|T191|PT|C3249|NCI|Acute Myeloid Leukemia without Maturation|9873/3
C0026998|T191|SY|TCGA|NCI|Acute Myeloid Leukemia without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|AML without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|FAB M1|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Granulocytic Leukemia|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Granulocytic Leukemia without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Myeloblastic Leukemia|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Myeloblastic Leukemia without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Myelocytic Leukemia|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Myelocytic Leukemia without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Myelogenous Leukemia|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Myelogenous Leukemia without Maturation|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Myeloid Leukemia|9873/3
C0026998|T191|SY|C3249|NCI|M1 Acute Myeloid Leukemia without Maturation|9873/3
C0026998|T191|PT|C3249|NCI_NICHD|Acute Myeloid Leukemia without Maturation|9873/3
C0026998|T191|AB|Xa3Ea|RCD|Acute myelo leuk without matn|9873/3
C0026998|T191|PT|Xa3Ea|RCD|Acute myeloblastic leukaemia without maturation|9873/3
C0026998|T191|AB|Xa3Ea|RCD|M1 - Acut myel leuk -no maturn|9873/3
C0026998|T191|SY|Xa3Ea|RCD|M1 - Acute myeloblastic leukaemia without maturation|9873/3
C0026998|T191|PT|Xa3Ea|RCDAE|Acute myeloblastic leukemia without maturation|9873/3
C0026998|T191|SY|Xa3Ea|RCDAE|M1 - Acute myeloblastic leukemia without maturation|9873/3
C0026998|T191|SYGB|103690005|SNOMEDCT_US|Acute granulocytic leukaemia without maturation|9873/3
C0026998|T191|SY|103690005|SNOMEDCT_US|Acute granulocytic leukemia without maturation|9873/3
C0026998|T191|SYGB|103690005|SNOMEDCT_US|Acute myeloblastic leukaemia without maturation|9873/3
C0026998|T191|OAP|285766002|SNOMEDCT_US|Acute myeloblastic leukaemia without maturation|9873/3
C0026998|T191|OAP|285766002|SNOMEDCT_US|Acute myeloblastic leukemia without maturation|9873/3
C0026998|T191|SY|103690005|SNOMEDCT_US|Acute myeloblastic leukemia without maturation|9873/3
C0026998|T191|SYGB|103690005|SNOMEDCT_US|Acute myelocytic leukaemia without maturation|9873/3
C0026998|T191|SY|103690005|SNOMEDCT_US|Acute myelocytic leukemia without maturation|9873/3
C0026998|T191|SYGB|359640008|SNOMEDCT_US|Acute myelogenous leukaemia without maturation|9873/3
C0026998|T191|SYGB|103690005|SNOMEDCT_US|Acute myelogenous leukaemia without maturation|9873/3
C0026998|T191|OAP|359636004|SNOMEDCT_US|Acute myelogenous leukaemia without maturation, FAB M1|9873/3
C0026998|T191|SY|103690005|SNOMEDCT_US|Acute myelogenous leukemia without maturation|9873/3
C0026998|T191|SY|359640008|SNOMEDCT_US|Acute myelogenous leukemia without maturation|9873/3
C0026998|T191|IS|127223004|SNOMEDCT_US|Acute myelogenous leukemia without maturation, FAB M1|9873/3
C0026998|T191|OAP|359636004|SNOMEDCT_US|Acute myelogenous leukemia without maturation, FAB M1|9873/3
C0026998|T191|PTGB|103690005|SNOMEDCT_US|Acute myeloid leukaemia without maturation|9873/3
C0026998|T191|PTGB|359640008|SNOMEDCT_US|Acute myeloid leukaemia without maturation, FAB M1|9873/3
C0026998|T191|OAP|127223004|SNOMEDCT_US|Acute myeloid leukaemia without maturation, FAB M1|9873/3
C0026998|T191|PT|103690005|SNOMEDCT_US|Acute myeloid leukemia without maturation|9873/3
C0026998|T191|OAP|127223004|SNOMEDCT_US|Acute myeloid leukemia without maturation, FAB M1|9873/3
C0026998|T191|PT|359640008|SNOMEDCT_US|Acute myeloid leukemia without maturation, FAB M1|9873/3
C0026998|T191|SY|103690005|SNOMEDCT_US|FAB M1|9873/3
C0026998|T191|OAS|285766002|SNOMEDCT_US|M1 - Acute myeloblastic leukaemia without maturation|9873/3
C0026998|T191|SYGB|359640008|SNOMEDCT_US|M1 - Acute myeloblastic leukaemia without maturation|9873/3
C0026998|T191|OAS|285766002|SNOMEDCT_US|M1 - Acute myeloblastic leukemia without maturation|9873/3
C0026998|T191|SY|359640008|SNOMEDCT_US|M1 - Acute myeloblastic leukemia without maturation|9873/3
C1879321|T191|ET|C92.0|ICD10CM|Acute myeloblastic leukemia M2|9874/3
C1879321|T191|PT|230921|MEDCIN|acute myelogenous leukemia with maturation|9874/3
C1879321|T191|SY|230921|MEDCIN|AML with maturation|9874/3
C1879321|T191|ET|D015470|MSH|Acute Myeloid Leukemia with Maturation|9874/3
C1879321|T191|PEP|D015470|MSH|Leukemia, Myeloid, Acute, M2|9874/3
C1879321|T191|ET|D015470|MSH|Myeloid Leukemia, Acute, M2|9874/3
C1879321|T191|SY|C3250|NCI|Acute M2 Myeloid Leukemia|9874/3
C1879321|T191|SY|C3250|NCI|Acute Myeloblastic Leukemia with Maturation|9874/3
C1879321|T191|SY|C3250|NCI|Acute Myelocytic Leukemia with Maturation|9874/3
C1879321|T191|SY|C3250|NCI|Acute Myelogenous Leukemia with Maturation|9874/3
C1879321|T191|PT|C3250|NCI|Acute Myeloid Leukemia with Maturation|9874/3
C1879321|T191|SY|TCGA|NCI|Acute Myeloid Leukemia with Maturation|9874/3
C1879321|T191|SY|C3250|NCI|AML with Maturation|9874/3
C1879321|T191|SY|C3250|NCI|FAB M2|9874/3
C1879321|T191|SY|C3250|NCI|M2 Acute Granulocytic Leukemia|9874/3
C1879321|T191|SY|C3250|NCI|M2 Acute Myeloblastic Leukemia|9874/3
C1879321|T191|SY|C3250|NCI|M2 Acute Myeloblastic Leukemia with Maturation|9874/3
C1879321|T191|SY|C3250|NCI|M2 Acute Myelocytic Leukemia with Maturation|9874/3
C1879321|T191|SY|C3250|NCI|M2 Acute Myelogenous Leukemia|9874/3
C1879321|T191|SY|C3250|NCI|M2 Acute Myelogenous Leukemia with Maturation|9874/3
C1879321|T191|SY|C3250|NCI|M2 Acute Myeloid Leukemia|9874/3
C1879321|T191|SY|C3250|NCI|M2 Acute Myeloid Leukemia with Maturation|9874/3
C1879321|T191|PT|C3250|NCI_NICHD|Acute Myeloid Leukemia with Maturation|9874/3
C1879321|T191|AB|Xa3Ec|RCD|Acute myelo leuk with matn|9874/3
C1879321|T191|PT|Xa3Ec|RCD|Acute myeloblastic leukaemia with maturation|9874/3
C1879321|T191|AB|Xa3Ec|RCD|M2 - Ac myel leuk with maturn|9874/3
C1879321|T191|SY|Xa3Ec|RCD|M2 - Acute myeloblastic leukaemia with maturation|9874/3
C1879321|T191|PT|Xa3Ec|RCDAE|Acute myeloblastic leukemia with maturation|9874/3
C1879321|T191|SY|Xa3Ec|RCDAE|M2 - Acute myeloblastic leukemia with maturation|9874/3
C1879321|T191|SYGB|103691009|SNOMEDCT_US|Acute granulocytic leukaemia with maturation|9874/3
C1879321|T191|SY|103691009|SNOMEDCT_US|Acute granulocytic leukemia with maturation|9874/3
C1879321|T191|SYGB|103691009|SNOMEDCT_US|Acute myeloblastic leukaemia with maturation|9874/3
C1879321|T191|OAP|285768001|SNOMEDCT_US|Acute myeloblastic leukaemia with maturation|9874/3
C1879321|T191|OAP|285768001|SNOMEDCT_US|Acute myeloblastic leukemia with maturation|9874/3
C1879321|T191|SY|103691009|SNOMEDCT_US|Acute myeloblastic leukemia with maturation|9874/3
C1879321|T191|SYGB|103691009|SNOMEDCT_US|Acute myelocytic leukaemia with maturation|9874/3
C1879321|T191|SY|103691009|SNOMEDCT_US|Acute myelocytic leukemia with maturation|9874/3
C1879321|T191|SYGB|103691009|SNOMEDCT_US|Acute myelogenous leukaemia with maturation|9874/3
C1879321|T191|OAP|359645003|SNOMEDCT_US|Acute myelogenous leukaemia with maturation, FAB M2|9874/3
C1879321|T191|SY|103691009|SNOMEDCT_US|Acute myelogenous leukemia with maturation|9874/3
C1879321|T191|IS|127224005|SNOMEDCT_US|Acute myelogenous leukemia with maturation, FAB M2|9874/3
C1879321|T191|OAP|359645003|SNOMEDCT_US|Acute myelogenous leukemia with maturation, FAB M2|9874/3
C1879321|T191|OF|359645003|SNOMEDCT_US|Acute myelogenous leukemia with maturation, FAB M2|9874/3
C1879321|T191|PTGB|103691009|SNOMEDCT_US|Acute myeloid leukaemia with maturation|9874/3
C1879321|T191|PTGB|359648001|SNOMEDCT_US|Acute myeloid leukaemia with maturation, FAB M2|9874/3
C1879321|T191|OAP|127224005|SNOMEDCT_US|Acute myeloid leukaemia with maturation, FAB M2|9874/3
C1879321|T191|PT|103691009|SNOMEDCT_US|Acute myeloid leukemia with maturation|9874/3
C1879321|T191|OAP|127224005|SNOMEDCT_US|Acute myeloid leukemia with maturation, FAB M2|9874/3
C1879321|T191|PT|359648001|SNOMEDCT_US|Acute myeloid leukemia with maturation, FAB M2|9874/3
C1879321|T191|SY|103691009|SNOMEDCT_US|FAB M2|9874/3
C1879321|T191|OAS|285768001|SNOMEDCT_US|M2 - Acute myeloblastic leukaemia with maturation|9874/3
C1879321|T191|SYGB|359648001|SNOMEDCT_US|M2 - Acute myeloblastic leukaemia with maturation|9874/3
C1879321|T191|SY|359648001|SNOMEDCT_US|M2 - Acute myeloblastic leukemia with maturation|9874/3
C1879321|T191|OAS|285768001|SNOMEDCT_US|M2 - Acute myeloblastic leukemia with maturation|9874/3
C0023473|T191|PT|BI00304|BI|chronic myelogenous leukemia|9875/3
C0023473|T191|AB|BI00304|BI|cml|9875/3
C0023473|T191|PT|0003456|CCPSS|LEUKEMIA CHRONIC MYELOGENOUS|9875/3
C0023473|T191|SY|0000007345|CHV|chronic granulocytic leukaemia|9875/3
C0023473|T191|SY|0000007345|CHV|chronic granulocytic leukemia|9875/3
C0023473|T191|SY|0000007345|CHV|chronic myelocytic leukemia|9875/3
C0023473|T191|SY|0000007345|CHV|chronic myelogenous leukaemia|9875/3
C0023473|T191|SY|0000007345|CHV|chronic myelogenous leukemia|9875/3
C0023473|T191|SY|0000007345|CHV|chronic myeloid leukaemia|9875/3
C0023473|T191|SY|0000007345|CHV|chronic myeloid leukemia|9875/3
C0023473|T191|SY|0000007345|CHV|chronic myeloid leukemias|9875/3
C0023473|T191|SY|0000007345|CHV|cml|9875/3
C0023473|T191|PT|U000138|COSTAR|CHRONIC GRANULOCYTIC LEUKEMIA|9875/3
C0023473|T191|ET|2004-1700|CSP|chronic granulocytic leukemia|9875/3
C0023473|T191|ET|2004-1700|CSP|chronic myelocytic leukemia|9875/3
C0023473|T191|PT|2004-1700|CSP|chronic myelogenous leukemia|9875/3
C0023473|T191|ET|2004-1700|CSP|chronic myeloid leukemia|9875/3
C0023473|T191|ET|2004-1700|CSP|CML|9875/3
C0023473|T191|PT|LEUKEMIA CHRON MYELO|CST|CHRONIC MYELOCYTIC LEUKEMIA|9875/3
C0023473|T191|GT|LEUKEMIA CHRON MYELO|CST|LEUKEMIA MYELOCYTIC CHRONIC|9875/3
C0023473|T191|SY|NOCODE|DXP|CML|9875/3
C0023473|T191|SY|NOCODE|DXP|LEUKEMIA, GRANULOCYTIC, CHRONIC|9875/3
C0023473|T191|DI|U001052|DXP|LEUKEMIA, MYELOCYTIC, CHRONIC|9875/3
C0023473|T191|SY|NOCODE|DXP|LEUKEMIA, MYELOGENOUS, CHRONIC|9875/3
C0023473|T191|SY|NOCODE|DXP|LEUKEMIA, MYELOID, CHRONIC|9875/3
C0023473|T191|SY|HP:0005506|HPO|Chronic myelocytic leukemia|9875/3
C0023473|T191|PT|HP:0005506|HPO|Chronic myelogenous leukemia|9875/3
C0023473|T191|SY|HP:0005506|HPO|Chronic myeloid leukemia|9875/3
C0023473|T191|PT|C92.1|ICD10|Chronic myeloid leukaemia|9875/3
C0023473|T191|PT|C92.1|ICD10AE|Chronic myeloid leukemia|9875/3
C0023473|T191|HT|205.1|ICD9CM|Myeloid leukemia, chronic|9875/3
C0023473|T191|PT|MTHU016669|ICPC2ICD10ENG|chronic; myelosis|9875/3
C0023473|T191|PT|MTHU032697|ICPC2ICD10ENG|granulocytic; leukemia, chronic|9875/3
C0023473|T191|PT|MTHU044757|ICPC2ICD10ENG|leukemia; granulocytic, chronic|9875/3
C0023473|T191|PT|MTHU044782|ICPC2ICD10ENG|leukemia; myelocytic, chronic|9875/3
C0023473|T191|PT|MTHU044786|ICPC2ICD10ENG|leukemia; myeloid, chronic|9875/3
C0023473|T191|PT|MTHU050843|ICPC2ICD10ENG|myelocytic; leukemia, chronic|9875/3
C0023473|T191|PT|MTHU050857|ICPC2ICD10ENG|myeloid; leukemia, chronic|9875/3
C0023473|T191|PT|MTHU050919|ICPC2ICD10ENG|myelosis; chronic|9875/3
C0023473|T191|PTN|B73005|ICPC2P|chronic myeloid leukaemia|9875/3
C0023473|T191|MTH_PTN|B73005|ICPC2P|chronic myeloid leukemia|9875/3
C0023473|T191|PT|B73005|ICPC2P|Leukaemia;chronic myeloid|9875/3
C0023473|T191|MTH_PT|B73005|ICPC2P|Leukemia;chronic myeloid|9875/3
C0023473|T191|PT|sh2004008307|LCH_NW|Chronic myeloid leukemia|9875/3
C0023473|T191|LA|LA26791-6|LNC|Chronic myelogenous leukemia|9875/3
C0023473|T191|LLT|10008904|MDR|Chronic granulocytic leukaemia|9875/3
C0023473|T191|LLT|10008905|MDR|Chronic granulocytic leukemia|9875/3
C0023473|T191|LLT|10058245|MDR|Chronic myelocytic leukaemia|9875/3
C0023473|T191|LLT|10009011|MDR|Chronic myelocytic leukemia|9875/3
C0023473|T191|LLT|10058246|MDR|Chronic myelogenous leukaemia|9875/3
C0023473|T191|LLT|10009012|MDR|Chronic myelogenous leukemia|9875/3
C0023473|T191|LLT|10009013|MDR|Chronic myeloid leukaemia|9875/3
C0023473|T191|PT|10009013|MDR|Chronic myeloid leukaemia|9875/3
C0023473|T191|LLT|10009015|MDR|Chronic myeloid leukemia|9875/3
C0023473|T191|MTH_PT|10009013|MDR|Chronic myeloid leukemia|9875/3
C0023473|T191|LLT|10009700|MDR|CML|9875/3
C0023473|T191|LLT|10058247|MDR|Leukaemia myelocytic chronic|9875/3
C0023473|T191|HT|10024296|MDR|Leukaemias chronic myeloid|9875/3
C0023473|T191|LLT|10024347|MDR|Leukemia myelocytic chronic|9875/3
C0023473|T191|MTH_HT|10024296|MDR|Leukemias chronic myeloid|9875/3
C0023473|T191|LLT|10028553|MDR|Myeloid leukaemia, chronic|9875/3
C0023473|T191|LLT|10028558|MDR|Myeloid leukemia, chronic|9875/3
C0023473|T191|PT|31475|MEDCIN|chronic myelogenous leukemia|9875/3
C1292771|T191|PT|230914|MEDCIN|chronic myelogenous leukemia - BCR/ABL positive|9875/3
C1292771|T191|SY|230914|MEDCIN|chronic myelogenous leukemia BCR/ABL positive|9875/3
C0023473|T191|ET|5624|MEDLINEPLUS|Chronic Granulocytic Leukemia|9875/3
C0023473|T191|SY|5624|MEDLINEPLUS|Chronic granulocytic leukemia|9875/3
C0023473|T191|ET|5624|MEDLINEPLUS|Chronic Myelogenous Leukemia|9875/3
C0023473|T191|SY|5624|MEDLINEPLUS|Chronic myelogenous leukemia|9875/3
C0023473|T191|PT|5624|MEDLINEPLUS|Chronic Myeloid Leukemia|9875/3
C0023473|T191|SY|5624|MEDLINEPLUS|CML|9875/3
C0023473|T191|ET|5624|MEDLINEPLUS|CML|9875/3
C0023473|T191|ET|5624|MEDLINEPLUS|Leukemia, Myeloid, Chronic|9875/3
C0023473|T191|PM|D015464|MSH|Chronic Granulocytic Leukemia|9875/3
C0023473|T191|PM|D015464|MSH|Chronic Granulocytic Leukemias|9875/3
C0023473|T191|PM|D015464|MSH|Chronic Myelocytic Leukemia|9875/3
C0023473|T191|PM|D015464|MSH|Chronic Myelocytic Leukemias|9875/3
C0023473|T191|PM|D015464|MSH|Chronic Myelogenous Leukemia|9875/3
C0023473|T191|PM|D015464|MSH|Chronic Myelogenous Leukemias|9875/3
C0023473|T191|PM|D015464|MSH|Chronic Myeloid Leukemia|9875/3
C0023473|T191|PM|D015464|MSH|Chronic Myeloid Leukemias|9875/3
C0023473|T191|ET|D015464|MSH|Granulocytic Leukemia, Chronic|9875/3
C0023473|T191|PM|D015464|MSH|Granulocytic Leukemias, Chronic|9875/3
C0023473|T191|DEV|D015464|MSH|LEUKEMIA PHILA POS|9875/3
C0023473|T191|PM|D015464|MSH|Leukemia, Chronic Granulocytic|9875/3
C0023473|T191|PM|D015464|MSH|Leukemia, Chronic Myelocytic|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Chronic Myelogenous|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Chronic Myeloid|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Granulocytic, Chronic|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myelocytic, Chronic|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myelogenous, Chronic|9875/3
C0023473|T191|MH|D015464|MSH|Leukemia, Myelogenous, Chronic, BCR-ABL Positive|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myelogenous, Ph1 Positive|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myelogenous, Ph1-Positive|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Chronic|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Ph1 Positive|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Ph1-Positive|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Philadelphia Positive|9875/3
C0023473|T191|ET|D015464|MSH|Leukemia, Myeloid, Philadelphia-Positive|9875/3
C0023473|T191|PM|D015464|MSH|Leukemia, Ph1-Positive Myelogenous|9875/3
C0023473|T191|PM|D015464|MSH|Leukemia, Ph1-Positive Myeloid|9875/3
C0023473|T191|PM|D015464|MSH|Leukemia, Philadelphia-Positive Myeloid|9875/3
C0023473|T191|PM|D015464|MSH|Leukemias, Chronic Granulocytic|9875/3
C0023473|T191|PM|D015464|MSH|Leukemias, Chronic Myelocytic|9875/3
C0023473|T191|PM|D015464|MSH|Leukemias, Chronic Myelogenous|9875/3
C0023473|T191|PM|D015464|MSH|Leukemias, Chronic Myeloid|9875/3
C0023473|T191|PM|D015464|MSH|Leukemias, Ph1-Positive Myelogenous|9875/3
C0023473|T191|PM|D015464|MSH|Leukemias, Ph1-Positive Myeloid|9875/3
C0023473|T191|PM|D015464|MSH|Leukemias, Philadelphia-Positive Myeloid|9875/3
C0023473|T191|ET|D015464|MSH|Myelocytic Leukemia, Chronic|9875/3
C0023473|T191|PM|D015464|MSH|Myelocytic Leukemias, Chronic|9875/3
C0023473|T191|ET|D015464|MSH|Myelogenous Leukemia, Chronic|9875/3
C0023473|T191|PM|D015464|MSH|Myelogenous Leukemia, Ph1 Positive|9875/3
C0023473|T191|ET|D015464|MSH|Myelogenous Leukemia, Ph1-Positive|9875/3
C0023473|T191|PM|D015464|MSH|Myelogenous Leukemias, Chronic|9875/3
C0023473|T191|PM|D015464|MSH|Myelogenous Leukemias, Ph1-Positive|9875/3
C0023473|T191|ET|D015464|MSH|Myeloid Leukemia, Chronic|9875/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemia, Ph1 Positive|9875/3
C0023473|T191|ET|D015464|MSH|Myeloid Leukemia, Ph1-Positive|9875/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemia, Philadelphia Positive|9875/3
C0023473|T191|ET|D015464|MSH|Myeloid Leukemia, Philadelphia-Positive|9875/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemias, Chronic|9875/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemias, Ph1-Positive|9875/3
C0023473|T191|PM|D015464|MSH|Myeloid Leukemias, Philadelphia-Positive|9875/3
C0023473|T191|PM|D015464|MSH|Ph1-Positive Myelogenous Leukemia|9875/3
C0023473|T191|PM|D015464|MSH|Ph1-Positive Myelogenous Leukemias|9875/3
C0023473|T191|PM|D015464|MSH|Ph1-Positive Myeloid Leukemia|9875/3
C0023473|T191|PM|D015464|MSH|Ph1-Positive Myeloid Leukemias|9875/3
C0023473|T191|PM|D015464|MSH|Philadelphia-Positive Myeloid Leukemia|9875/3
C0023473|T191|PM|D015464|MSH|Philadelphia-Positive Myeloid Leukemias|9875/3
C0023473|T191|PN|NOCODE|MTH|Myeloid Leukemia, Chronic|9875/3
C0023473|T191|SY|C3174|NCI|BCR-ABL Positive Chronic Myelogenous Leukemia|9875/3
C0023473|T191|SY|C3174|NCI|Chronic Granulocytic Leukemia|9875/3
C0023473|T191|SY|C3174|NCI|Chronic Myelocytic Leukemia|9875/3
C0023473|T191|SY|C3174|NCI|Chronic Myelogenous Leukemia|9875/3
C0023473|T191|SY|TCGA|NCI|Chronic Myelogenous Leukemia, BCR-ABL1 Positive|9875/3
C0023473|T191|PT|C3174|NCI|Chronic Myelogenous Leukemia, BCR-ABL1 Positive|9875/3
C0023473|T191|SY|C3174|NCI|Chronic Myelogenous Leukemias|9875/3
C0023473|T191|SY|C3174|NCI|Chronic Myeloid Leukemia|9875/3
C0023473|T191|AB|C3174|NCI|CML|9875/3
C0023473|T191|SY|C3174|NCI|CML - Chronic Myelogenous Leukemia|9875/3
C0023473|T191|PT|C3174|NCI_CPTAC|Chronic Myelogenous Leukemia, BCR-ABL1 Positive|9875/3
C0023473|T191|SY|C3174|NCI_CTRP|Chronic Myelogenous Leukemia, BCR-ABL1 Positive|9875/3
C0023473|T191|PT|CDR0000046754|NCI_NCI-GLOSS|chronic granulocytic leukemia|9875/3
C0023473|T191|PT|CDR0000044901|NCI_NCI-GLOSS|chronic myelogenous leukemia|9875/3
C0023473|T191|PT|CDR0000046755|NCI_NCI-GLOSS|chronic myeloid leukemia|9875/3
C0023473|T191|PT|CDR0000044382|NCI_NCI-GLOSS|CML|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|CGL|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|chronic granulocytic leukemia|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|chronic myelocytic leukemia|9875/3
C0023473|T191|PT|CDR0000037900|PDQ|chronic myelogenous leukemia|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|Chronic Myelogenous Leukemias|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|Chronic Myeloid Leukemia|9875/3
C0023473|T191|AB|CDR0000037900|PDQ|CML|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|CML - Chronic Myelogenous Leukemia|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|granulocytic leukemia, chronic|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|leukemia, chronic myelogenous|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|myelocytic leukemia, chronic|9875/3
C0023473|T191|SY|CDR0000037900|PDQ|myelogenous leukemia, chronic|9875/3
C0023473|T191|PT|R0121663|QMR|LEUKEMIA CHRONIC MYELOCYTIC|9875/3
C0023473|T191|AB|B651.|RCD|CGL - Chronic granul leukaemia|9875/3
C0023473|T191|SY|B651.|RCD|CGL - Chronic granulocytic leukaemia|9875/3
C0023473|T191|SY|B651.|RCD|Chronic granulocytic leukaemia|9875/3
C0023473|T191|PT|B651.|RCD|Chronic myeloid leukaemia|9875/3
C0023473|T191|OP|B651z|RCD|Chronic myeloid leukaemia NOS|9875/3
C0023473|T191|AB|B651.|RCD|CML - Chronic myeloid leukaem|9875/3
C0023473|T191|SY|B651.|RCD|CML - Chronic myeloid leukaemia|9875/3
C0023473|T191|AB|B651.|RCDAE|CGL - Chronic granul leukemia|9875/3
C0023473|T191|SY|B651.|RCDAE|CGL - Chronic granulocytic leukemia|9875/3
C0023473|T191|SY|B651.|RCDAE|Chronic granulocytic leukemia|9875/3
C0023473|T191|PT|B651.|RCDAE|Chronic myeloid leukemia|9875/3
C0023473|T191|OP|B651z|RCDAE|Chronic myeloid leukemia NOS|9875/3
C0023473|T191|SY|B651.|RCDAE|CML - Chronic myeloid leukemia|9875/3
C0023473|T191|OP|BBr63|RCDSA|Chronic myeloid leukemia|9875/3
C0023473|T191|OP|BBr63|RCDSY|Chronic myeloid leukaemia|9875/3
C0023473|T191|SYGB|92818009|SNOMEDCT_US|CGL - Chronic granulocytic leukaemia|9875/3
C0023473|T191|SY|92818009|SNOMEDCT_US|CGL - Chronic granulocytic leukemia|9875/3
C0023473|T191|SYGB|63364005|SNOMEDCT_US|Chronic granulocytic leukaemia|9875/3
C1292771|T191|SYGB|128825002|SNOMEDCT_US|Chronic granulocytic leukaemia, BCR/ABL|9875/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic granulocytic leukemia|9875/3
C1292771|T191|SY|128825002|SNOMEDCT_US|Chronic granulocytic leukemia, BCR/ABL|9875/3
C0023473|T191|SYGB|92818009|SNOMEDCT_US|Chronic myelocytic leukaemia|9875/3
C0023473|T191|SYGB|63364005|SNOMEDCT_US|Chronic myelocytic leukaemia|9875/3
C0023473|T191|SY|92818009|SNOMEDCT_US|Chronic myelocytic leukemia|9875/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic myelocytic leukemia|9875/3
C0023473|T191|SYGB|63364005|SNOMEDCT_US|Chronic myelogenous leukaemia|9875/3
C1292771|T191|PTGB|128825002|SNOMEDCT_US|Chronic myelogenous leukaemia, BCR/ABL positive|9875/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic myelogenous leukemia|9875/3
C1292771|T191|PT|128825002|SNOMEDCT_US|Chronic myelogenous leukemia, BCR/ABL positive|9875/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic myelogenous leukemia, no ICD-O subtype|9875/3
C0023473|T191|SY|63364005|SNOMEDCT_US|Chronic myelogenous leukemia, no International Classification of Diseases for Oncology subtype|9875/3
C0023473|T191|PTGB|92818009|SNOMEDCT_US|Chronic myeloid leukaemia|9875/3
C0023473|T191|PTGB|63364005|SNOMEDCT_US|Chronic myeloid leukaemia|9875/3
C0023473|T191|OAP|154592009|SNOMEDCT_US|Chronic myeloid leukaemia|9875/3
C0023473|T191|OF|154592009|SNOMEDCT_US|Chronic myeloid leukaemia|9875/3
C0023473|T191|OAP|188735005|SNOMEDCT_US|Chronic myeloid leukaemia NOS|9875/3
C0023473|T191|SYGB|92818009|SNOMEDCT_US|Chronic myeloid leukaemia, disease|9875/3
C0023473|T191|PT|92818009|SNOMEDCT_US|Chronic myeloid leukemia|9875/3
C0023473|T191|PT|63364005|SNOMEDCT_US|Chronic myeloid leukemia|9875/3
C0023473|T191|OAP|154592009|SNOMEDCT_US|Chronic myeloid leukemia|9875/3
C0023473|T191|OAP|188735005|SNOMEDCT_US|Chronic myeloid leukemia NOS|9875/3
C0023473|T191|SY|92818009|SNOMEDCT_US|Chronic myeloid leukemia, disease|9875/3
C0023473|T191|SYGB|92818009|SNOMEDCT_US|CML - Chronic myeloid leukaemia|9875/3
C0023473|T191|SY|92818009|SNOMEDCT_US|CML - Chronic myeloid leukemia|9875/3
C1292772|T191|PT|C92.2|ICD10|Subacute myeloid leukaemia|9876/3
C1292772|T191|PT|C92.2|ICD10AE|Subacute myeloid leukemia|9876/3
C1292772|T191|AB|C92.2|ICD10CM|Atypical chronic myeloid leukemia, BCR/ABL-negative|9876/3
C1292772|T191|HT|C92.2|ICD10CM|Atypical chronic myeloid leukemia, BCR/ABL-negative|9876/3
C1292772|T191|ET|C92.20|ICD10CM|Atypical chronic myeloid leukemia, BCR/ABL-negative NOS|9876/3
C1292772|T191|HT|205.2|ICD9CM|Myeloid leukemia, subacute|9876/3
C1292772|T191|PT|MTHU032698|ICPC2ICD10ENG|granulocytic; leukemia, subacute|9876/3
C1292772|T191|PT|MTHU044758|ICPC2ICD10ENG|leukemia; granulocytic, subacute|9876/3
C1292772|T191|PT|MTHU044787|ICPC2ICD10ENG|leukemia; myeloid, subacute|9876/3
C1292772|T191|PT|MTHU050858|ICPC2ICD10ENG|myeloid; leukemia, subacute|9876/3
C1292772|T191|PT|MTHU050924|ICPC2ICD10ENG|myelosis; subacute|9876/3
C1292772|T191|PT|MTHU071162|ICPC2ICD10ENG|subacute; myelosis|9876/3
C1292772|T191|LLT|10028554|MDR|Myeloid leukaemia, subacute|9876/3
C1292772|T191|LLT|10028559|MDR|Myeloid leukemia, subacute|9876/3
C1292772|T191|LLT|10042292|MDR|Subacute myeloid leukaemia|9876/3
C1292772|T191|LLT|10054651|MDR|Subacute myeloid leukemia|9876/3
C1292772|T191|PT|350015|MEDCIN|Atypical chronic myeloid leukemia|9876/3
C1292772|T191|SY|99746|MEDCIN|leukemia myelogenous subacute|9876/3
C1292772|T191|PT|99746|MEDCIN|subacute myelogenous leukemia|9876/3
C1292772|T191|ET|D054438|MSH|Atypical Chronic Myeloid Leukemia|9876/3
C1292772|T191|ET|D054438|MSH|Chronic Myeloid Leukemia, Atypical|9876/3
C1292772|T191|DEV|D054438|MSH|LEUKEMIA PHILA NEG|9876/3
C1292772|T191|ET|D054438|MSH|Leukemia, Myelogenous, Ph1 Negative|9876/3
C1292772|T191|ET|D054438|MSH|Leukemia, Myelogenous, Ph1-Negative|9876/3
C1292772|T191|ET|D054438|MSH|Leukemia, Myeloid, Chronic, Atypical|9876/3
C1292772|T191|MH|D054438|MSH|Leukemia, Myeloid, Chronic, Atypical, BCR-ABL Negative|9876/3
C1292772|T191|ET|D054438|MSH|Leukemia, Myeloid, Ph1 Negative|9876/3
C1292772|T191|ET|D054438|MSH|Leukemia, Myeloid, Ph1-Negative|9876/3
C1292772|T191|ET|D054438|MSH|Leukemia, Myeloid, Philadelphia Negative|9876/3
C1292772|T191|ET|D054438|MSH|Leukemia, Myeloid, Philadelphia-Negative|9876/3
C1292772|T191|PM|D054438|MSH|Leukemia, Ph1-Negative Myelogenous|9876/3
C1292772|T191|PM|D054438|MSH|Leukemia, Ph1-Negative Myeloid|9876/3
C1292772|T191|PM|D054438|MSH|Leukemia, Philadelphia-Negative Myeloid|9876/3
C1292772|T191|PM|D054438|MSH|Leukemias, Ph1-Negative Myelogenous|9876/3
C1292772|T191|PM|D054438|MSH|Leukemias, Ph1-Negative Myeloid|9876/3
C1292772|T191|PM|D054438|MSH|Leukemias, Philadelphia-Negative Myeloid|9876/3
C1292772|T191|PM|D054438|MSH|Myelogenous Leukemia, Ph1 Negative|9876/3
C1292772|T191|ET|D054438|MSH|Myelogenous Leukemia, Ph1-Negative|9876/3
C1292772|T191|PM|D054438|MSH|Myelogenous Leukemias, Ph1-Negative|9876/3
C1292772|T191|PM|D054438|MSH|Myeloid Leukemia, Ph1 Negative|9876/3
C1292772|T191|ET|D054438|MSH|Myeloid Leukemia, Ph1-Negative|9876/3
C1292772|T191|PM|D054438|MSH|Myeloid Leukemia, Philadelphia Negative|9876/3
C1292772|T191|ET|D054438|MSH|Myeloid Leukemia, Philadelphia-Negative|9876/3
C1292772|T191|PM|D054438|MSH|Myeloid Leukemias, Ph1-Negative|9876/3
C1292772|T191|PM|D054438|MSH|Myeloid Leukemias, Philadelphia-Negative|9876/3
C1292772|T191|PM|D054438|MSH|Ph1-Negative Myelogenous Leukemia|9876/3
C1292772|T191|PM|D054438|MSH|Ph1-Negative Myelogenous Leukemias|9876/3
C1292772|T191|PM|D054438|MSH|Ph1-Negative Myeloid Leukemia|9876/3
C1292772|T191|PM|D054438|MSH|Ph1-Negative Myeloid Leukemias|9876/3
C1292772|T191|PM|D054438|MSH|Philadelphia-Negative Myeloid Leukemia|9876/3
C1292772|T191|PM|D054438|MSH|Philadelphia-Negative Myeloid Leukemias|9876/3
C1292772|T191|PN|NOCODE|MTH|Leukemia, Myeloid, Chronic, Atypical, BCR-ABL Negative|9876/3
C1292772|T191|AB|C3519|NCI|aCML|9876/3
C1292772|T191|SY|C3519|NCI|Atypical Chronic Myeloid Leukemia|9876/3
C1292772|T191|PT|C3519|NCI|Atypical Chronic Myeloid Leukemia, BCR-ABL1 Negative|9876/3
C1292772|T191|SY|TCGA|NCI|Atypical Chronic Myeloid Leukemia, BCR-ABL1 Negative|9876/3
C1292772|T191|SY|C3519|NCI|Atypical CML|9876/3
C1292772|T191|PT|C3176|NCI|Philadelphia-Negative Myelogenous Leukemia|9876/3
C1292772|T191|OP|C3519|NCI|Subacute Granulocytic Leukemia|9876/3
C1292772|T191|OP|C3519|NCI|Subacute Myelogenous Leukemia|9876/3
C1292772|T191|SY|C3519|NCI|Subacute Myeloid Leukemia|9876/3
C1292772|T191|DN|C3519|NCI_CTRP|Atypical Chronic Myeloid Leukemia, BCR-ABL1 Negative|9876/3
C1292772|T191|AB|CDR0000335175|PDQ|aCML|9876/3
C1292772|T191|SY|CDR0000335175|PDQ|atypical chronic myeloid leukemia|9876/3
C1292772|T191|PT|CDR0000335175|PDQ|atypical chronic myeloid leukemia, BCR-ABL1 negative|9876/3
C1292772|T191|AB|CDR0000335175|PDQ|atypical CML|9876/3
C1292772|T191|IS|CDR0000335175|PDQ|subacute granulocytic leukemia|9876/3
C1292772|T191|IS|CDR0000335175|PDQ|subacute myelogenous leukemia|9876/3
C1292772|T191|SY|CDR0000335175|PDQ|subacute myeloid leukemia|9876/3
C1292772|T191|AB|Xa0SX|RCD|Atypic chron myeloid leukaemia|9876/3
C1292772|T191|PT|Xa0SX|RCD|Atypical chronic myeloid leukaemia|9876/3
C1292772|T191|PT|B652.|RCD|Subacute myeloid leukaemia|9876/3
C1292772|T191|AB|Xa0SX|RCDAE|Atypic chron myeloid leukemia|9876/3
C1292772|T191|PT|Xa0SX|RCDAE|Atypical chronic myeloid leukemia|9876/3
C1292772|T191|PT|B652.|RCDAE|Subacute myeloid leukemia|9876/3
C1292772|T191|PT|BBr62|RCDSA|Subacute myeloid leukemia|9876/3
C1292772|T191|PT|BBr62|RCDSY|Subacute myeloid leukaemia|9876/3
C1292772|T191|PTGB|277589003|SNOMEDCT_US|Atypical chronic myeloid leukaemia|9876/3
C1292772|T191|PTGB|128826001|SNOMEDCT_US|Atypical chronic myeloid leukaemia, BCR/ABL negative|9876/3
C1292772|T191|PT|277589003|SNOMEDCT_US|Atypical chronic myeloid leukemia|9876/3
C1292772|T191|PT|128826001|SNOMEDCT_US|Atypical chronic myeloid leukemia, BCR/ABL negative|9876/3
C1292772|T191|IS|74326002|SNOMEDCT_US|Subacute granulocytic leukemia|9876/3
C1292772|T191|IS|74326002|SNOMEDCT_US|Subacute myelogenous leukemia|9876/3
C1292772|T191|PTGB|188736006|SNOMEDCT_US|Subacute myeloid leukaemia|9876/3
C1292772|T191|OAP|95278004|SNOMEDCT_US|Subacute myeloid leukaemia|9876/3
C1292772|T191|OAP|74326002|SNOMEDCT_US|Subacute myeloid leukaemia|9876/3
C1292772|T191|IS|74326002|SNOMEDCT_US|Subacute myeloid leukaemia -RETIRED-|9876/3
C1292772|T191|IS|95278004|SNOMEDCT_US|Subacute myeloid leukaemia -RETIRED-|9876/3
C1292772|T191|OAP|74326002|SNOMEDCT_US|Subacute myeloid leukemia|9876/3
C1292772|T191|OAP|95278004|SNOMEDCT_US|Subacute myeloid leukemia|9876/3
C1292772|T191|PT|188736006|SNOMEDCT_US|Subacute myeloid leukemia|9876/3
C1292772|T191|OF|74326002|SNOMEDCT_US|Subacute myeloid leukemia -RETIRED-|9876/3
C1292772|T191|IS|74326002|SNOMEDCT_US|Subacute myeloid leukemia -RETIRED-|9876/3
C1292772|T191|IS|95278004|SNOMEDCT_US|Subacute myeloid leukemia -RETIRED-|9876/3
C1292772|T191|OF|95278004|SNOMEDCT_US|Subacute myeloid leukemia -RETIRED-|9876/3
C0023465|T191|SY|0000007342|CHV|acute monoblastic leukemia|9891/3
C0023465|T191|SY|0000058163|CHV|acute monoblastic leukemia|9891/3
C0023465|T191|PT|0000058163|CHV|acute monocytic leukemia|9891/3
C0023465|T191|PT|0000007342|CHV|acute monocytic leukemia|9891/3
C0023465|T191|PT|2004-2820|CSP|acute monocytic leukemia|9891/3
C0023465|T191|PT|LEUKEMIA ACUTE MONO|CST|ACUTE MONOBLASTIC LEUKEMIA|9891/3
C0023465|T191|GT|LEUKEMIA ACUTE MONO|CST|LEUKEMIA MONOBLASTIC ACUTE|9891/3
C0023465|T191|DI|U001044|DXP|LEUKEMIA, ACUTE MONOCYTIC|9891/3
C0023465|T191|SY|HP:0004845|HPO|Acute monoblastic leukemia|9891/3
C0023465|T191|PT|HP:0004845|HPO|Acute monocytic leukemia|9891/3
C0023465|T191|SY|HP:0004845|HPO|AML-M5|9891/3
C0023465|T191|SY|HP:0004845|HPO|AMoL|9891/3
C3831784|T191|PT|C93.0|ICD10|Acute monocytic leukaemia|9891/3
C3831784|T191|PT|C93.0|ICD10AE|Acute monocytic leukemia|9891/3
C3831784|T191|AB|C93.0|ICD10CM|Acute monoblastic/monocytic leukemia|9891/3
C3831784|T191|HT|C93.0|ICD10CM|Acute monoblastic/monocytic leukemia|9891/3
C3831784|T191|ET|C93.00|ICD10CM|Acute monoblastic/monocytic leukemia NOS|9891/3
C3831784|T191|ET|C93.0|ICD10CM|AML M5|9891/3
C0023465|T191|HT|206.0|ICD9CM|Monocytic leukemia, acute|9891/3
C0023465|T191|PT|MTHU050292|ICPC2ICD10ENG|monocytic; leukemia, acute|9891/3
C0023465|T191|PT|10000871|MDR|Acute monocytic leukaemia|9891/3
C0023465|T191|LLT|10000871|MDR|Acute monocytic leukaemia|9891/3
C0023465|T191|LLT|10000873|MDR|Acute monocytic leukemia|9891/3
C0023465|T191|MTH_PT|10000871|MDR|Acute monocytic leukemia|9891/3
C0023465|T191|LLT|10027890|MDR|Monocytic leukaemia, acute|9891/3
C0023465|T191|LLT|10027895|MDR|Monocytic leukemia, acute|9891/3
C3831784|T191|PT|338571|MEDCIN|acute monoblastic/monocytic leukemia|9891/3
C0023465|T191|PT|97733|MEDCIN|acute monocytic leukemia|9891/3
C0023465|T191|SY|97733|MEDCIN|leukemia monocytic acute|9891/3
C3831784|T191|SY|338571|MEDCIN|leukemia monocytic/monoblastic acute|9891/3
C0023465|T191|PM|D007948|MSH|Acute Monoblastic Leukemia|9891/3
C0023465|T191|PM|D007948|MSH|Acute Monoblastic Leukemias|9891/3
C0023465|T191|PM|D007948|MSH|Acute Monocytic Leukemia|9891/3
C0023465|T191|PM|D007948|MSH|Acute Monocytic Leukemias|9891/3
C0023465|T191|DSV|D007948|MSH|LEUKEMIA MYELOID ACUTE M 05|9891/3
C0023465|T191|ET|D007948|MSH|Leukemia, Acute Monocytic|9891/3
C0023465|T191|ET|D007948|MSH|Leukemia, Monoblastic, Acute|9891/3
C0023465|T191|MH|D007948|MSH|Leukemia, Monocytic, Acute|9891/3
C0023465|T191|ET|D007948|MSH|Leukemia, Myeloid, Acute, M5|9891/3
C0023465|T191|ET|D007948|MSH|Leukemia, Myeloid, Schilling Type|9891/3
C0023465|T191|ET|D007948|MSH|Leukemia, Myeloid, Schilling-Type|9891/3
C0023465|T191|PM|D007948|MSH|Leukemia, Schilling-Type Myeloid|9891/3
C0023465|T191|PM|D007948|MSH|Leukemias, Acute Monoblastic|9891/3
C0023465|T191|PM|D007948|MSH|Leukemias, Acute Monocytic|9891/3
C0023465|T191|ET|D007948|MSH|Monoblastic Leukemia, Acute|9891/3
C0023465|T191|PM|D007948|MSH|Monoblastic Leukemias, Acute|9891/3
C0023465|T191|ET|D007948|MSH|Monocytic Leukemia, Acute|9891/3
C0023465|T191|PM|D007948|MSH|Monocytic Leukemias, Acute|9891/3
C0023465|T191|DSV|D007948|MSH|MYELOID LEUKEMIA ACUTE M 05|9891/3
C0023465|T191|ET|D007948|MSH|Myeloid Leukemia, Acute, M5|9891/3
C0023465|T191|PM|D007948|MSH|Myeloid Leukemia, Schilling Type|9891/3
C0023465|T191|ET|D007948|MSH|Myeloid Leukemia, Schilling-Type|9891/3
C0023465|T191|PM|D007948|MSH|Schilling-Type Myeloid Leukemia|9891/3
C0023465|T191|PN|NOCODE|MTH|Acute monocytic leukemia|9891/3
C3831784|T191|PN|NOCODE|MTH|Acute monocytic/monoblastic leukemia|9891/3
C1318544|T191|PN|NOCODE|MTH|M5b Acute differentiated monocytic leukemia|9891/3
C3831784|T191|PT|C7318|NCI|Acute Monoblastic and Monocytic Leukemia|9891/3
C3831784|T191|SY|TCGA|NCI|Acute Monoblastic and Monocytic Leukemia|9891/3
C3831784|T191|SY|C7318|NCI|Acute Monoblastic Leukemia and Acute Monocytic Leukemia|9891/3
C1318544|T191|PT|C4861|NCI|Acute Monocytic Leukemia|9891/3
C3831784|T191|SY|C7318|NCI|Acute Myeloid Leukemia M5|9891/3
C1318544|T191|SY|C4861|NCI|Monocytic Leukemia|9891/3
C1318544|T191|PT|C4861|NCI_CDISC|LEUKEMIA, MONOCYTIC, MALIGNANT|9891/3
C1318544|T191|SY|C4861|NCI_CDISC|Monocytic Leukemia|9891/3
C3831784|T191|PT|C7318|NCI_CPTAC|Acute Monoblastic and Monocytic Leukemia|9891/3
C1318544|T191|PT|C4861|NCI_CPTAC|Acute Monocytic Leukemia|9891/3
C3831784|T191|PT|C7318|NCI_NICHD|Acute Monoblastic and Monocytic Leukemia|9891/3
C0023465|T191|PT|Xa0Sl|RCD|Acute monoblastic leukaemia|9891/3
C0023465|T191|PT|B660.|RCD|Acute monocytic leukaemia|9891/3
C0023465|T191|SY|Xa0Sl|RCD|Acute monocytoid leukaemia|9891/3
C1318544|T191|AB|B660.|RCD|M5b - Acute monocytic leukaem|9891/3
C1318544|T191|SY|B660.|RCD|M5b - Acute monocytic leukaemia|9891/3
C0023465|T191|PT|Xa0Sl|RCDAE|Acute monoblastic leukemia|9891/3
C0023465|T191|PT|B660.|RCDAE|Acute monocytic leukemia|9891/3
C0023465|T191|SY|Xa0Sl|RCDAE|Acute monocytoid leukemia|9891/3
C1318544|T191|SY|B660.|RCDAE|M5b - Acute monocytic leukemia|9891/3
C0023465|T191|PT|BBr91|RCDSA|Acute monocytic leukemia|9891/3
C0023465|T191|PT|BBr91|RCDSY|Acute monocytic leukaemia|9891/3
C3831784|T191|PTGB|703818007|SNOMEDCT_US|Acute monoblastic and monocytic leukaemia|9891/3
C3831784|T191|PT|703818007|SNOMEDCT_US|Acute monoblastic and monocytic leukemia|9891/3
C0023465|T191|SYGB|22331004|SNOMEDCT_US|Acute monoblastic leukaemia|9891/3
C0023465|T191|SY|22331004|SNOMEDCT_US|Acute monoblastic leukemia|9891/3
C0023465|T191|PTGB|413441006|SNOMEDCT_US|Acute monocytic leukaemia|9891/3
C0023465|T191|PTGB|22331004|SNOMEDCT_US|Acute monocytic leukaemia|9891/3
C0023465|T191|OAS|91859000|SNOMEDCT_US|Acute monocytic leukaemia|9891/3
C0023465|T191|OAP|91859000|SNOMEDCT_US|Acute monocytic leukaemia, FAB M5|9891/3
C1318544|T191|SYGB|413441006|SNOMEDCT_US|Acute monocytic leukaemia, FAB M5b|9891/3
C1318544|T191|PT|413441006|SNOMEDCT_US|Acute monocytic leukemia|9891/3
C0023465|T191|OAS|91859000|SNOMEDCT_US|Acute monocytic leukemia|9891/3
C0023465|T191|PT|22331004|SNOMEDCT_US|Acute monocytic leukemia|9891/3
C0023465|T191|OAP|91859000|SNOMEDCT_US|Acute monocytic leukemia, FAB M5|9891/3
C1318544|T191|SY|413441006|SNOMEDCT_US|Acute monocytic leukemia, FAB M5b|9891/3
C0023465|T191|SY|22331004|SNOMEDCT_US|Acute monocytic leukemia, morphology|9891/3
C3831784|T191|PTGB|413442004|SNOMEDCT_US|Acute monocytic/monoblastic leukaemia|9891/3
C3831784|T191|PT|413442004|SNOMEDCT_US|Acute monocytic/monoblastic leukemia|9891/3
C0023465|T191|SY|22331004|SNOMEDCT_US|FAB M5|9891/3
C1318544|T191|SY|22331004|SNOMEDCT_US|FAB M5B|9891/3
C1318544|T191|OAS|91859000|SNOMEDCT_US|M5b - Acute monocytic leukaemia|9891/3
C1318544|T191|SYGB|413441006|SNOMEDCT_US|M5b - Acute monocytic leukaemia|9891/3
C1318544|T191|SY|413441006|SNOMEDCT_US|M5b - Acute monocytic leukemia|9891/3
C1318544|T191|OAS|91859000|SNOMEDCT_US|M5b - Acute monocytic leukemia|9891/3
C1292773|T191|AB|C92.A|ICD10CM|Acute myeloid leukemia with multilineage dysplasia|9895/3
C1292773|T191|HT|C92.A|ICD10CM|Acute myeloid leukemia with multilineage dysplasia|9895/3
C1292773|T191|ET|C92.A0|ICD10CM|Acute myeloid leukemia with multilineage dysplasia NOS|9895/3
C1292773|T191|PT|230922|MEDCIN|acute myelogenous leukemia with multilineage dysplasia|9895/3
C1292773|T191|SY|230922|MEDCIN|AML with multilineage dysplasia|9895/3
C1292773|T191|PN|NOCODE|MTH|Acute myeloid leukemia with multilineage dysplasia|9895/3
C2825139|T191|PN|NOCODE|MTH|Acute Myeloid Leukemia with Myelodysplasia-Related Changes|9895/3
C1292773|T191|SY|TCGA|NCI|Acute Myeloid Leukemia with Multilineage Dysplasia|9895/3
C1292773|T191|PT|C9289|NCI|Acute Myeloid Leukemia with Multilineage Dysplasia|9895/3
C2825139|T191|PT|C7600|NCI|Acute Myeloid Leukemia with Myelodysplasia-Related Changes|9895/3
C2825139|T191|SY|TCGA|NCI|Acute Myeloid Leukemia with Myelodysplasia-Related Changes|9895/3
C1292773|T191|SY|C9289|NCI|AML with Multilineage Dysplasia|9895/3
C2825139|T191|SY|C7600|NCI|AML with Myelodysplasia-Related Changes|9895/3
C1292773|T191|SY|C9289|NCI|De novo Acute Myeloid Leukemia with Multilineage Dysplasia|9895/3
C1292773|T191|PT|C9289|NCI_CPTAC|Acute Myeloid Leukemia with Multilineage Dysplasia|9895/3
C2825139|T191|PT|C7600|NCI_NICHD|Acute Myeloid Leukemia with Myelodysplasia-Related Changes|9895/3
C2825139|T191|SY|C7600|NCI_NICHD|AML with Myelodysplasia-Related Changes|9895/3
C1292773|T191|SYGB|128827005|SNOMEDCT_US|Acute myeloid leukaemia with multilineage dysplasia|9895/3
C1292773|T191|SYGB|445448008|SNOMEDCT_US|Acute myeloid leukaemia with multilineage dysplasia|9895/3
C1275662|T191|PTGB|397341000|SNOMEDCT_US|Acute myeloid leukaemia with multilineage dysplasia following a myelodysplastic syndrome or myelodysplastic syndrome/myeloproliferative disorder|9895/3
C1275663|T191|PTGB|397342007|SNOMEDCT_US|Acute myeloid leukaemia with multilineage dysplasia without antecedent myelodysplastic syndrome|9895/3
C2825139|T191|PTGB|128827005|SNOMEDCT_US|Acute myeloid leukaemia with myelodysplasia-related changes|9895/3
C2825139|T191|PTGB|445448008|SNOMEDCT_US|Acute myeloid leukaemia with myelodysplasia-related changes|9895/3
C2825139|T191|SYGB|128827005|SNOMEDCT_US|Acute myeloid leukaemia without prior myelodysplastic syndrome|9895/3
C1292773|T191|SY|445448008|SNOMEDCT_US|Acute myeloid leukemia with multilineage dysplasia|9895/3
C1292773|T191|SY|128827005|SNOMEDCT_US|Acute myeloid leukemia with multilineage dysplasia|9895/3
C1275662|T191|PT|397341000|SNOMEDCT_US|Acute myeloid leukemia with multilineage dysplasia following a myelodysplastic syndrome or myelodysplastic syndrome/myeloproliferative disorder|9895/3
C1275663|T191|PT|397342007|SNOMEDCT_US|Acute myeloid leukemia with multilineage dysplasia without antecedent myelodysplastic syndrome|9895/3
C2825139|T191|PT|128827005|SNOMEDCT_US|Acute myeloid leukemia with myelodysplasia-related changes|9895/3
C2825139|T191|PT|445448008|SNOMEDCT_US|Acute myeloid leukemia with myelodysplasia-related changes|9895/3
C2825139|T191|SY|128827005|SNOMEDCT_US|Acute myeloid leukemia without prior myelodysplastic syndrome|9895/3
C1275662|T191|SY|397341000|SNOMEDCT_US|AML with multilineage dysplasia following a myelodysplastic syndrome or myelodysplastic syndrome/myeloproliferative disorder|9895/3
C1275663|T191|SY|397342007|SNOMEDCT_US|AML with multilineage dysplasia without antecedent myelodysplastic syndrome|9895/3
C1292775|T191|AB|C92.6|ICD10CM|Acute myeloid leukemia with 11q23-abnormality|9897/3
C1292775|T191|HT|C92.6|ICD10CM|Acute myeloid leukemia with 11q23-abnormality|9897/3
C1292775|T191|ET|C92.60|ICD10CM|Acute myeloid leukemia with 11q23-abnormality NOS|9897/3
C1292775|T191|PN|NOCODE|MTH|Acute myeloid leukemia, 11q23 abnormalities|9897/3
C2919692|T191|SY|C82403|NCI|Acute Myeloid Leukemia with 11q23 Abnormalities|9897/3
C2919692|T191|SY|C82403|NCI|Acute Myeloid Leukemia with MLL Abnormalities|9897/3
C2825116|T191|PT|C6924|NCI|Acute Myeloid Leukemia with Variant MLL Translocations|9897/3
C2825116|T191|SY|TCGA|NCI|Acute Myeloid Leukemia with Variant MLL Translocations|9897/3
C2825116|T191|PT|C6924|NCI_NICHD|Acute Myeloid Leukemia with Variant MLL Translocations|9897/3
C2825116|T191|SY|C6924|NCI_NICHD|AML with Variant MLL Translocations|9897/3
C2919692|T191|SYGB|444911000|SNOMEDCT_US|Acute myeloid leukaemia with 11q23 abnormality|9897/3
C1292775|T191|PTGB|128829008|SNOMEDCT_US|Acute myeloid leukaemia, 11q23 abnormalities|9897/3
C1292775|T191|SYGB|128829008|SNOMEDCT_US|Acute myeloid leukaemia, MLL|9897/3
C2919692|T191|SY|444911000|SNOMEDCT_US|Acute myeloid leukemia with 11q23 abnormality|9897/3
C1292775|T191|PT|128829008|SNOMEDCT_US|Acute myeloid leukemia, 11q23 abnormalities|9897/3
C1292775|T191|SY|128829008|SNOMEDCT_US|Acute myeloid leukemia, MLL|9897/3
C1834582|T191|SY|HP:0005534|HPO|TMD|9898/1
C1834582|T191|SY|HP:0005534|HPO|Transient leukemia of Down syndrome|9898/1
C1834582|T191|SY|HP:0005534|HPO|Transient myeloproliferative disorder|9898/1
C1834582|T191|PT|HP:0005534|HPO|Transient myeloproliferative syndrome|9898/1
C1834582|T191|CE|C563551|MSH|Leukemia, Transient|9898/1
C1834582|T191|NM|C563551|MSH|Myeloproliferative Syndrome, Transient|9898/1
C1834582|T191|CE|C563551|MSH|Transient Abnormal Myelopoiesis|9898/1
C1834582|T191|PN|NOCODE|MTH|MYELOPROLIFERATIVE SYNDROME, TRANSIENT|9898/1
C1834582|T191|AB|C82339|NCI|TAM|9898/1
C1834582|T191|PT|C82339|NCI|Transient Abnormal Myelopoiesis Associated with Down Syndrome|9898/1
C1834582|T191|SY|C82339|NCI|Transient Myeloproliferative Disorder|9898/1
C1834582|T191|PT|C82339|NCI_NICHD|Transient Abnormal Myelopoiesis|9898/1
C1834582|T191|SY|C82339|NCI_NICHD|Transient Myeloproliferative Disorder|9898/1
C1834582|T191|PT|721307000|SNOMEDCT_US|Transient abnormal myelopoiesis|9898/1
C1834582|T191|PT|450934005|SNOMEDCT_US|Transient abnormal myelopoiesis|9898/1
C2825149|T191|PT|C43223|NCI|Myeloid Leukemia Associated with Down Syndrome|9898/3
C2825149|T191|PT|C43223|NCI_NICHD|Acute Myeloid Leukemia Occurring in Children with Down syndrome|9898/3
C2825149|T191|SY|C43223|NCI_NICHD|Acute Myeloid Leukemia with GATA1 Mutations|9898/3
C2825149|T191|SY|C43223|NCI_NICHD|AML Occurring in Children with Down Syndrome|9898/3
C2825149|T191|PTGB|450935006|SNOMEDCT_US|Myeloid leukaemia associated with Down Syndrome|9898/3
C2825149|T191|PT|450935006|SNOMEDCT_US|Myeloid leukemia associated with Down Syndrome|9898/3
C0023462|T191|SY|0000007341|CHV|acute megakaryoblastic leukemia|9910/3
C0023462|T191|PT|0000007341|CHV|acute megakaryocytic leukemia|9910/3
C0023462|T191|PT|0000058164|CHV|megakaryoblastic leukemia|9910/3
C0023462|T191|SY|0000058164|CHV|megakaryocytic leukemia|9910/3
C0023462|T191|SY|0000058164|CHV|megakaryocytic myelosis|9910/3
C0023462|T191|ET|0446-2826|CSP|megakaryocytic leukemia|9910/3
C0023462|T191|DI|U001049|DXP|LEUKEMIA, MEGAKARYOCYTIC|9910/3
C0023462|T191|PT|HP:0006733|HPO|Acute megakaryocytic leukemia|9910/3
C0023462|T191|SY|HP:0006733|HPO|AMegL|9910/3
C0023462|T191|PT|C94.2|ICD10|Acute megakaryoblastic leukaemia|9910/3
C0023462|T191|PT|C94.2|ICD10AE|Acute megakaryoblastic leukemia|9910/3
C0023462|T191|AB|C94.2|ICD10CM|Acute megakaryoblastic leukemia|9910/3
C0023462|T191|HT|C94.2|ICD10CM|Acute megakaryoblastic leukemia|9910/3
C0023462|T191|ET|C94.20|ICD10CM|Acute megakaryoblastic leukemia NOS|9910/3
C0023462|T191|ET|C94.2|ICD10CM|Acute megakaryocytic leukemia|9910/3
C0023462|T191|ET|C94.2|ICD10CM|Acute myeloid leukemia M7|9910/3
C0023462|T191|HT|207.2|ICD9CM|Megakaryocytic leukemia|9910/3
C0023462|T191|PT|MTHU044770|ICPC2ICD10ENG|leukemia; megakaryocytic|9910/3
C0023462|T191|PT|MTHU044802|ICPC2ICD10ENG|leukemia; thrombocytic|9910/3
C0023462|T191|PT|MTHU048035|ICPC2ICD10ENG|megakaryocytic; leukemia|9910/3
C0023462|T191|PT|MTHU048037|ICPC2ICD10ENG|megakaryocytic; myelosis|9910/3
C0023462|T191|PT|MTHU050922|ICPC2ICD10ENG|myelosis; megakaryocytic|9910/3
C0023462|T191|PT|MTHU075503|ICPC2ICD10ENG|thrombocytic; leukemia|9910/3
C0023462|T191|LLT|10000859|MDR|Acute megakaryoblastic leukaemia|9910/3
C0023462|T191|LLT|10060556|MDR|Acute megakaryoblastic leukemia|9910/3
C0023462|T191|LLT|10000860|MDR|Acute megakaryocytic leukaemia|9910/3
C0023462|T191|PT|10000860|MDR|Acute megakaryocytic leukaemia|9910/3
C0023462|T191|LLT|10000861|MDR|Acute megakaryocytic leukemia|9910/3
C0023462|T191|MTH_PT|10000860|MDR|Acute megakaryocytic leukemia|9910/3
C0023462|T191|LLT|10027121|MDR|Megakaryocytic leukaemia|9910/3
C0023462|T191|LLT|10027122|MDR|Megakaryocytic leukaemia NOS|9910/3
C0023462|T191|LLT|10027124|MDR|Megakaryocytic leukemia|9910/3
C0023462|T191|MTH_LLT|10027122|MDR|Megakaryocytic leukemia NOS|9910/3
C0023462|T191|PT|230925|MEDCIN|acute megakaryoblastic leukemia|9910/3
C0023462|T191|SY|230925|MEDCIN|leukemia acute megakaryoblastic|9910/3
C0023462|T191|SY|31479|MEDCIN|leukemia megakaryocytic|9910/3
C0023462|T191|PT|31479|MEDCIN|megakaryocytic leukemia|9910/3
C0023462|T191|PM|D007947|MSH|Acute Megakaryoblastic Leukemia|9910/3
C0023462|T191|PM|D007947|MSH|Acute Megakaryoblastic Leukemias|9910/3
C0023462|T191|PM|D007947|MSH|Acute Megakaryocytic Leukemia|9910/3
C0023462|T191|PM|D007947|MSH|Acute Megakaryocytic Leukemias|9910/3
C0023462|T191|DSV|D007947|MSH|LEUKEMIA MYELOID ACUTE M 07|9910/3
C0023462|T191|PM|D007947|MSH|Leukemia, Acute Megakaryoblastic|9910/3
C0023462|T191|PM|D007947|MSH|Leukemia, Acute Megakaryocytic|9910/3
C0023462|T191|MH|D007947|MSH|Leukemia, Megakaryoblastic, Acute|9910/3
C0023462|T191|ET|D007947|MSH|Leukemia, Megakaryocytic|9910/3
C0023462|T191|ET|D007947|MSH|Leukemia, Megakaryocytic, Acute|9910/3
C0023462|T191|ET|D007947|MSH|Leukemia, Myeloid, Acute, M7|9910/3
C0023462|T191|PM|D007947|MSH|Leukemias, Acute Megakaryoblastic|9910/3
C0023462|T191|PM|D007947|MSH|Leukemias, Acute Megakaryocytic|9910/3
C0023462|T191|PM|D007947|MSH|Leukemias, Megakaryocytic|9910/3
C0023462|T191|ET|D007947|MSH|Megakaryoblastic Leukemia, Acute|9910/3
C0023462|T191|PM|D007947|MSH|Megakaryoblastic Leukemias, Acute|9910/3
C0023462|T191|ET|D007947|MSH|Megakaryocytic Leukemia|9910/3
C0023462|T191|ET|D007947|MSH|Megakaryocytic Leukemia, Acute|9910/3
C0023462|T191|PM|D007947|MSH|Megakaryocytic Leukemias|9910/3
C0023462|T191|PM|D007947|MSH|Megakaryocytic Leukemias, Acute|9910/3
C0023462|T191|DSV|D007947|MSH|MYELOID LEUKEMIA ACUTE M 07|9910/3
C0023462|T191|ET|D007947|MSH|Myeloid Leukemia, Acute, M7|9910/3
C0023462|T191|PN|NOCODE|MTH|Acute Megakaryocytic Leukemias|9910/3
C0023462|T191|ET|207.2|MTHICD9|Megakaryocytic myelosis|9910/3
C0023462|T191|ET|207.2|MTHICD9|Thrombocytic leukemia|9910/3
C0023462|T191|SY|C3170|NCI|Acute M7 Myeloid Leukemia|9910/3
C0023462|T191|SY|TCGA|NCI|Acute Megakaryoblastic Leukemia|9910/3
C0023462|T191|PT|C3170|NCI|Acute Megakaryoblastic Leukemia|9910/3
C0023462|T191|SY|C3170|NCI|Acute Megakaryocytic Leukemia|9910/3
C0023462|T191|SY|C3170|NCI|FAB M7|9910/3
C0023462|T191|SY|C3170|NCI_CDISC|Acute M7 Myeloid Leukemia|9910/3
C0023462|T191|SY|C3170|NCI_CDISC|Acute Megakaryocytic Leukemia|9910/3
C0023462|T191|SY|C3170|NCI_CDISC|Fab M7|9910/3
C0023462|T191|PT|C3170|NCI_CDISC|LEUKEMIA, MEGAKARYOCYTIC, MALIGNANT|9910/3
C0023462|T191|PT|C3170|NCI_CPTAC|Acute Megakaryoblastic Leukemia|9910/3
C0023462|T191|PT|C3170|NCI_NICHD|Acute Megakaryoblastic Leukemia|9910/3
C0023462|T191|SY|C3170|NCI_NICHD|AMKL|9910/3
C0023462|T191|AB|Xa0Sm|RCD|Acute megakaryoblast leukaemia|9910/3
C0023462|T191|PT|Xa0Sm|RCD|Acute megakaryoblastic leukaemia|9910/3
C0023462|T191|SY|Xa0Sm|RCD|M7 - Acute megakaryoblastic leukaemia|9910/3
C0023462|T191|AB|Xa0Sm|RCD|M7-Acute megakaryoblas leukaem|9910/3
C0023462|T191|OP|B672.|RCD|Megakaryocytic leukaemia|9910/3
C0023462|T191|PT|BBrA2|RCD|Megakaryocytic myelosis|9910/3
C0023462|T191|IS|B672.|RCD|Thrombocytic leukaemia|9910/3
C0023462|T191|AB|Xa0Sm|RCDAE|Acute megakaryoblast leukemia|9910/3
C0023462|T191|PT|Xa0Sm|RCDAE|Acute megakaryoblastic leukemia|9910/3
C0023462|T191|SY|Xa0Sm|RCDAE|M7 - Acute megakaryoblastic leukemia|9910/3
C0023462|T191|OP|B672.|RCDAE|Megakaryocytic leukemia|9910/3
C0023462|T191|IS|B672.|RCDAE|Thrombocytic leukemia|9910/3
C0023462|T191|OP|BBrA5|RCDSA|Acute megakaryoblastic leukemia|9910/3
C0023462|T191|PT|BBrA1|RCDSA|Megakaryocytic leukemia|9910/3
C0023462|T191|SY|BBrA1|RCDSA|Thrombocytic leukemia|9910/3
C0023462|T191|OA|BBrA5|RCDSY|Acut megakaryoblast leukaem|9910/3
C0023462|T191|OP|BBrA5|RCDSY|Acute megakaryoblastic leukaemia|9910/3
C0023462|T191|PT|BBrA1|RCDSY|Megakaryocytic leukaemia|9910/3
C0023462|T191|SY|BBrA1|RCDSY|Thrombocytic leukaemia|9910/3
C0023462|T191|PTGB|52220008|SNOMEDCT_US|Acute megakaryoblastic leukaemia|9910/3
C0023462|T191|PTGB|277602003|SNOMEDCT_US|Acute megakaryoblastic leukaemia|9910/3
C0023462|T191|OAP|94149003|SNOMEDCT_US|Acute megakaryoblastic leukaemia, FAB M7|9910/3
C0023462|T191|SYGB|277602003|SNOMEDCT_US|Acute megakaryoblastic leukaemia, FAB M7|9910/3
C0023462|T191|SYGB|52220008|SNOMEDCT_US|Acute megakaryoblastic leukaemia, morphology|9910/3
C0023462|T191|PT|52220008|SNOMEDCT_US|Acute megakaryoblastic leukemia|9910/3
C0023462|T191|PT|277602003|SNOMEDCT_US|Acute megakaryoblastic leukemia|9910/3
C0023462|T191|SY|277602003|SNOMEDCT_US|Acute megakaryoblastic leukemia, FAB M7|9910/3
C0023462|T191|OAP|94149003|SNOMEDCT_US|Acute megakaryoblastic leukemia, FAB M7|9910/3
C0023462|T191|SY|52220008|SNOMEDCT_US|Acute megakaryoblastic leukemia, morphology|9910/3
C0023462|T191|SY|52220008|SNOMEDCT_US|FAB M7|9910/3
C0023462|T191|SYGB|277602003|SNOMEDCT_US|M7 - Acute megakaryoblastic leukaemia|9910/3
C0023462|T191|SY|277602003|SNOMEDCT_US|M7 - Acute megakaryoblastic leukemia|9910/3
C0023462|T191|SY|52220008|SNOMEDCT_US|Malignant megakaryocytosis|9910/3
C0023462|T191|SYGB|52220008|SNOMEDCT_US|Megakaryoblastic leukaemia|9910/3
C0023462|T191|SY|52220008|SNOMEDCT_US|Megakaryoblastic leukemia|9910/3
C0023462|T191|PTGB|188754005|SNOMEDCT_US|Megakaryocytic leukaemia|9910/3
C0023462|T191|SYGB|52220008|SNOMEDCT_US|Megakaryocytic leukaemia|9910/3
C0023462|T191|IS|277602003|SNOMEDCT_US|Megakaryocytic leukaemia|9910/3
C0023462|T191|OAS|94149003|SNOMEDCT_US|Megakaryocytic leukaemia|9910/3
C0023462|T191|OAS|94149003|SNOMEDCT_US|Megakaryocytic leukemia|9910/3
C0023462|T191|PT|188754005|SNOMEDCT_US|Megakaryocytic leukemia|9910/3
C0023462|T191|SY|52220008|SNOMEDCT_US|Megakaryocytic leukemia|9910/3
C0023462|T191|IS|277602003|SNOMEDCT_US|Megakaryocytic leukemia|9910/3
C0023462|T191|SY|52220008|SNOMEDCT_US|Megakaryocytic myelosis|9910/3
C0023462|T191|SYGB|188754005|SNOMEDCT_US|Thrombocytic leukaemia|9910/3
C0023462|T191|SY|188754005|SNOMEDCT_US|Thrombocytic leukemia|9910/3
C1336735|T191|LLT|10066355|MDR|Treatment related acute myeloid leukaemia|9920/3
C1336735|T191|LLT|10066353|MDR|Treatment related acute myeloid leukemia|9920/3
C1292776|T191|SY|366677|MEDCIN|acute therapy related myeloid leukemia and myelodysplastic syndrome|9920/3
C1292776|T191|PT|366677|MEDCIN|Therapy related acute myeloid leukemia and myelodysplastic syndrome|9920/3
C1292776|T191|SY|C27912|NCI|Acute Myeloid Leukaemias and Myelodysplastic Syndromes, Therapy-Related|9920/3
C1336735|T191|AB|C8252|NCI|t-AML|9920/3
C1336735|T191|PT|C8252|NCI|Therapy-Related Acute Myeloid Leukemia|9920/3
C1292776|T191|SY|C27912|NCI|Therapy-Related Acute Myeloid Leukemia and Myelodysplastic Syndrome|9920/3
C1292776|T191|SY|C27912|NCI|Therapy-Related AML and MDS|9920/3
C1292776|T191|SY|TCGA|NCI|Therapy-Related Myeloid Neoplasm|9920/3
C1292776|T191|PT|C27912|NCI|Therapy-Related Myeloid Neoplasm|9920/3
C1336735|T191|SY|C8252|NCI|Treatment Related Acute Myelocytic Leukemia|9920/3
C1336735|T191|SY|C8252|NCI|Treatment Related Acute Myelogenous Leukemia|9920/3
C1336735|T191|SY|C8252|NCI|Treatment Related Acute Myeloid Leukemia|9920/3
C1336735|T191|SY|C8252|NCI|Treatment Related AML|9920/3
C1336735|T191|SY|C8252|NCI|Treatment-Related Acute Myelocytic Leukemia|9920/3
C1336735|T191|SY|C8252|NCI|Treatment-Related Acute Myelogenous Leukemia|9920/3
C1336735|T191|SY|C8252|NCI|Treatment-related Acute Myeloid Leukemia|9920/3
C1336735|T191|SY|C8252|NCI|Treatment-Related AML|9920/3
C1336735|T191|PT|10066353|NCI_CTEP-SDC|Treatment related acute myeloid leukemia|9920/3
C1336735|T191|SY|10066353|NCI_CTEP-SDC|Treatment related AML|9920/3
C1336735|T191|DN|C8252|NCI_CTRP|High-Grade Treatment-Related Myeloid Neoplasm|9920/3
C1292776|T191|PT|C27912|NCI_NICHD|Therapy-Related Myeloid Neoplasm|9920/3
C1292776|T191|PTGB|721306009|SNOMEDCT_US|Therapy related acute myeloid leukaemia and myelodysplastic syndrome|9920/3
C1292776|T191|PT|721306009|SNOMEDCT_US|Therapy related acute myeloid leukemia and myelodysplastic syndrome|9920/3
C1292776|T191|PTGB|128830003|SNOMEDCT_US|Therapy-related acute myeloid leukaemia and myelodysplastic syndrome|9920/3
C1292776|T191|PT|128830003|SNOMEDCT_US|Therapy-related acute myeloid leukemia and myelodysplastic syndrome|9920/3
C4721505|T191|SY|0000017245|CHV|myeloid sarcoma|9930/3
C4721505|T191|SY|NOCODE|DXP|CANCER, GREEN|9930/3
C4721505|T191|SY|NOCODE|DXP|CHLOROLEUKEMIA|9930/3
C4721505|T191|DI|U000330|DXP|CHLOROMA|9930/3
C4721505|T191|SY|NOCODE|DXP|CHLOROMYELOMA|9930/3
C4721505|T191|SY|NOCODE|DXP|CHLOROSARCOMA|9930/3
C4721505|T191|PT|C92.3|ICD10|Myeloid sarcoma|9930/3
C4721505|T191|ET|C92.3|ICD10CM|Chloroma|9930/3
C4721505|T191|HT|C92.3|ICD10CM|Myeloid sarcoma|9930/3
C4721505|T191|AB|C92.3|ICD10CM|Myeloid sarcoma|9930/3
C4721505|T191|ET|C92.30|ICD10CM|Myeloid sarcoma NOS|9930/3
C4721505|T191|HT|205.3|ICD9CM|Myeloid sarcoma|9930/3
C4721505|T191|PT|MTHU016222|ICPC2ICD10ENG|chloroma|9930/3
C4721505|T191|PT|MTHU050859|ICPC2ICD10ENG|myeloid; sarcoma|9930/3
C4721505|T191|PT|MTHU050912|ICPC2ICD10ENG|myelosarcoma|9930/3
C4721505|T191|PT|MTHU065924|ICPC2ICD10ENG|sarcoma; myeloid|9930/3
C4721505|T191|PT|sh85024568|LCH_NW|Chloroma|9930/3
C4721505|T191|LLT|10008583|MDR|Chloroma|9930/3
C4721505|T191|PT|10008583|MDR|Chloroma|9930/3
C4721505|T191|LLT|10028562|MDR|Myeloid sarcoma|9930/3
C4721505|T191|PT|97882|MEDCIN|chloroma|9930/3
C4721505|T191|SY|97881|MEDCIN|leukemia myeloid sarcoma|9930/3
C4721505|T191|SY|97882|MEDCIN|leukemia myeloid sarcoma chloroma|9930/3
C4721505|T191|PT|97881|MEDCIN|myeloid sarcoma|9930/3
C4721505|T191|ET|D023981|MSH|Chloroma|9930/3
C4721505|T191|PM|D023981|MSH|Chloromas|9930/3
C4721505|T191|ET|D023981|MSH|Extramedullary Myeloid Cell Tumor|9930/3
C4721505|T191|ET|D023981|MSH|Myeloid Cell Tumor, Extramedullary|9930/3
C4721505|T191|ET|D023981|MSH|Myeloid Sarcoma|9930/3
C4721505|T191|PM|D023981|MSH|Myeloid Sarcomas|9930/3
C4721505|T191|MH|D023981|MSH|Sarcoma, Myeloid|9930/3
C4721505|T191|PM|D023981|MSH|Sarcomas, Myeloid|9930/3
C4721505|T191|PN|NOCODE|MTH|Sarcoma, Myeloid|9930/3
C4721505|T191|ET|205.3|MTHICD9|Chloroma|9930/3
C4721505|T191|SY|C3520|NCI|Chloroma|9930/3
C4721505|T191|SY|C3520|NCI|Extramedullary Myeloid Tumor|9930/3
C4721505|T191|PT|C3520|NCI|Myeloid Sarcoma|9930/3
C4721505|T191|SY|TCGA|NCI|Myeloid Sarcoma|9930/3
C4721505|T191|SY|C3520|NCI_CDISC|Chloroma|9930/3
C4721505|T191|SY|C3520|NCI_CDISC|Extramedullary Myeloid Tumor|9930/3
C4721505|T191|PT|C3520|NCI_CDISC|SARCOMA, MYELOID, MALIGNANT|9930/3
C4721505|T191|PT|C3520|NCI_CPTAC|Myeloid Sarcoma|9930/3
C4721505|T191|PT|CDR0000335063|NCI_NCI-GLOSS|chloroma|9930/3
C4721505|T191|PT|C3520|NCI_NICHD|Myeloid Sarcoma|9930/3
C4721505|T191|PT|B653.|RCD|Myeloid sarcoma|9930/3
C4721505|T191|OP|B653z|RCD|Myeloid sarcoma NOS|9930/3
C4721505|T191|OP|BBrA3|RCDSY|Myeloid sarcoma|9930/3
C4721505|T191|PT|188737002|SNOMEDCT_US|Chloroma|9930/3
C4721505|T191|SY|35287006|SNOMEDCT_US|Chloroma|9930/3
C4721505|T191|PT|35287006|SNOMEDCT_US|Myeloid sarcoma|9930/3
C4721505|T191|PT|94719007|SNOMEDCT_US|Myeloid sarcoma|9930/3
C4721505|T191|OAP|188739004|SNOMEDCT_US|Myeloid sarcoma NOS|9930/3
C4721505|T191|SY|94719007|SNOMEDCT_US|Myeloid sarcoma, disease|9930/3
C4721505|T191|SY|35287006|SNOMEDCT_US|Myeloid sarcoma, morphology|9930/3
C0334674|T191|PT|0000030020|CHV|acute myelofibrosis|9931/3
C0334674|T191|PT|C94.5|ICD10|Acute myelofibrosis|9931/3
C0334674|T191|PT|C94.4|ICD10|Acute panmyelosis|9931/3
C0334674|T191|ET|C94.4|ICD10CM|Acute myelofibrosis|9931/3
C0334674|T191|ET|C94.40|ICD10CM|Acute myelofibrosis NOS|9931/3
C0334674|T191|ET|C94.40|ICD10CM|Acute panmyelosis NOS|9931/3
C0334674|T191|AB|C94.4|ICD10CM|Acute panmyelosis with myelofibrosis|9931/3
C0334674|T191|HT|C94.4|ICD10CM|Acute panmyelosis with myelofibrosis|9931/3
C0334674|T191|PT|MTHU003165|ICPC2ICD10ENG|acute; myelofibrosis|9931/3
C0334674|T191|PT|MTHU050849|ICPC2ICD10ENG|myelofibrosis; acute|9931/3
C0334674|T191|LLT|10000879|MDR|Acute myelofibrosis|9931/3
C0334674|T191|PT|350342|MEDCIN|Acute myelofibrosis|9931/3
C0334674|T191|PT|311876|MEDCIN|acute panmyelosis|9931/3
C0334674|T191|PT|230928|MEDCIN|acute panmyelosis with myelofibrosis|9931/3
C0334674|T191|SY|350342|MEDCIN|myelofibrosis acute|9931/3
C0334674|T191|PN|NOCODE|MTH|Acute panmyelosis with myelofibrosis|9931/3
C0334674|T191|ET|238.7|MTHICD9|Acute panmyelosis|9931/3
C0334674|T191|SY|C4344|NCI|Acute Myelofibrosis|9931/3
C0334674|T191|SY|C4344|NCI|Acute Myelosclerosis|9931/3
C0334674|T191|SY|C4344|NCI|Acute Panmyelosis|9931/3
C0334674|T191|PT|C4344|NCI|Acute Panmyelosis with Myelofibrosis|9931/3
C0334674|T191|SY|TCGA|NCI|Acute Panmyelosis with Myelofibrosis|9931/3
C0334674|T191|AB|C4344|NCI|APMF|9931/3
C0334674|T191|PT|Xa0So|RCD|Acute myelofibrosis|9931/3
C0334674|T191|PT|B674.|RCD|Acute panmyelosis|9931/3
C0334674|T191|OP|BBrA7|RCDSY|Acute myelofibrosis|9931/3
C0334674|T191|PT|BBs1.|RCDSY|Acute panmyelosis|9931/3
C0334674|T191|OAP|21721006|SNOMEDCT_US|Acute myelofibrosis|9931/3
C0334674|T191|SY|80570006|SNOMEDCT_US|Acute myelofibrosis|9931/3
C0334674|T191|OAP|188757003|SNOMEDCT_US|Acute myelofibrosis|9931/3
C0334674|T191|SY|109991003|SNOMEDCT_US|Acute myelofibrosis|9931/3
C0334674|T191|OF|188757003|SNOMEDCT_US|Acute myelofibrosis|9931/3
C0334674|T191|OF|21721006|SNOMEDCT_US|Acute myelofibrosis -RETIRED-|9931/3
C0334674|T191|IS|21721006|SNOMEDCT_US|Acute myelofibrosis -RETIRED-|9931/3
C0334674|T191|SY|80570006|SNOMEDCT_US|Acute myelosclerosis|9931/3
C0334674|T191|OAP|188756007|SNOMEDCT_US|Acute panmyelosis|9931/3
C0334674|T191|SY|80570006|SNOMEDCT_US|Acute panmyelosis|9931/3
C0334674|T191|PT|80570006|SNOMEDCT_US|Acute panmyelosis with myelofibrosis|9931/3
C0334674|T191|PT|109991003|SNOMEDCT_US|Acute panmyelosis with myelofibrosis|9931/3
C0023443|T191|SD|NEO063|CCSR_10|Leukemia - hairy cell|9940/3
C0023443|T191|SY|0000007335|CHV|cell hairy leukemia|9940/3
C0023443|T191|SY|0000007335|CHV|cells hairy leukemia|9940/3
C0023443|T191|SY|0000007335|CHV|hairy cell leukaemia|9940/3
C0023443|T191|PT|0000007335|CHV|hairy cell leukemia|9940/3
C0023443|T191|SY|0000007335|CHV|hairy-cell leukaemia|9940/3
C0023443|T191|SY|0000007335|CHV|hairy-cell leukemia|9940/3
C0023443|T191|SY|0000007335|CHV|leukaemia hairy cell|9940/3
C0023443|T191|SY|0000007335|CHV|leukemia hairy cell|9940/3
C0023443|T191|PT|U000334|COSTAR|HAIRY CELL LEUKEMIA|9940/3
C0023443|T191|PT|2004-1799|CSP|hairy cell leukemia|9940/3
C0023443|T191|ET|2004-1799|CSP|hairy T cell leukemia|9940/3
C0023443|T191|SY|NOCODE|DXP|HAIRY CELL LEUKEMIA|9940/3
C0023443|T191|DI|U001666|DXP|RETICULOENDOTHELIOSIS, LEUKEMIC|9940/3
C0023443|T191|PT|C91.4|ICD10|Hairy-cell leukaemia|9940/3
C0023443|T191|PT|C91.4|ICD10AE|Hairy-cell leukemia|9940/3
C0023443|T191|HT|C91.4|ICD10CM|Hairy cell leukemia|9940/3
C0023443|T191|AB|C91.4|ICD10CM|Hairy cell leukemia|9940/3
C0023443|T191|ET|C91.40|ICD10CM|Hairy cell leukemia NOS|9940/3
C0023443|T191|ET|C91.4|ICD10CM|Leukemic reticuloendotheliosis|9940/3
C0023443|T191|HT|202.4|ICD9CM|Leukemic reticuloendotheliosis|9940/3
C0023443|T191|PT|MTHU044759|ICPC2ICD10ENG|leukemia; hairy cell|9940/3
C0023443|T191|PT|MTHU044803|ICPC2ICD10ENG|leukemic; reticuloendotheliosis|9940/3
C0023443|T191|PT|MTHU064351|ICPC2ICD10ENG|reticuloendotheliosis; leukemic|9940/3
C0023443|T191|PT|U002667|LCH|Leukemia, Hairy cell|9940/3
C0023443|T191|PT|sh85076294|LCH_NW|Leukemia, Hairy cell|9940/3
C0023443|T191|LLT|10019053|MDR|Hairy cell leukaemia|9940/3
C0023443|T191|PT|10019053|MDR|Hairy cell leukaemia|9940/3
C0023443|T191|LLT|10019055|MDR|Hairy cell leukemia|9940/3
C0023443|T191|MTH_PT|10019053|MDR|Hairy cell leukemia|9940/3
C0023443|T191|LLT|10024326|MDR|Leukaemic reticuloendotheliosis|9940/3
C0023443|T191|LLT|10024362|MDR|Leukemic reticuloendotheliosis|9940/3
C0023443|T191|PT|33858|MEDCIN|hairy cell leukemia|9940/3
C0023443|T191|SY|33858|MEDCIN|hairy-cell leukemia|9940/3
C0023443|T191|SY|33858|MEDCIN|leukemia hairy-cell|9940/3
C0023443|T191|ET|5620|MEDLINEPLUS|Hairy Cell Leukemia|9940/3
C0023443|T191|ET|D007943|MSH|Hairy Cell Leukemia|9940/3
C0023443|T191|PM|D007943|MSH|Hairy Cell Leukemias|9940/3
C0023443|T191|MH|D007943|MSH|Leukemia, Hairy Cell|9940/3
C0023443|T191|PM|D007943|MSH|Leukemias, Hairy Cell|9940/3
C0023443|T191|PM|D007943|MSH|Leukemic Reticuloendothelioses|9940/3
C0023443|T191|ET|D007943|MSH|Leukemic Reticuloendotheliosis|9940/3
C0023443|T191|PM|D007943|MSH|Reticuloendothelioses, Leukemic|9940/3
C0023443|T191|ET|D007943|MSH|Reticuloendotheliosis, Leukemic|9940/3
C0023443|T191|SY|NOCODE|MTH|HAIRY CELL LEUKEMIA|9940/3
C0023443|T191|PN|NOCODE|MTH|Hairy Cell Leukemia|9940/3
C0023443|T191|ET|202.4|MTHICD9|Hairy-cell leukemia|9940/3
C0023443|T191|SY|TCGA|NCI|Hairy Cell Leukemia|9940/3
C0023443|T191|PT|C7402|NCI|Hairy Cell Leukemia|9940/3
C0023443|T191|AB|C7402|NCI|HCL|9940/3
C0023443|T191|SY|C7402|NCI|Leukemic Reticuloendotheliosis|9940/3
C0023443|T191|PT|C7402|NCI_CPTAC|Hairy Cell Leukemia|9940/3
C0023443|T191|PT|10019053|NCI_CTEP-SDC|Hairy cell leukemia|9940/3
C0023443|T191|DN|C7402|NCI_CTRP|Hairy Cell Leukemia|9940/3
C0023443|T191|PT|CDR0000045159|NCI_NCI-GLOSS|hairy cell leukemia|9940/3
C0023443|T191|PT|CDR0000039065|PDQ|hairy cell leukemia|9940/3
C0023443|T191|AB|CDR0000039065|PDQ|HCL|9940/3
C0023443|T191|SY|CDR0000039065|PDQ|leukemia, hairy cell|9940/3
C0023443|T191|ET|CDR0000039065|PDQ|Leukemia, hairy cell|9940/3
C0023443|T191|SY|CDR0000039065|PDQ|Leukemic Reticuloendotheliosis|9940/3
C0023443|T191|PT|R0121664|QMR|LEUKEMIA HAIRY CELL|9940/3
C0023443|T191|PT|B624.|RCD|Hairy cell leukaemia|9940/3
C0023443|T191|SY|B624.|RCD|HCL - Hairy cell leukaemia|9940/3
C0023443|T191|AB|B624.|RCD|Leukaem reticuloendotheliosis|9940/3
C0023443|T191|OA|B6240|RCD|Leukaem.reticuloend.-unsp.site|9940/3
C0023443|T191|OA|B624z|RCD|Leukaemic reticuloendoth. NOS|9940/3
C0023443|T191|SY|B624.|RCD|Leukaemic reticuloendotheliosis|9940/3
C0023443|T191|OP|B624z|RCD|Leukaemic reticuloendotheliosis NOS|9940/3
C0023443|T191|OP|B6240|RCD|Leukaemic reticuloendotheliosis of unspecified sites|9940/3
C0023443|T191|SY|B624.|RCD|LRE - Leukaemic reticuloendotheliosis|9940/3
C0023443|T191|AB|B624.|RCD|LRE-Leuk reticuloendotheliosis|9940/3
C0023443|T191|PT|B624.|RCDAE|Hairy cell leukemia|9940/3
C0023443|T191|SY|B624.|RCDAE|HCL - Hairy cell leukemia|9940/3
C0023443|T191|OA|B624z|RCDAE|Leukemic reticuloendoth. NOS|9940/3
C0023443|T191|SY|B624.|RCDAE|Leukemic reticuloendotheliosis|9940/3
C0023443|T191|OP|B624z|RCDAE|Leukemic reticuloendotheliosis NOS|9940/3
C0023443|T191|OP|B6240|RCDAE|Leukemic reticuloendotheliosis of unspecified sites|9940/3
C0023443|T191|SY|B624.|RCDAE|LRE - Leukemic reticuloendotheliosis|9940/3
C0023443|T191|IS|BBrA8|RCDSA|Hairy cell leukemia|9940/3
C0023443|T191|OP|BBrA8|RCDSA|Leukemic reticuloendotheliosis|9940/3
C0023443|T191|IS|BBrA8|RCDSY|Hairy cell leukaemia|9940/3
C0023443|T191|OA|BBrA8|RCDSY|Leukaem reticuloendothelsis|9940/3
C0023443|T191|OP|BBrA8|RCDSY|Leukaemic reticuloendotheliosis|9940/3
C0023443|T191|PTGB|54087003|SNOMEDCT_US|Hairy cell leukaemia|9940/3
C0023443|T191|SYGB|118613001|SNOMEDCT_US|Hairy cell leukaemia|9940/3
C0023443|T191|PT|54087003|SNOMEDCT_US|Hairy cell leukemia|9940/3
C0023443|T191|SY|118613001|SNOMEDCT_US|Hairy cell leukemia|9940/3
C0023443|T191|SYGB|118613001|SNOMEDCT_US|HCL - Hairy cell leukaemia|9940/3
C0023443|T191|SY|118613001|SNOMEDCT_US|HCL - Hairy cell leukemia|9940/3
C0023443|T191|SYGB|54087003|SNOMEDCT_US|Leukaemic reticuloendotheliosis|9940/3
C0023443|T191|OAP|85228003|SNOMEDCT_US|Leukaemic reticuloendotheliosis|9940/3
C0023443|T191|IS|85228003|SNOMEDCT_US|Leukaemic reticuloendotheliosis -RETIRED-|9940/3
C0023443|T191|OAP|188653005|SNOMEDCT_US|Leukaemic reticuloendotheliosis NOS|9940/3
C0023443|T191|OAP|188644003|SNOMEDCT_US|Leukaemic reticuloendotheliosis of unspecified sites|9940/3
C0023443|T191|OAP|85228003|SNOMEDCT_US|Leukemic reticuloendotheliosis|9940/3
C0023443|T191|SY|54087003|SNOMEDCT_US|Leukemic reticuloendotheliosis|9940/3
C0023443|T191|OF|85228003|SNOMEDCT_US|Leukemic reticuloendotheliosis -RETIRED-|9940/3
C0023443|T191|IS|85228003|SNOMEDCT_US|Leukemic reticuloendotheliosis -RETIRED-|9940/3
C0023443|T191|OAP|188653005|SNOMEDCT_US|Leukemic reticuloendotheliosis NOS|9940/3
C0023443|T191|OAP|188644003|SNOMEDCT_US|Leukemic reticuloendotheliosis of unspecified sites|9940/3
C0023443|T191|SYGB|118613001|SNOMEDCT_US|LRE - Leukaemic reticuloendotheliosis|9940/3
C0023443|T191|SY|118613001|SNOMEDCT_US|LRE - Leukemic reticuloendotheliosis|9940/3
C0023443|T191|PT|1771|WHO|HAIRY CELL LEUKAEMIA|9940/3
C0023480|T191|SY|0000007347|CHV|chronic myelomonocytic leukaemia|9945/3
C0023480|T191|SY|0000007347|CHV|chronic myelomonocytic leukemia|9945/3
C0023480|T191|PT|0000007347|CHV|cmml|9945/3
C0023480|T191|PT|HP:0012325|HPO|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|AB|C93.1|ICD10CM|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|HT|C93.1|ICD10CM|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|ET|C93.10|ICD10CM|Chronic myelomonocytic leukemia NOS|9945/3
C0023480|T191|PT|MTHU044790|ICPC2ICD10ENG|leukemia; myelomonocytic, chronic|9945/3
C0023480|T191|PT|MTHU050874|ICPC2ICD10ENG|myelomonocytic; leukemia, chronic|9945/3
C0023480|T191|PT|10009018|MDR|Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|LLT|10009018|MDR|Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|LLT|10054350|MDR|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|MTH_PT|10009018|MDR|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|PT|35942|MEDCIN|chronic myelomonocytic leukemia|9945/3
C0023480|T191|SY|35942|MEDCIN|CMML|9945/3
C0023480|T191|PM|D015477|MSH|Chronic Myelomonocytic Leukemia|9945/3
C0023480|T191|PM|D015477|MSH|Chronic Myelomonocytic Leukemias|9945/3
C0023480|T191|PM|D015477|MSH|Leukemia, Chronic Myelomonocytic|9945/3
C0023480|T191|MH|D015477|MSH|Leukemia, Myelomonocytic, Chronic|9945/3
C0023480|T191|PM|D015477|MSH|Leukemias, Chronic Myelomonocytic|9945/3
C0023480|T191|ET|D015477|MSH|Myelomonocytic Leukemia, Chronic|9945/3
C0023480|T191|PM|D015477|MSH|Myelomonocytic Leukemias, Chronic|9945/3
C0023480|T191|PN|NOCODE|MTH|Leukemia, Myelomonocytic, Chronic|9945/3
C0023480|T191|PT|C3178|NCI|Chronic Myelomonocytic Leukemia|9945/3
C0023480|T191|SY|TCGA|NCI|Chronic Myelomonocytic Leukemia|9945/3
C0023480|T191|AB|C3178|NCI|CMML|9945/3
C0023480|T191|PT|C3178|NCI_CPTAC|Chronic Myelomonocytic Leukemia|9945/3
C0023480|T191|PT|10009018|NCI_CTEP-SDC|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|SY|C3178|NCI_CTRP|Chronic Myelomonocytic Leukemia|9945/3
C0023480|T191|PT|CDR0000367436|NCI_NCI-GLOSS|chronic myelomonocytic leukemia|9945/3
C0023480|T191|PT|CDR0000367437|NCI_NCI-GLOSS|CMML|9945/3
C0023480|T191|PT|CDR0000040361|PDQ|chronic myelomonocytic leukemia|9945/3
C0023480|T191|AB|CDR0000040361|PDQ|CMML|9945/3
C0023480|T191|SY|CDR0000040361|PDQ|myelomonocytic leukemia, chronic|9945/3
C0023480|T191|AB|B691.|RCD|Chronic myelomonocyt leukaemia|9945/3
C0023480|T191|PT|B691.|RCD|Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|AB|B691.|RCD|CMML - Chron myelomonocyt leuk|9945/3
C0023480|T191|SY|B691.|RCD|CMML - Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|AB|B691.|RCDAE|Chronic myelomonocyt leukemia|9945/3
C0023480|T191|PT|B691.|RCDAE|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|SY|B691.|RCDAE|CMML - Chronic myelomonocytic leukemia|9945/3
C0023480|T191|OP|BBr68|RCDSA|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|OA|BBr68|RCDSY|Chrn myelomonocytic leukaem|9945/3
C0023480|T191|OP|BBr68|RCDSY|Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|OAP|188769006|SNOMEDCT_US|Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|OAP|79660002|SNOMEDCT_US|Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|PTGB|128831004|SNOMEDCT_US|Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|PTGB|127225006|SNOMEDCT_US|Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|IS|79660002|SNOMEDCT_US|Chronic myelomonocytic leukaemia -RETIRED-|9945/3
C0023480|T191|PT|127225006|SNOMEDCT_US|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|OAP|79660002|SNOMEDCT_US|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|OAP|188769006|SNOMEDCT_US|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|PT|128831004|SNOMEDCT_US|Chronic myelomonocytic leukemia|9945/3
C0023480|T191|OF|79660002|SNOMEDCT_US|Chronic myelomonocytic leukemia -RETIRED-|9945/3
C0023480|T191|IS|79660002|SNOMEDCT_US|Chronic myelomonocytic leukemia -RETIRED-|9945/3
C0023480|T191|OAS|188769006|SNOMEDCT_US|CMML - Chronic myelomonocytic leukaemia|9945/3
C0023480|T191|OAS|188769006|SNOMEDCT_US|CMML - Chronic myelomonocytic leukemia|9945/3
C0349639|T191|SY|0000031274|CHV|jmml|9946/3
C0349639|T191|SY|0000031274|CHV|juvenile myelomonocytic leukemia|9946/3
C0349639|T191|PT|HP:0012209|HPO|Juvenile myelomonocytic leukemia|9946/3
C0349639|T191|HT|C93.3|ICD10CM|Juvenile myelomonocytic leukemia|9946/3
C0349639|T191|AB|C93.3|ICD10CM|Juvenile myelomonocytic leukemia|9946/3
C0349639|T191|ET|C93.30|ICD10CM|Juvenile myelomonocytic leukemia NOS|9946/3
C0349639|T191|LLT|10023248|MDR|Juvenile chronic myeloid leukaemia|9946/3
C0349639|T191|LLT|10060498|MDR|Juvenile chronic myeloid leukemia|9946/3
C0349639|T191|LLT|10023249|MDR|Juvenile chronic myelomonocytic leukaemia|9946/3
C0349639|T191|PT|10023249|MDR|Juvenile chronic myelomonocytic leukaemia|9946/3
C0349639|T191|LLT|10054439|MDR|Juvenile chronic myelomonocytic leukemia|9946/3
C0349639|T191|MTH_PT|10023249|MDR|Juvenile chronic myelomonocytic leukemia|9946/3
C0349639|T191|PT|350014|MEDCIN|Juvenile chronic myeloid leukemia|9946/3
C0349639|T191|PT|230929|MEDCIN|juvenile myelomonocytic leukemia|9946/3
C0349639|T191|SY|230929|MEDCIN|leukemia juvenile myelomonocytic|9946/3
C0349639|T191|ET|D054429|MSH|Juvenile Chronic Myelogenous Leukemia|9946/3
C0349639|T191|ET|D054429|MSH|Juvenile Myelomonocytic Leukemia|9946/3
C0349639|T191|PM|D054429|MSH|Juvenile Myelomonocytic Leukemias|9946/3
C0349639|T191|ET|D054429|MSH|Leukemia, Juvenile Myelomonocytic|9946/3
C0349639|T191|MH|D054429|MSH|Leukemia, Myelomonocytic, Juvenile|9946/3
C0349639|T191|PM|D054429|MSH|Myelomonocytic Leukemia, Juvenile|9946/3
C0349639|T191|PM|D054429|MSH|Myelomonocytic Leukemias, Juvenile|9946/3
C0349639|T191|PN|NOCODE|MTH|Juvenile Myelomonocytic Leukemia|9946/3
C0349639|T191|AB|C9233|NCI|JCML|9946/3
C0349639|T191|AB|C9233|NCI|JMML|9946/3
C0349639|T191|OP|C9233|NCI|Juvenile Chronic Myelogenous Leukemia|9946/3
C0349639|T191|OP|C9233|NCI|Juvenile Chronic Myeloid Leukemia|9946/3
C0349639|T191|PT|C9233|NCI|Juvenile Myelomonocytic Leukemia|9946/3
C0349639|T191|SY|TCGA|NCI|Juvenile Myelomonocytic Leukemia|9946/3
C0349639|T191|PT|C9233|NCI_CPTAC|Juvenile Myelomonocytic Leukemia|9946/3
C0349639|T191|PT|10023249|NCI_CTEP-SDC|Juvenile myelomonocytic leukemia|9946/3
C0349639|T191|DN|C9233|NCI_CTRP|Juvenile Myelomonocytic Leukemia|9946/3
C0349639|T191|PT|CDR0000450126|NCI_NCI-GLOSS|JMML|9946/3
C0349639|T191|PT|CDR0000045048|NCI_NCI-GLOSS|juvenile myelomonocytic leukemia|9946/3
C0349639|T191|SY|C9233|NCI_NICHD|Chronic Myelomonocytic Leukemia|9946/3
C0349639|T191|SY|C9233|NCI_NICHD|JMML|9946/3
C0349639|T191|PT|C9233|NCI_NICHD|Juvenile Myelomonocytic Leukemia|9946/3
C0349639|T191|AB|CDR0000038439|PDQ|JCML|9946/3
C0349639|T191|SY|CDR0000038439|PDQ|JMML|9946/3
C0349639|T191|AB|CDR0000038439|PDQ|JMML|9946/3
C0349639|T191|IS|CDR0000038439|PDQ|juvenile chronic myelogenous leukemia|9946/3
C0349639|T191|SY|CDR0000038439|PDQ|juvenile chronic myelogenous leukemia|9946/3
C0349639|T191|SY|CDR0000038439|PDQ|juvenile chronic myeloid leukemia|9946/3
C0349639|T191|IS|CDR0000038439|PDQ|juvenile chronic myeloid leukemia|9946/3
C0349639|T191|PT|CDR0000038439|PDQ|juvenile myelomonocytic leukemia|9946/3
C0349639|T191|SY|CDR0000038439|PDQ|myelomonocytic leukemia, juvenile|9946/3
C0349639|T191|AB|Xa0SV|RCD|JCML - Juv chron myel leukaem|9946/3
C0349639|T191|SY|Xa0SV|RCD|JCML - Juvenile chronic myeloid leukaemia|9946/3
C0349639|T191|AB|Xa0SV|RCD|Juv chronic myeloid leukaemia|9946/3
C0349639|T191|PT|Xa0SV|RCD|Juvenile chronic myeloid leukaemia|9946/3
C0349639|T191|SY|Xa0SV|RCDAE|JCML - Juvenile chronic myeloid leukemia|9946/3
C0349639|T191|AB|Xa0SV|RCDAE|Juv chronic myeloid leukemia|9946/3
C0349639|T191|PT|Xa0SV|RCDAE|Juvenile chronic myeloid leukemia|9946/3
C0349639|T191|SYGB|277587001|SNOMEDCT_US|JCML - Juvenile chronic myeloid leukaemia|9946/3
C0349639|T191|SY|277587001|SNOMEDCT_US|JCML - Juvenile chronic myeloid leukemia|9946/3
C0349639|T191|PTGB|277587001|SNOMEDCT_US|Juvenile chronic myeloid leukaemia|9946/3
C0349639|T191|PT|277587001|SNOMEDCT_US|Juvenile chronic myeloid leukemia|9946/3
C0349639|T191|SYGB|128832006|SNOMEDCT_US|Juvenile chronic myelomonocytic leukaemia|9946/3
C0349639|T191|SY|128832006|SNOMEDCT_US|Juvenile chronic myelomonocytic leukemia|9946/3
C0349639|T191|PTGB|445227008|SNOMEDCT_US|Juvenile myelomonocytic leukaemia|9946/3
C0349639|T191|PTGB|128832006|SNOMEDCT_US|Juvenile myelomonocytic leukaemia|9946/3
C0349639|T191|PT|445227008|SNOMEDCT_US|Juvenile myelomonocytic leukemia|9946/3
C0349639|T191|PT|128832006|SNOMEDCT_US|Juvenile myelomonocytic leukemia|9946/3
C1292777|T191|ET|C94.8|ICD10CM|Aggressive NK-cell leukemia|9948/3
C1292777|T191|LLT|10028811|MDR|Natural killer-cell leukaemia|9948/3
C1292777|T191|PT|10028811|MDR|Natural killer-cell leukaemia|9948/3
C1292777|T191|LLT|10054481|MDR|Natural killer-cell leukemia|9948/3
C1292777|T191|MTH_PT|10028811|MDR|Natural killer-cell leukemia|9948/3
C1292777|T191|LLT|10029429|MDR|NK-cell leukaemia|9948/3
C1292777|T191|LLT|10029430|MDR|NK-cell leukemia|9948/3
C1292777|T191|PT|366679|MEDCIN|Aggressive natural killer-cell leukemia|9948/3
C1292777|T191|PT|230930|MEDCIN|aggressive NK-cell leukemia|9948/3
C1292777|T191|SY|230930|MEDCIN|leukemia aggressive NK-cell|9948/3
C1292777|T191|PN|NOCODE|MTH|Aggressive natural killer-cell leukemia|9948/3
C1292777|T191|PT|C8647|NCI|Aggressive NK-Cell Leukemia|9948/3
C1292777|T191|SY|TCGA|NCI|Aggressive NK-Cell Leukemia|9948/3
C1292777|T191|SY|C8647|NCI|Aggressive NK-Cell Leukemia/Lymphoma|9948/3
C1292777|T191|SY|C8647|NCI|Natural Killer Cell Leukemia|9948/3
C1292777|T191|SY|C8647|NCI|NK Cell Leukemia|9948/3
C1292777|T191|SY|C8647|NCI|NK-Cell Leukemia|9948/3
C1292777|T191|DN|C8647|NCI_CTRP|Aggressive NK-Cell Leukemia|9948/3
C1292777|T191|PT|CDR0000671058|PDQ|aggressive NK-cell leukemia|9948/3
C1292777|T191|PTGB|721310007|SNOMEDCT_US|Aggressive natural killer-cell leukaemia|9948/3
C1292777|T191|SYGB|128833001|SNOMEDCT_US|Aggressive natural killer-cell leukaemia|9948/3
C1292777|T191|PT|721310007|SNOMEDCT_US|Aggressive natural killer-cell leukemia|9948/3
C1292777|T191|SY|128833001|SNOMEDCT_US|Aggressive natural killer-cell leukemia|9948/3
C1292777|T191|SYGB|128833001|SNOMEDCT_US|Aggressive NK cell leukaemia|9948/3
C1292777|T191|SY|128833001|SNOMEDCT_US|Aggressive NK cell leukemia|9948/3
C1292777|T191|PTGB|128833001|SNOMEDCT_US|Aggressive NK-cell leukaemia|9948/3
C1292777|T191|PT|128833001|SNOMEDCT_US|Aggressive NK-cell leukemia|9948/3
C0032463|T191|NP|0000023087|AOD|polycythemia vera|9950/3
C0032463|T191|AB|BI00325|BI|p vera|9950/3
C0032463|T191|PT|BI00325|BI|polycythemia vera|9950/3
C0032463|T191|PT|0042418|CCPSS|POLYCYTHEMIA VERA|9950/3
C0032463|T191|SY|0000009911|CHV|erythraemia|9950/3
C0032463|T191|SY|0000009911|CHV|erythremia|9950/3
C0032463|T191|SY|0000009911|CHV|erythrocythemia|9950/3
C0032463|T191|SY|0000009911|CHV|osler's disease|9950/3
C0032463|T191|SY|0000009911|CHV|p vera|9950/3
C0032463|T191|SY|0000009911|CHV|polycythaemia rubra vera|9950/3
C0032463|T191|SY|0000009911|CHV|polycythaemia vera|9950/3
C0032463|T191|SY|0000009911|CHV|polycythemia ruba vera|9950/3
C0032463|T191|SY|0000009911|CHV|polycythemia rubra vera|9950/3
C0032463|T191|PT|0000009911|CHV|polycythemia vera|9950/3
C0032463|T191|SY|0000009911|CHV|primary polycythemia|9950/3
C0032463|T191|SY|0000009911|CHV|proliferative polycythemia|9950/3
C0032463|T191|SY|0000009911|CHV|splenomegalic polycythemia|9950/3
C0032463|T191|SY|0000009911|CHV|vaquez's disease|9950/3
C0032463|T191|PT|NOCODE|COSTAR|Polycythemia Vera|9950/3
C0032463|T191|PT|2004-0979|CSP|polycythemia vera|9950/3
C0032463|T191|SY|NOCODE|DXP|ERYTHREMIA|9950/3
C0032463|T191|SY|NOCODE|DXP|OSLER-VAQUEZ DISEASE|9950/3
C0032463|T191|SY|NOCODE|DXP|POLYCYTHEMIA VERA|9950/3
C0032463|T191|DI|U001549|DXP|POLYCYTHEMIA, PRIMARY|9950/3
C0032463|T191|SY|NOCODE|DXP|POLYCYTHEMIA, SPLENOMEGALIC|9950/3
C0032463|T191|SY|NOCODE|DXP|VAQUEZ-OSLER DISEASE|9950/3
C0032463|T191|PT|D45|ICD10|Polycythaemia vera|9950/3
C0032463|T191|PT|D45|ICD10AE|Polycythemia vera|9950/3
C0032463|T191|PT|D45|ICD10CM|Polycythemia vera|9950/3
C0032463|T191|AB|D45|ICD10CM|Polycythemia vera|9950/3
C0032463|T191|PT|238.4|ICD9CM|Polycythemia vera|9950/3
C0032463|T191|AB|238.4|ICD9CM|Polycythemia vera|9950/3
C0032463|T191|PT|MTHU027038|ICPC2ICD10ENG|erythremia|9950/3
C0032463|T191|PT|MTHU056041|ICPC2ICD10ENG|Osler-Vaquez|9950/3
C0032463|T191|PT|MTHU060919|ICPC2ICD10ENG|polycythemia; rubra vera|9950/3
C0032463|T191|PT|MTHU060922|ICPC2ICD10ENG|polycythemia; vera|9950/3
C0032463|T191|PT|MTHU065159|ICPC2ICD10ENG|rubra; polycythemia rubra vera|9950/3
C0032463|T191|PT|MTHU079103|ICPC2ICD10ENG|Vaquez-Osler|9950/3
C0032463|T191|PT|MTHU079591|ICPC2ICD10ENG|vera; polycythemia|9950/3
C0032463|T191|PTN|B75004|ICPC2P|polycythaemia rubra vera|9950/3
C0032463|T191|PT|B75004|ICPC2P|Polycythaemia rubra vera|9950/3
C0032463|T191|MTH_PT|B75004|ICPC2P|Polycythemia rubra vera|9950/3
C0032463|T191|MTH_PTN|B75004|ICPC2P|polycythemia rubra vera|9950/3
C0032463|T191|PT|U003754|LCH|Polycythemia vera|9950/3
C0032463|T191|PT|sh85104611|LCH_NW|Polycythemia vera|9950/3
C0032463|T191|LLT|10036056|MDR|Polycythaemia rubra vera|9950/3
C0032463|T191|PT|10036057|MDR|Polycythaemia vera|9950/3
C0032463|T191|LLT|10036057|MDR|Polycythaemia vera|9950/3
C0032463|T191|LLT|10036060|MDR|Polycythemia rubra vera|9950/3
C0032463|T191|LLT|10036061|MDR|Polycythemia vera|9950/3
C0032463|T191|MTH_PT|10036057|MDR|Polycythemia vera|9950/3
C0032463|T191|LLT|10036725|MDR|Primary polycythaemia|9950/3
C0032463|T191|LLT|10036726|MDR|Primary polycythemia|9950/3
C0032463|T191|LLT|10064071|MDR|Vaquez's disease|9950/3
C0032463|T191|PT|30372|MEDCIN|polycythemia vera|9950/3
C0032463|T191|PM|D011087|MSH|Disease, Osler-Vaquez|9950/3
C0032463|T191|ET|D011087|MSH|Erythremia|9950/3
C0032463|T191|PM|D011087|MSH|Erythremias|9950/3
C0032463|T191|DEV|D011087|MSH|OSLER VAQUEZ DIS|9950/3
C0032463|T191|PM|D011087|MSH|Osler Vaquez Disease|9950/3
C0032463|T191|ET|D011087|MSH|Osler-Vaquez Disease|9950/3
C0032463|T191|ET|D011087|MSH|Polycythemia Ruba Vera|9950/3
C0032463|T191|PM|D011087|MSH|Polycythemia Ruba Veras|9950/3
C0032463|T191|ET|D011087|MSH|Polycythemia Rubra Vera|9950/3
C0032463|T191|PM|D011087|MSH|Polycythemia Rubra Veras|9950/3
C0032463|T191|MH|D011087|MSH|Polycythemia Vera|9950/3
C0032463|T191|PM|D011087|MSH|Polycythemia, Primary|9950/3
C0032463|T191|PM|D011087|MSH|Polycythemias, Primary|9950/3
C0032463|T191|ET|D011087|MSH|Primary Polycythemia|9950/3
C0032463|T191|PM|D011087|MSH|Primary Polycythemias|9950/3
C0032463|T191|PM|D011087|MSH|Ruba Vera, Polycythemia|9950/3
C0032463|T191|PM|D011087|MSH|Ruba Veras, Polycythemia|9950/3
C0032463|T191|PM|D011087|MSH|Vera, Polycythemia Ruba|9950/3
C0032463|T191|PM|D011087|MSH|Vera, Polycythemia Rubra|9950/3
C0032463|T191|PM|D011087|MSH|Veras, Polycythemia Ruba|9950/3
C0032463|T191|PM|D011087|MSH|Veras, Polycythemia Rubra|9950/3
C0032463|T191|PN|NOCODE|MTH|Polycythemia Vera|9950/3
C0032463|T191|SY|C3336|NCI|Polycythemia Rubra Vera|9950/3
C0032463|T191|PT|C3336|NCI|Polycythemia Vera|9950/3
C0032463|T191|SY|TCGA|NCI|Polycythemia Vera|9950/3
C0032463|T191|PT|C3336|NCI_CPTAC|Polycythemia Vera|9950/3
C0032463|T191|PT|10036061|NCI_CTEP-SDC|Polycythemia vera|9950/3
C0032463|T191|DN|C3336|NCI_CTRP|Polycythemia Vera|9950/3
C0032463|T191|PT|CDR0000426418|NCI_NCI-GLOSS|polycythemia vera|9950/3
C0032463|T191|PT|C3336|NCI_NICHD|Polycythemia Vera|9950/3
C0032463|T191|SY|CDR0000039350|PDQ|p.vera|9950/3
C0032463|T191|SY|CDR0000039350|PDQ|polycythaemia vera|9950/3
C0032463|T191|SY|CDR0000039350|PDQ|polycythemia ruba vera|9950/3
C0032463|T191|SY|CDR0000039350|PDQ|polycythemia rubra vera|9950/3
C0032463|T191|PT|CDR0000039350|PDQ|polycythemia vera|9950/3
C0032463|T191|SY|CDR0000039350|PDQ|PV|9950/3
C0032463|T191|PT|R0121727|QMR|POLYCYTHEMIA VERA|9950/3
C0032463|T191|PT|Xa0eC|RCD|Erythraemia|9950/3
C0032463|T191|PT|B934.|RCD|Polycythaemia rubra vera|9950/3
C0032463|T191|SY|B934.|RCD|Polycythaemia vera|9950/3
C0032463|T191|SY|B934.|RCD|PPP - Primary proliferative polycythaemia|9950/3
C0032463|T191|AB|B934.|RCD|PPP-Primary prolif polycythaem|9950/3
C0032463|T191|AB|B934.|RCD|Prim proliferat polycythaemia|9950/3
C0032463|T191|SY|B934.|RCD|Primary proliferative polycythaemia|9950/3
C0032463|T191|SY|B934.|RCD|PRV - Polycythaemia rubra vera|9950/3
C0032463|T191|PT|Xa0eC|RCDAE|Erythremia|9950/3
C0032463|T191|PT|B934.|RCDAE|Polycythemia rubra vera|9950/3
C0032463|T191|SY|B934.|RCDAE|Polycythemia vera|9950/3
C0032463|T191|SY|B934.|RCDAE|PPP - Primary proliferative polycythemia|9950/3
C0032463|T191|AB|B934.|RCDAE|Prim proliferat polycythemia|9950/3
C0032463|T191|SY|B934.|RCDAE|Primary proliferative polycythemia|9950/3
C0032463|T191|SY|B934.|RCDAE|PRV - Polycythemia rubra vera|9950/3
C0032463|T191|IS|BBs0.|RCDSA|Polycythemia rubra vera|9950/3
C0032463|T191|OP|BBs0.|RCDSA|Polycythemia vera|9950/3
C0032463|T191|IS|BBs0.|RCDSY|Polycythaemia rubra vera|9950/3
C0032463|T191|OP|BBs0.|RCDSY|Polycythaemia vera|9950/3
C0032463|T191|OAP|278190000|SNOMEDCT_US|Erythraemia|9950/3
C0032463|T191|OAP|278190000|SNOMEDCT_US|Erythremia|9950/3
C0032463|T191|SY|109992005|SNOMEDCT_US|Osler-Vaquez syndrome|9950/3
C0032463|T191|SY|109992005|SNOMEDCT_US|Osler's disease|9950/3
C0032463|T191|SYGB|128841001|SNOMEDCT_US|Polycythaemia rubra vera|9950/3
C0032463|T191|SYGB|109992005|SNOMEDCT_US|Polycythaemia rubra vera|9950/3
C0032463|T191|OAS|154644004|SNOMEDCT_US|Polycythaemia rubra vera|9950/3
C0032463|T191|OAS|269652000|SNOMEDCT_US|Polycythaemia rubra vera|9950/3
C0032463|T191|PTGB|128841001|SNOMEDCT_US|Polycythaemia vera|9950/3
C0032463|T191|OAP|31569001|SNOMEDCT_US|Polycythaemia vera|9950/3
C0032463|T191|OAS|154644004|SNOMEDCT_US|Polycythaemia vera|9950/3
C0032463|T191|OAS|269652000|SNOMEDCT_US|Polycythaemia vera|9950/3
C0032463|T191|SYGB|109992005|SNOMEDCT_US|Polycythaemia vera|9950/3
C0032463|T191|IS|31569001|SNOMEDCT_US|Polycythaemia vera -RETIRED-|9950/3
C0032463|T191|IS|31569001|SNOMEDCT_US|Polycythemia rubra vera|9950/3
C0032463|T191|SY|109992005|SNOMEDCT_US|Polycythemia rubra vera|9950/3
C0032463|T191|OAS|269652000|SNOMEDCT_US|Polycythemia rubra vera|9950/3
C0032463|T191|OAS|154644004|SNOMEDCT_US|Polycythemia rubra vera|9950/3
C0032463|T191|SY|128841001|SNOMEDCT_US|Polycythemia rubra vera|9950/3
C0032463|T191|OAP|31569001|SNOMEDCT_US|Polycythemia vera|9950/3
C0032463|T191|OAS|154644004|SNOMEDCT_US|Polycythemia vera|9950/3
C0032463|T191|PT|128841001|SNOMEDCT_US|Polycythemia vera|9950/3
C0032463|T191|OAS|269652000|SNOMEDCT_US|Polycythemia vera|9950/3
C0032463|T191|SY|109992005|SNOMEDCT_US|Polycythemia vera|9950/3
C0032463|T191|IS|31569001|SNOMEDCT_US|Polycythemia vera -RETIRED-|9950/3
C0032463|T191|OF|31569001|SNOMEDCT_US|Polycythemia vera -RETIRED-|9950/3
C0032463|T191|SYGB|109992005|SNOMEDCT_US|PPP - Primary proliferative polycythaemia|9950/3
C0032463|T191|SY|109992005|SNOMEDCT_US|PPP - Primary proliferative polycythemia|9950/3
C0032463|T191|SYGB|109992005|SNOMEDCT_US|Primary polycythaemia|9950/3
C0032463|T191|SYGB|109992005|SNOMEDCT_US|Primary proliferative polycythaemia|9950/3
C0032463|T191|SY|109992005|SNOMEDCT_US|Primary proliferative polycythemia|9950/3
C0032463|T191|SYGB|128841001|SNOMEDCT_US|Proliferative polycythaemia|9950/3
C0032463|T191|SY|128841001|SNOMEDCT_US|Proliferative polycythemia|9950/3
C0032463|T191|SYGB|109992005|SNOMEDCT_US|PRV - Polycythaemia rubra vera|9950/3
C0032463|T191|SY|109992005|SNOMEDCT_US|PRV - Polycythemia rubra vera|9950/3
C0032463|T191|SY|109992005|SNOMEDCT_US|Vaquez's disease|9950/3
C1292778|T191|PT|D47.1|ICD10|Chronic myeloproliferative disease|9960/3
C1292778|T191|AB|D47.1|ICD10CM|Chronic myeloproliferative disease|9960/3
C1292778|T191|PT|D47.1|ICD10CM|Chronic myeloproliferative disease|9960/3
C1292778|T191|PT|338489|MEDCIN|chronic myeloproliferative syndrome|9960/3
C1292778|T191|SY|338489|MEDCIN|myeloproliferative syndrome chronic|9960/3
C1292778|T191|PN|NOCODE|MTH|Chronic myeloproliferative disorder|9960/3
C1292778|T191|ET|238.7|MTHICD9|Chronic myeloproliferative disease NOS|9960/3
C1292778|T191|SY|C4345|NCI|Chronic Myeloproliferative Disease|9960/3
C1292778|T191|SY|C4345|NCI|Chronic Myeloproliferative Disorder|9960/3
C1292778|T191|SY|C4345|NCI|Chronic Myeloproliferative Neoplasm|9960/3
C1292778|T191|AB|C4345|NCI|CMPD|9960/3
C1292778|T191|SY|MPN-SAF|NCI|MPD|9960/3
C1292778|T191|AB|C4345|NCI|MPN|9960/3
C1292778|T191|SY|C4345|NCI|Myeloproliferative Disease|9960/3
C1292778|T191|SY|C4345|NCI|Myeloproliferative Disorder|9960/3
C1292778|T191|PT|C4345|NCI|Myeloproliferative Neoplasm|9960/3
C1292778|T191|SY|C4345|NCI|Myeloproliferative Tumor|9960/3
C1292778|T191|PT|C4345|NCI_CPTAC|Myeloproliferative Neoplasm|9960/3
C1292778|T191|DN|C4345|NCI_CTRP|Chronic Myeloproliferative Disease|9960/3
C1292778|T191|PT|CDR0000045210|NCI_NCI-GLOSS|myeloproliferative disorder|9960/3
C1292778|T191|SY|CDR0000039347|PDQ|chronic myeloproliferative disease|9960/3
C1292778|T191|SY|CDR0000039347|PDQ|chronic myeloproliferative disorders|9960/3
C1292778|T191|PT|CDR0000039347|PDQ|chronic myeloproliferative neoplasms|9960/3
C1292778|T191|AB|CDR0000039347|PDQ|CMPD|9960/3
C1292778|T191|OA|BBs2.|RCD|Chron myeloproliferative dis|9960/3
C1292778|T191|OP|BBs2.|RCD|Chronic myeloproliferative disease|9960/3
C1292778|T191|SY|128842008|SNOMEDCT_US|Chronic myeloproliferative disease|9960/3
C1292778|T191|IS|20921005|SNOMEDCT_US|Chronic myeloproliferative disease -RETIRED-|9960/3
C1292778|T191|OF|20921005|SNOMEDCT_US|Chronic myeloproliferative disease -RETIRED-|9960/3
C1292778|T191|SY|128842008|SNOMEDCT_US|Chronic myeloproliferative disease, no ICD-O subtype|9960/3
C1292778|T191|SY|128842008|SNOMEDCT_US|Chronic myeloproliferative disease, no International Classification of Diseases for Oncology subtype|9960/3
C1292778|T191|SY|115248004|SNOMEDCT_US|Chronic myeloproliferative disorder|9960/3
C1292778|T191|SY|128842008|SNOMEDCT_US|Chronic myeloproliferative disorder|9960/3
C1292778|T191|PT|115248004|SNOMEDCT_US|Myeloproliferative neoplasm|9960/3
C1292778|T191|PT|128842008|SNOMEDCT_US|Myeloproliferative neoplasm, no ICD-O subtype|9960/3
C0001815|T191|PT|1008871|CCPSS|MYELOID METAPLASIA AGNOGENIC|9961/3
C0001815|T191|PT|0000000825|CHV|agnogenic myeloid metaplasia|9961/3
C0001815|T191|SY|0000000825|CHV|aleukemic myelosis|9961/3
C0001815|T191|PT|0000042711|CHV|idiopathic myelofibrosis|9961/3
C0001815|T191|SY|0000021389|CHV|metaplasia myelofibrosis myeloid|9961/3
C0001815|T191|SY|0000042711|CHV|myelofibrosis idiopathic|9961/3
C0001815|T191|SY|0000042712|CHV|myelofibrosis primary|9961/3
C0001815|T191|PT|0000021389|CHV|myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|PT|0000042712|CHV|primary myelofibrosis|9961/3
C0001815|T191|GT|MARROW HYPERPLASIA|CST|MYELOSIS NONLEUKEMIC|9961/3
C0001815|T191|FI|U000410|DXP|BONE MARROW FIBROSIS|9961/3
C0001815|T191|SY|NOCODE|DXP|MOS|9961/3
C0001815|T191|SY|NOCODE|DXP|MYELOFIBROSIS|9961/3
C0001815|T191|SY|NOCODE|DXP|MYELOFIBROSIS AND MYELOID METAPLASIA|9961/3
C0001815|T191|SY|NOCODE|DXP|MYELOID METAPLASIA, AGNOGENIC|9961/3
C0001815|T191|SY|NOCODE|DXP|MYELOSCLEROSIS|9961/3
C0001815|T191|SY|NOCODE|DXP|MYELOSIS, ALEUKEMIC|9961/3
C0001815|T191|ET|D47.4|ICD10CM|Chronic idiopathic myelofibrosis|9961/3
C0001815|T191|AB|238.76|ICD9CM|Myelofi w myelo metaplas|9961/3
C0001815|T191|PT|238.76|ICD9CM|Myelofibrosis with myeloid metaplasia|9961/3
C0001815|T191|PT|MTHU004928|ICPC2ICD10ENG|aleukemic; myelosis|9961/3
C0001815|T191|PT|MTHU050861|ICPC2ICD10ENG|myeloid metaplasia; myelosclerosis|9961/3
C0001815|T191|PT|MTHU050916|ICPC2ICD10ENG|myelosclerosis; with myeloid metaplasia|9961/3
C0001815|T191|PT|MTHU050918|ICPC2ICD10ENG|myelosis; aleukemic|9961/3
C0001815|T191|PT|MTHU050923|ICPC2ICD10ENG|myelosis; nonleukemic|9961/3
C0001815|T191|PT|MTHU053301|ICPC2ICD10ENG|nonleukemic; myelosis|9961/3
C0001815|T191|LLT|10077161|MDR|Primary myelofibrosis|9961/3
C0001815|T191|PT|10077161|MDR|Primary myelofibrosis|9961/3
C0001815|T191|PT|311875|MEDCIN|idiopathic myelofibrosis|9961/3
C0001815|T191|PT|30306|MEDCIN|myelofibrosis with myeloid metaplasia|9961/3
C0001815|T191|PT|98887|MEDCIN|myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|PT|311873|MEDCIN|primary myelofibrosis|9961/3
C0001815|T191|ET|D055728|MSH|Agnogenic Myeloid Metaplasia|9961/3
C0001815|T191|PM|D055728|MSH|Agnogenic Myeloid Metaplasias|9961/3
C0001815|T191|PM|D055728|MSH|Bone Marrow Fibroses|9961/3
C0001815|T191|ET|D055728|MSH|Bone Marrow Fibrosis|9961/3
C0001815|T191|ET|D055728|MSH|Chronic Idiopathic Myelofibrosis|9961/3
C0001815|T191|PM|D055728|MSH|Fibroses, Bone Marrow|9961/3
C0001815|T191|ET|D055728|MSH|Fibrosis, Bone Marrow|9961/3
C0001815|T191|ET|D055728|MSH|Idiopathic Myelofibrosis|9961/3
C0001815|T191|PM|D055728|MSH|Metaplasia, Agnogenic Myeloid|9961/3
C0001815|T191|PM|D055728|MSH|Metaplasia, Myeloid|9961/3
C0001815|T191|PM|D055728|MSH|Metaplasias, Agnogenic Myeloid|9961/3
C0001815|T191|PM|D055728|MSH|Metaplasias, Myeloid|9961/3
C0001815|T191|PM|D055728|MSH|Myelofibroses|9961/3
C0001815|T191|PM|D055728|MSH|Myelofibroses, Primary|9961/3
C0001815|T191|ET|D055728|MSH|Myelofibrosis|9961/3
C0001815|T191|ET|D055728|MSH|Myelofibrosis With Myeloid Metaplasia|9961/3
C0001815|T191|PM|D055728|MSH|Myelofibrosis, Primary|9961/3
C0001815|T191|ET|D055728|MSH|Myeloid Metaplasia|9961/3
C0001815|T191|PM|D055728|MSH|Myeloid Metaplasia, Agnogenic|9961/3
C0001815|T191|PM|D055728|MSH|Myeloid Metaplasias|9961/3
C0001815|T191|PM|D055728|MSH|Myeloid Metaplasias, Agnogenic|9961/3
C0001815|T191|PM|D055728|MSH|Myeloscleroses|9961/3
C0001815|T191|ET|D055728|MSH|Myelosclerosis|9961/3
C0001815|T191|PM|D055728|MSH|Myeloses, Nonleukemic|9961/3
C0001815|T191|ET|D055728|MSH|Myelosis, Nonleukemic|9961/3
C0001815|T191|PM|D055728|MSH|Nonleukemic Myeloses|9961/3
C0001815|T191|PM|D055728|MSH|Nonleukemic Myelosis|9961/3
C0001815|T191|PM|D055728|MSH|Primary Myelofibroses|9961/3
C0001815|T191|MH|D055728|MSH|Primary Myelofibrosis|9961/3
C0001815|T191|SY|NOCODE|MTH|MYELOSIS NON-LEUKEMIC|9961/3
C0001815|T191|PN|NOCODE|MTH|Primary Myelofibrosis|9961/3
C0001815|T191|ET|238.76|MTHICD9|Agnogenic myeloid metaplasia|9961/3
C0001815|T191|ET|205.8|MTHICD9|Aleukemic myelosis|9961/3
C0001815|T191|ET|238.76|MTHICD9|Myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|ET|238.76|MTHICD9|Primary myelofibrosis|9961/3
C0001815|T191|SY|C2862|NCI|Agnogenic Myeloid Metaplasia|9961/3
C0001815|T191|AB|C2862|NCI|AMM|9961/3
C0001815|T191|SY|C2862|NCI|Chronic Idiopathic Myelofibrosis|9961/3
C0001815|T191|AB|C2862|NCI|CIMF|9961/3
C0001815|T191|SY|C2862|NCI|Idiopathic Bone Marrow Fibrosis|9961/3
C0001815|T191|SY|C2862|NCI|Idiopathic Myelofibrosis|9961/3
C0001815|T191|SY|C2862|NCI|Myelosclerosis with Myeloid Metaplasia|9961/3
C0001815|T191|SY|TCGA|NCI|Primary Myelofibrosis|9961/3
C0001815|T191|PT|C2862|NCI|Primary Myelofibrosis|9961/3
C0001815|T191|PT|C2862|NCI_CPTAC|Primary Myelofibrosis|9961/3
C0001815|T191|PT|10028537|NCI_CTEP-SDC|Chronic idiopathic myelofibrosis|9961/3
C0001815|T191|DN|C2862|NCI_CTRP|Primary Myelofibrosis|9961/3
C0001815|T191|PT|CDR0000306486|NCI_NCI-GLOSS|agnogenic myeloid metaplasia|9961/3
C0001815|T191|PT|CDR0000306487|NCI_NCI-GLOSS|chronic idiopathic myelofibrosis|9961/3
C0001815|T191|PT|CDR0000306490|NCI_NCI-GLOSS|idiopathic myelofibrosis|9961/3
C0001815|T191|PT|CDR0000306489|NCI_NCI-GLOSS|myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|SY|CDR0000039357|PDQ|agnogenic myeloid metaplasia|9961/3
C0001815|T191|AB|CDR0000039357|PDQ|AMM|9961/3
C0001815|T191|LV|CDR0000039357|PDQ|chronic idiopathic myelofibrosis|9961/3
C0001815|T191|SY|CDR0000039357|PDQ|chronic idiopathic myelofibrosis|9961/3
C0001815|T191|SY|CDR0000039357|PDQ|idiopathic bone marrow fibrosis|9961/3
C0001815|T191|SY|CDR0000039357|PDQ|idiopathic myelofibrosis|9961/3
C0001815|T191|OP|CDR0000042965|PDQ|idiopathic myelofibrosis|9961/3
C0001815|T191|SY|CDR0000039357|PDQ|myelofibrosis with myeloid metaplasia|9961/3
C0001815|T191|SY|CDR0000039357|PDQ|myeloid metaplasia, agnogenic|9961/3
C0001815|T191|SY|CDR0000039357|PDQ|myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|PT|CDR0000039357|PDQ|primary myelofibrosis|9961/3
C0001815|T191|OP|CDR0000042966|PDQ|primary myelofibrosis|9961/3
C0001815|T191|PT|R0121457|QMR|MYELOID METAPLASIA <PRIMARY MYELOFIBROSIS>|9961/3
C0001815|T191|SY|XaBBt|RCD|Megakaryocytic myelosclerosis|9961/3
C0001815|T191|AB|XaBBt|RCD|Myeloscleros + myeloid metapl|9961/3
C0001815|T191|PT|XaBBt|RCD|Myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|AB|BBs3.|RCDSY|Myeloscleros.+myeloid metap|9961/3
C0001815|T191|PT|BBs3.|RCDSY|Myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|SY|52967002|SNOMEDCT_US|Agnogenic myeloid metaplasia|9961/3
C0001815|T191|SY|128843003|SNOMEDCT_US|Agnogenic myeloid metaplasia|9961/3
C0001815|T191|SY|128843003|SNOMEDCT_US|Chronic idiopathic myelofibrosis|9961/3
C0001815|T191|SY|128843003|SNOMEDCT_US|Myelofibrosis as a result of myeloproliferative disease|9961/3
C0001815|T191|SY|307651005|SNOMEDCT_US|Myelofibrosis with myeloid metaplasia|9961/3
C0001815|T191|SY|128843003|SNOMEDCT_US|Myelofibrosis with myeloid metaplasia|9961/3
C0001815|T191|IS|22265001|SNOMEDCT_US|Myelofibrosis with myeloid metaplasia|9961/3
C0001815|T191|OAP|22265001|SNOMEDCT_US|Myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|OF|188773009|SNOMEDCT_US|Myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|PT|307651005|SNOMEDCT_US|Myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|PT|128843003|SNOMEDCT_US|Myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|OAP|188773009|SNOMEDCT_US|Myelosclerosis with myeloid metaplasia|9961/3
C0001815|T191|IS|22265001|SNOMEDCT_US|Myelosclerosis with myeloid metaplasia -RETIRED-|9961/3
C0001815|T191|OF|22265001|SNOMEDCT_US|Myelosclerosis with myeloid metaplasia -RETIRED-|9961/3
C0001815|T191|SY|128843003|SNOMEDCT_US|Primary myelofibrosis|9961/3
C0001815|T191|SY|307651005|SNOMEDCT_US|Primary myelofibrosis|9961/3
C0001815|T191|IT|0562|WHO|MYELOSIS NON-LEUKAEMIC|9961/3
C0040028|T047|SY|BI00328|BI|essential thrombocytosis|9962/3
C0040028|T047|PT|0057573|CCPSS|THROMBOCYTOSIS ESSENTIAL|9962/3
C0040028|T047|SY|0000012220|CHV|essential thrombocythaemia|9962/3
C0040028|T047|PT|0000012220|CHV|essential thrombocythemia|9962/3
C0040028|T047|PT|0000031201|CHV|essential thrombocytosis|9962/3
C0040028|T047|SY|0000012220|CHV|idiopathic thrombocythemia|9962/3
C0040028|T047|SY|0000012220|CHV|primary thrombocythemia|9962/3
C0040028|T047|SY|0000012220|CHV|thrombocythemia essential|9962/3
C0040028|T047|SY|0000031201|CHV|thrombocytosis essential|9962/3
C0040028|T047|PT|U000257|COSTAR|ESSENTIAL THROMBOCYTHEMIA|9962/3
C0040028|T047|ET|0446-2826|CSP|essential thrombocythemia|9962/3
C0040028|T047|PT|0446-2826|CSP|hemorrhagic thrombocythemia|9962/3
C0040028|T047|ET|0446-2826|CSP|idiopathic thrombocythemia|9962/3
C0040028|T047|ET|0446-2826|CSP|primary thrombocythemia|9962/3
C0040028|T047|SY|NOCODE|DXP|THROMBOCYTHEMIA, ESSENTIAL, WITH HEMORRHAGIC DIATHESIS|9962/3
C0040028|T047|DI|U001846|DXP|THROMBOCYTHEMIA, HEMORRHAGIC|9962/3
C0040028|T047|SY|NOCODE|DXP|THROMBOCYTHEMIA, IDIOPATHIC|9962/3
C0040028|T047|SY|NOCODE|DXP|THROMBOCYTHEMIA, PRIMARY HEMORRHAGIC|9962/3
C0040028|T047|PT|D75.2|ICD10|Essential thrombocytosis|9962/3
C0040028|T047|ET|D47.3|ICD10CM|Essential thrombocytosis|9962/3
C0040028|T047|ET|D47.3|ICD10CM|Idiopathic hemorrhagic thrombocythemia|9962/3
C0040028|T047|PT|238.71|ICD9CM|Essential thrombocythemia|9962/3
C0040028|T047|AB|238.71|ICD9CM|Essntial thrombocythemia|9962/3
C0040028|T047|PT|MTHU075538|ICPC2ICD10ENG|thrombocytosis; essential|9962/3
C0040028|T047|PTN|B83015|ICPC2P|essential thrombocytosis|9962/3
C0040028|T047|PT|B83015|ICPC2P|Thrombocytosis;essential|9962/3
C0040028|T047|LLT|10015493|MDR|Essential thrombocythaemia|9962/3
C0040028|T047|PT|10015493|MDR|Essential thrombocythaemia|9962/3
C0040028|T047|LLT|10015494|MDR|Essential thrombocythemia|9962/3
C0040028|T047|MTH_PT|10015493|MDR|Essential thrombocythemia|9962/3
C0040028|T047|LLT|10015495|MDR|Essential thrombocytosis|9962/3
C0040028|T047|OL|10021217|MDR|Ideopathic thrombocytosis|9962/3
C0040028|T047|LLT|10053263|MDR|Idiopathic thrombocytosis|9962/3
C0040028|T047|PT|311866|MEDCIN|essential hemorrhagic thrombocythemia|9962/3
C0040028|T047|PT|91365|MEDCIN|essential thrombocythemia|9962/3
C0040028|T047|PT|30300|MEDCIN|essential thrombocytosis|9962/3
C0040028|T047|PT|98886|MEDCIN|idiopathic thrombocythemia|9962/3
C0040028|T047|PT|311867|MEDCIN|primary thrombocytosis|9962/3
C0040028|T047|PM|D013920|MSH|Essential Thrombocythemia|9962/3
C0040028|T047|PM|D013920|MSH|Essential Thrombocythemias|9962/3
C0040028|T047|ET|D013920|MSH|Hemorrhagic Thrombocythemia|9962/3
C0040028|T047|PM|D013920|MSH|Hemorrhagic Thrombocythemias|9962/3
C0040028|T047|PM|D013920|MSH|Idiopathic Thrombocythemia|9962/3
C0040028|T047|PM|D013920|MSH|Idiopathic Thrombocythemias|9962/3
C0040028|T047|ET|D013920|MSH|Primary Thrombocythemia|9962/3
C0040028|T047|PM|D013920|MSH|Primary Thrombocythemias|9962/3
C0040028|T047|PM|D013920|MSH|Primary Thrombocytoses|9962/3
C0040028|T047|PM|D013920|MSH|Primary Thrombocytosis|9962/3
C0040028|T047|MH|D013920|MSH|Thrombocythemia, Essential|9962/3
C0040028|T047|ET|D013920|MSH|Thrombocythemia, Hemorrhagic|9962/3
C0040028|T047|ET|D013920|MSH|Thrombocythemia, Idiopathic|9962/3
C0040028|T047|ET|D013920|MSH|Thrombocythemia, Primary|9962/3
C0040028|T047|PM|D013920|MSH|Thrombocythemias, Essential|9962/3
C0040028|T047|PM|D013920|MSH|Thrombocythemias, Hemorrhagic|9962/3
C0040028|T047|PM|D013920|MSH|Thrombocythemias, Idiopathic|9962/3
C0040028|T047|PM|D013920|MSH|Thrombocythemias, Primary|9962/3
C0040028|T047|PM|D013920|MSH|Thrombocytoses, Primary|9962/3
C0040028|T047|ET|D013920|MSH|Thrombocytosis, Primary|9962/3
C0040028|T047|PN|NOCODE|MTH|Thrombocythemia, Essential|9962/3
C0040028|T047|ET|238.71|MTHICD9|Essential hemorrhagic thrombocythemia|9962/3
C0040028|T047|ET|238.71|MTHICD9|Essential thrombocytosis|9962/3
C0040028|T047|ET|238.71|MTHICD9|Primary thrombocytosis|9962/3
C0040028|T047|SY|C3407|NCI|Essential Thrombocytemia|9962/3
C0040028|T047|PT|C3407|NCI|Essential Thrombocythemia|9962/3
C0040028|T047|SY|TCGA|NCI|Essential Thrombocythemia|9962/3
C0040028|T047|SY|C3407|NCI|Essential Thrombocytosis|9962/3
C0040028|T047|SY|C3407|NCI|Idiopathic Thrombocythemia|9962/3
C0040028|T047|SY|C3407|NCI|Primary Thrombocythemia|9962/3
C0040028|T047|SY|C3407|NCI|Primary Thrombocytosis|9962/3
C0040028|T047|PT|C3407|NCI_CPTAC|Essential Thrombocythemia|9962/3
C0040028|T047|PT|10015493|NCI_CTEP-SDC|Essential thrombocythemia|9962/3
C0040028|T047|DN|C3407|NCI_CTRP|Essential Thrombocythemia|9962/3
C0040028|T047|PT|CDR0000256562|NCI_NCI-GLOSS|essential thrombocythemia|9962/3
C0040028|T047|PT|CDR0000256561|NCI_NCI-GLOSS|essential thrombocytosis|9962/3
C0040028|T047|PT|C3407|NCI_NICHD|Essential Thrombocythemia|9962/3
C0040028|T047|SY|C3407|NCI_NICHD|Essential Thrombocytosis|9962/3
C0040028|T047|SY|C3407|NCI_NICHD|ET|9962/3
C0040028|T047|PT|CDR0000039361|PDQ|essential thrombocythemia|9962/3
C0040028|T047|SY|CDR0000039361|PDQ|hemorrhagic thrombocythemia|9962/3
C0040028|T047|SY|CDR0000039361|PDQ|idiopathic thrombocytosis|9962/3
C0040028|T047|SY|CDR0000039361|PDQ|primary thrombocytosis|9962/3
C0040028|T047|SY|CDR0000039361|PDQ|thrombocythemia, essential|9962/3
C0040028|T047|PT|R0121884|QMR|THROMBOCYTHEMIA IDIOPATHIC|9962/3
C0040028|T047|PT|X20FX|RCD|Essential thrombocythaemia|9962/3
C0040028|T047|OP|D3y0.|RCD|Essential thrombocytosis|9962/3
C0040028|T047|AB|X20FX|RCD|ET - Essent thrombocythaemia|9962/3
C0040028|T047|SY|X20FX|RCD|ET - Essential thrombocythaemia|9962/3
C0040028|T047|PT|XaBBu|RCD|Idiopathic thrombocythaemia|9962/3
C0040028|T047|PT|X20FX|RCDAE|Essential thrombocythemia|9962/3
C0040028|T047|AB|X20FX|RCDAE|ET - Essent thrombocythemia|9962/3
C0040028|T047|SY|X20FX|RCDAE|ET - Essential thrombocythemia|9962/3
C0040028|T047|PT|XaBBu|RCDAE|Idiopathic thrombocythemia|9962/3
C0040028|T047|PT|BBs4.|RCDSA|Idiopathic thrombocythemia|9962/3
C0040028|T047|PT|BBs4.|RCDSY|Idiopathic thrombocythaemia|9962/3
C0040028|T047|SYGB|128844009|SNOMEDCT_US|Essential haemorrhagic thrombocythaemia|9962/3
C0040028|T047|IS|65471002|SNOMEDCT_US|Essential hemorrhagic thrombocythemia|9962/3
C0040028|T047|SY|128844009|SNOMEDCT_US|Essential hemorrhagic thrombocythemia|9962/3
C0040028|T047|PTGB|128844009|SNOMEDCT_US|Essential thrombocythaemia|9962/3
C0040028|T047|PTGB|109994006|SNOMEDCT_US|Essential thrombocythaemia|9962/3
C0040028|T047|OAP|189513005|SNOMEDCT_US|Essential thrombocythaemia|9962/3
C0040028|T047|OAP|234499005|SNOMEDCT_US|Essential thrombocythaemia|9962/3
C0040028|T047|OF|189513005|SNOMEDCT_US|Essential thrombocythaemia|9962/3
C0040028|T047|OF|234499005|SNOMEDCT_US|Essential thrombocythaemia|9962/3
C0040028|T047|IS|65471002|SNOMEDCT_US|Essential thrombocythemia|9962/3
C0040028|T047|PT|109994006|SNOMEDCT_US|Essential thrombocythemia|9962/3
C0040028|T047|PT|128844009|SNOMEDCT_US|Essential thrombocythemia|9962/3
C0040028|T047|OAP|234499005|SNOMEDCT_US|Essential thrombocythemia|9962/3
C0040028|T047|OAP|189513005|SNOMEDCT_US|Essential thrombocythemia|9962/3
C0040028|T047|SY|109994006|SNOMEDCT_US|Essential thrombocytosis|9962/3
C0040028|T047|OAP|191333009|SNOMEDCT_US|Essential thrombocytosis|9962/3
C0040028|T047|OAS|234499005|SNOMEDCT_US|ET - Essential thrombocythaemia|9962/3
C0040028|T047|OAS|234499005|SNOMEDCT_US|ET - Essential thrombocythemia|9962/3
C0040028|T047|SYGB|128844009|SNOMEDCT_US|Idiopathic haemorrhagic thrombocythaemia|9962/3
C0040028|T047|IS|65471002|SNOMEDCT_US|Idiopathic hemorrhagic thrombocythemia|9962/3
C0040028|T047|SY|128844009|SNOMEDCT_US|Idiopathic hemorrhagic thrombocythemia|9962/3
C0040028|T047|OAP|65471002|SNOMEDCT_US|Idiopathic thrombocythaemia|9962/3
C0040028|T047|OAS|189508006|SNOMEDCT_US|Idiopathic thrombocythaemia|9962/3
C0040028|T047|OF|189514004|SNOMEDCT_US|Idiopathic thrombocythaemia|9962/3
C0040028|T047|SYGB|109994006|SNOMEDCT_US|Idiopathic thrombocythaemia|9962/3
C0040028|T047|OAP|307652003|SNOMEDCT_US|Idiopathic thrombocythaemia|9962/3
C0040028|T047|SYGB|128844009|SNOMEDCT_US|Idiopathic thrombocythaemia|9962/3
C0040028|T047|OAP|189514004|SNOMEDCT_US|Idiopathic thrombocythaemia|9962/3
C0040028|T047|IS|65471002|SNOMEDCT_US|Idiopathic thrombocythaemia -RETIRED-|9962/3
C0040028|T047|OAP|307652003|SNOMEDCT_US|Idiopathic thrombocythemia|9962/3
C0040028|T047|SY|109994006|SNOMEDCT_US|Idiopathic thrombocythemia|9962/3
C0040028|T047|OAP|189514004|SNOMEDCT_US|Idiopathic thrombocythemia|9962/3
C0040028|T047|SY|128844009|SNOMEDCT_US|Idiopathic thrombocythemia|9962/3
C0040028|T047|OAP|65471002|SNOMEDCT_US|Idiopathic thrombocythemia|9962/3
C0040028|T047|OAS|189508006|SNOMEDCT_US|Idiopathic thrombocythemia|9962/3
C0040028|T047|IS|65471002|SNOMEDCT_US|Idiopathic thrombocythemia -RETIRED-|9962/3
C0040028|T047|OF|65471002|SNOMEDCT_US|Idiopathic thrombocythemia -RETIRED-|9962/3
C0040028|T047|SYGB|128844009|SNOMEDCT_US|Primary thrombocythaemia|9962/3
C0040028|T047|SY|128844009|SNOMEDCT_US|Primary thrombocythemia|9962/3
C0023481|T191|ET|D47.1|ICD10CM|Chronic neutrophilic leukemia|9963/3
C0023481|T191|PT|230931|MEDCIN|chronic neutrophilic leukemia|9963/3
C0023481|T191|SY|230931|MEDCIN|leukemia chronic neutrophilic|9963/3
C0023481|T191|PM|D015467|MSH|Chronic Neutrophilic Leukemia|9963/3
C0023481|T191|PM|D015467|MSH|Chronic Neutrophilic Leukemias|9963/3
C0023481|T191|PM|D015467|MSH|Leukemia, Chronic Neutrophilic|9963/3
C0023481|T191|MH|D015467|MSH|Leukemia, Neutrophilic, Chronic|9963/3
C0023481|T191|PM|D015467|MSH|Leukemias, Chronic Neutrophilic|9963/3
C0023481|T191|ET|D015467|MSH|Neutrophilic Leukemia, Chronic|9963/3
C0023481|T191|PM|D015467|MSH|Neutrophilic Leukemias, Chronic|9963/3
C0023481|T191|PN|NOCODE|MTH|Chronic Neutrophilic Leukemia|9963/3
C0023481|T191|PT|C3179|NCI|Chronic Neutrophilic Leukemia|9963/3
C0023481|T191|SY|TCGA|NCI|Chronic Neutrophilic Leukemia|9963/3
C0023481|T191|SY|C3179|NCI|Neutrophilic Leukemia|9963/3
C0023481|T191|DN|C3179|NCI_CTRP|Chronic Neutrophilic Leukemia|9963/3
C0023481|T191|PT|CDR0000426409|NCI_NCI-GLOSS|chronic neutrophilic leukemia|9963/3
C0023481|T191|PT|CDR0000276485|PDQ|chronic neutrophilic leukemia|9963/3
C0023481|T191|SY|CDR0000276485|PDQ|neutrophilic leukemia|9963/3
C0023481|T191|PT|B6512|RCD|Chronic neutrophilic leukaemia|9963/3
C0023481|T191|PT|B6512|RCDAE|Chronic neutrophilic leukemia|9963/3
C0023481|T191|PTGB|188734009|SNOMEDCT_US|Chronic neutrophilic leukaemia|9963/3
C0023481|T191|PTGB|128834007|SNOMEDCT_US|Chronic neutrophilic leukaemia|9963/3
C0023481|T191|PT|188734009|SNOMEDCT_US|Chronic neutrophilic leukemia|9963/3
C0023481|T191|PT|128834007|SNOMEDCT_US|Chronic neutrophilic leukemia|9963/3
C0346421|T191|SY|0000031070|CHV|chronic eosinophilic leukemia|9964/3
C1540912|T047|PT|0000031070|CHV|hypereosinophilic syndrome|9964/3
C0206141|T047|ET|0427-6368|CSP|idiopathic hypereosinophilic syndrome|9964/3
C1540912|T047|DI|U000872|DXP|HYPEREOSINOPHILIC SYNDROME|9964/3
C0346421|T191|LLT|10065854|MDR|Chronic eosinophilic leukaemia|9964/3
C0346421|T191|PT|10065854|MDR|Chronic eosinophilic leukaemia|9964/3
C0346421|T191|MTH_PT|10065854|MDR|Chronic eosinophilic leukemia|9964/3
C0346421|T191|LLT|10065872|MDR|Chronic eosinophilic leukemia|9964/3
C1540912|T047|PT|10048643|MDR|Hypereosinophilic syndrome|9964/3
C1540912|T047|LLT|10048643|MDR|Hypereosinophilic syndrome|9964/3
C0346421|T191|PT|331704|MEDCIN|chronic eosinophilic leukemia|9964/3
C0346421|T191|SY|331704|MEDCIN|chronic leukemia eosinophilic|9964/3
C1540912|T047|PT|30380|MEDCIN|hypereosinophilic syndrome|9964/3
C1540912|T047|ET|4589|MEDLINEPLUS|Hypereosinophilic Syndrome|9964/3
C0346421|T191|PCE|C580364|MSH|Chronic Eosinophilic Leukemia|9964/3
C1540912|T047|MH|D017681|MSH|Hypereosinophilic Syndrome|9964/3
C0206141|T047|ET|D017681|MSH|Hypereosinophilic Syndrome, Idiopathic|9964/3
C1540912|T047|PM|D017681|MSH|Hypereosinophilic Syndromes|9964/3
C0206141|T047|PM|D017681|MSH|Hypereosinophilic Syndromes, Idiopathic|9964/3
C0206141|T047|PEP|D017681|MSH|Idiopathic Hypereosinophilic Syndrome|9964/3
C0206141|T047|PM|D017681|MSH|Idiopathic Hypereosinophilic Syndromes|9964/3
C1540912|T047|PM|D017681|MSH|Syndrome, Hypereosinophilic|9964/3
C0206141|T047|PM|D017681|MSH|Syndrome, Idiopathic Hypereosinophilic|9964/3
C1540912|T047|PM|D017681|MSH|Syndromes, Hypereosinophilic|9964/3
C0206141|T047|PM|D017681|MSH|Syndromes, Idiopathic Hypereosinophilic|9964/3
C0346421|T191|PN|NOCODE|MTH|Chronic eosinophilic leukemia|9964/3
C1540912|T047|PN|NOCODE|MTH|Hypereosinophilic syndrome|9964/3
C0206141|T047|PN|NOCODE|MTH|Idiopathic Hypereosinophilic Syndrome|9964/3
C0346421|T191|AB|C4563|NCI|CEL|9964/3
C0346421|T191|SY|C4563|NCI|Chronic Eosinophilic Leukemia|9964/3
C0346421|T191|SY|C4563|NCI|Chronic Eosinophilic Leukemia, NOS|9964/3
C0346421|T191|PT|C4563|NCI|Chronic Eosinophilic Leukemia, Not Otherwise Specified|9964/3
C0346421|T191|SY|TCGA|NCI|Chronic Eosinophilic Leukemia, Not Otherwise Specified|9964/3
C0346421|T191|SY|C4563|NCI|Eosinophilic Leukemia|9964/3
C1540912|T047|PT|C27038|NCI|Hypereosinophilic Syndrome|9964/3
C1540912|T047|SY|TCGA|NCI|Hypereosinophilic Syndrome|9964/3
C0346421|T191|SY|10065872|NCI_CTEP-SDC|CEL/Hypereosinophilic syndrome|9964/3
C0346421|T191|PT|10065872|NCI_CTEP-SDC|Chronic eosinophilic leukemia/hypereosinophilic syndrome|9964/3
C0346421|T191|DN|C4563|NCI_CTRP|Chronic Eosinophilic Leukemia|9964/3
C1540912|T047|DN|C27038|NCI_CTRP|Hypereosinophilic Syndrome|9964/3
C0346421|T191|PT|CDR0000426408|NCI_NCI-GLOSS|chronic eosinophilic leukemia|9964/3
C0346421|T191|PT|CDR0000276487|PDQ|chronic eosinophilic leukemia|9964/3
C0346421|T191|PT|B6510|RCD|Chronic eosinophilic leukaemia|9964/3
C1540912|T047|PT|X20Dr|RCD|Hypereosinophilic syndrome|9964/3
C0346421|T191|PT|B6510|RCDAE|Chronic eosinophilic leukemia|9964/3
C0346421|T191|PTGB|413836008|SNOMEDCT_US|Chronic eosinophilic leukaemia|9964/3
C0346421|T191|PTGB|188733003|SNOMEDCT_US|Chronic eosinophilic leukaemia|9964/3
C0346421|T191|SYGB|128835008|SNOMEDCT_US|Chronic eosinophilic leukaemia|9964/3
C0346421|T191|SY|128835008|SNOMEDCT_US|Chronic eosinophilic leukemia|9964/3
C0346421|T191|PT|188733003|SNOMEDCT_US|Chronic eosinophilic leukemia|9964/3
C0346421|T191|PT|413836008|SNOMEDCT_US|Chronic eosinophilic leukemia|9964/3
C0206141|T047|IS|423294001|SNOMEDCT_US|HES|9964/3
C1540912|T047|SY|393573009|SNOMEDCT_US|HES - hypereosinophilic syndrome|9964/3
C1540912|T047|PT|128835008|SNOMEDCT_US|Hypereosinophilic syndrome|9964/3
C1540912|T047|PT|393573009|SNOMEDCT_US|Hypereosinophilic syndrome|9964/3
C1540912|T047|OAS|26328002|SNOMEDCT_US|Hypereosinophilic syndrome|9964/3
C1540912|T047|OF|393573009|SNOMEDCT_US|Hypereosinophilic syndrome|9964/3
C0206141|T047|IS|423294001|SNOMEDCT_US|Hypereosinophilic syndrome|9964/3
C1540912|T047|SY|128835008|SNOMEDCT_US|Hypereosinophilic syndrome/chronic eosinophilic leukemia|9964/3
C0206141|T047|PT|423294001|SNOMEDCT_US|Idiopathic hypereosinophilic syndrome|9964/3
C0206141|T047|PT|414450004|SNOMEDCT_US|Idiopathic hypereosinophilic syndrome|9964/3
C2827360|T191|SY|C84275|NCI|Myeloid and Lymphoid Neoplasms with PDGFRA Rearrangement|9965/3
C2827360|T191|PT|C84275|NCI|Myeloid/Lymphoid Neoplasms with PDGFRA Rearrangement|9965/3
C2827360|T191|SY|450940003|SNOMEDCT_US|Myeloid and lymphoid neoplasms with PDGFRA rearrangement|9965/3
C2827360|T191|PT|450940003|SNOMEDCT_US|Myeloid or lymphoid neoplasm with alpha-type platelet-derived growth factor receptor gene rearrangement|9965/3
C2827360|T191|SY|450940003|SNOMEDCT_US|Myeloid or lymphoid neoplasm with PDGFRA rearrangement|9965/3
C2827361|T191|SY|C84276|NCI|Myeloid and Lymphoid Neoplasms with PDGFRB Rearrangement|9966/3
C2827361|T191|SY|C84276|NCI|Myeloid Neoplasms with PDGFRB Rearrangement|9966/3
C2827361|T191|PT|C84276|NCI|Myeloid/Lymphoid Neoplasms with PDGFRB Rearrangement|9966/3
C3472621|T191|OP|450941004|SNOMEDCT_US|Myeloid neoplasm with beta-type platelet-derived growth factor gene rearrangement|9966/3
C3472621|T191|PT|450941004|SNOMEDCT_US|Myeloid neoplasm with beta-type platelet-derived growth factor receptor gene rearrangement|9966/3
C3472621|T191|SY|450941004|SNOMEDCT_US|Myeloid neoplasm with PDGFRB rearrangement|9966/3
C2827362|T191|SY|C84277|NCI|8p11 Myeloproliferative Syndrome|9967/3
C2827362|T191|SY|C84277|NCI|8p11 Stem Cell Leukemia/Lymphoma Syndrome|9967/3
C2827362|T191|SY|C84277|NCI|8p11 Stem Cell Lymphoma/Leukemia Syndrome|9967/3
C2827362|T191|SY|C84277|NCI|8p11 Stem Cell Syndrome|9967/3
C2827362|T191|SY|C84277|NCI|Myeloid and Lymphoid Neoplasms with FGFR1 Rearrangement|9967/3
C2827362|T191|PT|C84277|NCI|Myeloid/Lymphoid Neoplasms with FGFR1 Rearrangement|9967/3
C3472622|T191|SY|450942006|SNOMEDCT_US|Myeloid or lymphoid neoplasm with FGFR1 abnormality|9967/3
C3472622|T191|PT|450942006|SNOMEDCT_US|Myeloid or lymphoid neoplasm with fibroblast growth factor receptor 1 abnormality|9967/3
C0024314|T191|SY|0000007624|CHV|diseases lymphoproliferative|9970/1
C0024314|T191|SY|0000007624|CHV|disorders lymphoproliferative|9970/1
C0024314|T191|SY|0000007624|CHV|duncan syndrome|9970/1
C0024314|T191|SY|0000007624|CHV|duncan's syndrome|9970/1
C0024314|T191|SY|0000007624|CHV|duncans syndrome|9970/1
C0024314|T191|SY|0000007624|CHV|lymphoproliferative disease|9970/1
C0024314|T191|PT|0000007624|CHV|lymphoproliferative disorder|9970/1
C0024314|T191|SY|0000007624|CHV|lymphoproliferative disorder nos|9970/1
C0024314|T191|SY|0000007624|CHV|lymphoproliferative disorders|9970/1
C0024314|T191|PT|HP:0005523|HPO|Lymphoproliferative disorder|9970/1
C0024314|T191|ET|HP:0005523|HPO|Lymphoproliferative disorders|9970/1
C0024314|T191|ET|D47.9|ICD10CM|Lymphoproliferative disease NOS|9970/1
C0024314|T191|PT|MTHU046871|ICPC2ICD10ENG|lymphoproliferative; disorder|9970/1
C0024314|T191|PT|U002767|LCH|Lymphoproliferative disorders|9970/1
C0024314|T191|PT|sh85079155|LCH_NW|Lymphoproliferative disorders|9970/1
C0024314|T191|LLT|10068350|MDR|Duncan syndrome|9970/1
C0024314|T191|PT|10061232|MDR|Lymphoproliferative disorder|9970/1
C0024314|T191|LLT|10061232|MDR|Lymphoproliferative disorder|9970/1
C0024314|T191|LLT|10025351|MDR|Lymphoproliferative disorder NOS|9970/1
C0024314|T191|PT|312073|MEDCIN|lymphoproliferative disease|9970/1
C0024314|T191|PM|D008232|MSH|Disorder, Lymphoproliferative|9970/1
C0024314|T191|PM|D008232|MSH|Disorders, Lymphoproliferative|9970/1
C0024314|T191|DEV|D008232|MSH|LYMPHOPROLIFERATIVE DIS|9970/1
C0024314|T191|PM|D008232|MSH|Lymphoproliferative Disorder|9970/1
C0024314|T191|MH|D008232|MSH|Lymphoproliferative Disorders|9970/1
C0024314|T191|PN|NOCODE|MTH|Lymphoproliferative Disorders|9970/1
C0024314|T191|PT|C9308|NCI|Lymphoproliferative Disorder|9970/1
C0024314|T191|DN|C9308|NCI_CTRP|Lymphoproliferative Disorder|9970/1
C0024314|T191|PT|CDR0000045767|NCI_NCI-GLOSS|lymphoproliferative disorder|9970/1
C0024314|T191|PT|CDR0000617669|PDQ|lymphoproliferative disorder|9970/1
C0024314|T191|ET|CDR0000617669|PDQ|Lymphoproliferative disorder|9970/1
C0024314|T191|SY|X20Ik|RCD|Duncan's syndrome|9970/1
C0024314|T191|PT|Xa0QI|RCD|Lymphoproliferative disorder|9970/1
C0024314|T191|SY|77121009|SNOMEDCT_US|Duncan's syndrome|9970/1
C0024314|T191|PT|84631004|SNOMEDCT_US|Lymphoproliferative disease|9970/1
C0024314|T191|SY|84631004|SNOMEDCT_US|Lymphoproliferative disease, no ICD-O subtype|9970/1
C0024314|T191|SY|84631004|SNOMEDCT_US|Lymphoproliferative disease, no International Classification of Diseases for Oncology subtype|9970/1
C0024314|T191|IS|84631004|SNOMEDCT_US|Lymphoproliferative disease, NOS|9970/1
C0024314|T191|PT|414629003|SNOMEDCT_US|Lymphoproliferative disorder|9970/1
C0024314|T191|PT|277466009|SNOMEDCT_US|Lymphoproliferative disorder|9970/1
C0432487|T191|AB|238.77|ICD9CM|Post tp lymphprolif dis|9971/1
C0432487|T191|LLT|10051358|MDR|Post transplant lymphoproliferative disorder|9971/1
C0432487|T191|PT|10051358|MDR|Post transplant lymphoproliferative disorder|9971/1
C0432487|T191|PN|NOCODE|MTH|Post-transplant lymphoproliferative disorder|9971/1
C0432487|T191|ET|238.77|MTHICD9|Post-transplant lymphoproliferative disorder|9971/1
C0432487|T191|ET|238.77|MTHICD9|PTLD|9971/1
C0432487|T191|PT|C4727|NCI|Post-Transplant Lymphoproliferative Disorder|9971/1
C0432487|T191|AB|C4727|NCI|PTLD|9971/1
C0432487|T191|DN|C4727|NCI_CTRP|Post-Transplant Lymphoproliferative Disorder|9971/1
C0432487|T191|PT|CDR0000468786|NCI_NCI-GLOSS|post-transplant lymphoproliferative disorder|9971/1
C0432487|T191|PT|CDR0000512811|NCI_NCI-GLOSS|PTLD|9971/1
C0432487|T191|PT|C4727|NCI_NICHD|Post-transplant Lymphoproliferative Disorder|9971/1
C0432487|T191|PT|CDR0000038607|PDQ|post-transplant lymphoproliferative disorder|9971/1
C0432487|T191|AB|CDR0000038607|PDQ|PTLD|9971/1
C0432487|T191|AB|X78FF|RCD|Post-transp lymphoprolif dis|9971/1
C0432487|T191|PT|X78FF|RCD|Post-transplant lymphoproliferative disorder|9971/1
C0432487|T191|SY|X78FF|RCD|PTLD - Post-transplant lymphoproliferative disorder|9971/1
C0432487|T191|AB|X78FF|RCD|PTLD-Post-trns lymphprolif dis|9971/1
C5190713|T191|PT|782919005|SNOMEDCT_US|Classical Hodgkin lymphoma type posttransplant lymphoproliferative disorder|9971/1
C0432487|T191|PT|254290004|SNOMEDCT_US|Lymphoproliferative disorder following transplantation|9971/1
C0432487|T191|PT|450943001|SNOMEDCT_US|Post transplant lymphoproliferative disorder|9971/1
C0432487|T191|SY|450943001|SNOMEDCT_US|Post transplant lymphoproliferative disorder, no ICD-O subtype|9971/1
C0432487|T191|SY|450943001|SNOMEDCT_US|Post transplant lymphoproliferative disorder, no International Classification of Diseases for Oncology subtype|9971/1
C0432487|T191|SY|254290004|SNOMEDCT_US|Post-transplant lymphoproliferative disorder|9971/1
C0432487|T191|OAP|127219007|SNOMEDCT_US|Post-transplantation lymphoproliferative syndrome|9971/1
C0432487|T191|SY|254290004|SNOMEDCT_US|Post-transplantation lymphoproliferative syndrome|9971/1
C0432487|T191|SY|450943001|SNOMEDCT_US|PTLD|9971/1
C0432487|T191|SY|254290004|SNOMEDCT_US|PTLD - Post-transplant lymphoproliferative disorder|9971/1
C4518573|T191|PT|733081008|SNOMEDCT_US|Reactive plasmacytic hyperplasia|9971/1
C1301361|T191|SY|C7183|NCI|Polymorphic B-Cell Lymphoma|9971/3
C1301361|T191|PT|C7183|NCI|Polymorphic Post-Transplant Lymphoproliferative Disorder|9971/3
C1301361|T191|SY|TCGA|NCI|Polymorphic Post-Transplant Lymphoproliferative Disorder|9971/3
C1301361|T191|SY|C7183|NCI|Polymorphic PTLD|9971/3
C1301361|T191|PT|762316003|SNOMEDCT_US|Polymorphic lymphoproliferative disorder following transplant|9971/3
C1301361|T191|OAP|450944007|SNOMEDCT_US|Polymorphic post transplant lymphoproliferative disorder|9971/3
C1301361|T191|SY|762316003|SNOMEDCT_US|Polymorphic post-transplant lymphoproliferative disorder|9971/3
C1301361|T191|PT|397351004|SNOMEDCT_US|Post-transplant lymphoproliferative disorder, polymorphic|9971/3
C1292778|T191|PT|D47.1|ICD10|Chronic myeloproliferative disease|9975/1
C1292778|T191|AB|D47.1|ICD10CM|Chronic myeloproliferative disease|9975/1
C1292778|T191|PT|D47.1|ICD10CM|Chronic myeloproliferative disease|9975/1
C1292778|T191|PT|338489|MEDCIN|chronic myeloproliferative syndrome|9975/1
C1292778|T191|SY|338489|MEDCIN|myeloproliferative syndrome chronic|9975/1
C1292778|T191|PN|NOCODE|MTH|Chronic myeloproliferative disorder|9975/1
C1292778|T191|ET|238.7|MTHICD9|Chronic myeloproliferative disease NOS|9975/1
C1292778|T191|SY|C4345|NCI|Chronic Myeloproliferative Disease|9975/1
C1292778|T191|SY|C4345|NCI|Chronic Myeloproliferative Disorder|9975/1
C1292778|T191|SY|C4345|NCI|Chronic Myeloproliferative Neoplasm|9975/1
C1292778|T191|AB|C4345|NCI|CMPD|9975/1
C1292778|T191|SY|MPN-SAF|NCI|MPD|9975/1
C1292778|T191|AB|C4345|NCI|MPN|9975/1
C2939461|T191|SY|C9290|NCI|Myeloid Malignancy|9975/1
C2939461|T191|PT|C9290|NCI|Myeloid Neoplasm|9975/1
C2939461|T191|SY|C9290|NCI|Myeloid Tumor|9975/1
C1292778|T191|SY|C4345|NCI|Myeloproliferative Disease|9975/1
C1292778|T191|SY|C4345|NCI|Myeloproliferative Disorder|9975/1
C1292778|T191|PT|C4345|NCI|Myeloproliferative Neoplasm|9975/1
C1292778|T191|SY|C4345|NCI|Myeloproliferative Tumor|9975/1
C2939461|T191|PT|C9290|NCI_CPTAC|Myeloid Neoplasm|9975/1
C1292778|T191|PT|C4345|NCI_CPTAC|Myeloproliferative Neoplasm|9975/1
C1292778|T191|DN|C4345|NCI_CTRP|Chronic Myeloproliferative Disease|9975/1
C2939461|T191|DN|C9290|NCI_CTRP|Myeloid Neoplasm|9975/1
C2939461|T191|PT|C9290|NCI_CTRP|Myeloid Neoplasm|9975/1
C1292778|T191|PT|CDR0000045210|NCI_NCI-GLOSS|myeloproliferative disorder|9975/1
C1292778|T191|SY|CDR0000039347|PDQ|chronic myeloproliferative disease|9975/1
C1292778|T191|SY|CDR0000039347|PDQ|chronic myeloproliferative disorders|9975/1
C1292778|T191|PT|CDR0000039347|PDQ|chronic myeloproliferative neoplasms|9975/1
C1292778|T191|AB|CDR0000039347|PDQ|CMPD|9975/1
C1292778|T191|OA|BBs2.|RCD|Chron myeloproliferative dis|9975/1
C1292778|T191|OP|BBs2.|RCD|Chronic myeloproliferative disease|9975/1
C1292778|T191|SY|128842008|SNOMEDCT_US|Chronic myeloproliferative disease|9975/1
C1292778|T191|IS|20921005|SNOMEDCT_US|Chronic myeloproliferative disease -RETIRED-|9975/1
C1292778|T191|OF|20921005|SNOMEDCT_US|Chronic myeloproliferative disease -RETIRED-|9975/1
C1292778|T191|SY|128842008|SNOMEDCT_US|Chronic myeloproliferative disease, no ICD-O subtype|9975/1
C1292778|T191|SY|128842008|SNOMEDCT_US|Chronic myeloproliferative disease, no International Classification of Diseases for Oncology subtype|9975/1
C1292778|T191|SY|115248004|SNOMEDCT_US|Chronic myeloproliferative disorder|9975/1
C1292778|T191|SY|128842008|SNOMEDCT_US|Chronic myeloproliferative disorder|9975/1
C2939461|T191|PT|414792005|SNOMEDCT_US|Myeloid neoplasm|9975/1
C1292778|T191|PT|115248004|SNOMEDCT_US|Myeloproliferative neoplasm|9975/1
C1292778|T191|PT|128842008|SNOMEDCT_US|Myeloproliferative neoplasm, no ICD-O subtype|9975/1
C1301355|T191|LA|LA26797-3|LNC|Myelodysplastic/myeloproliferative neoplasm|9975/3
C1301355|T191|SY|355240|MEDCIN|bone marrow neoplasm myelodysplastic / myeloproliferative disease|9975/3
C1328061|T191|SY|355241|MEDCIN|bone marrow neoplasm myelodysplastic / myeloproliferative disease unclassifiable|9975/3
C1301355|T191|PT|355240|MEDCIN|myelodysplastic / myeloproliferative disease|9975/3
C1328061|T191|PT|355241|MEDCIN|myelodysplastic / myeloproliferative neoplasm, unclassifiable|9975/3
C1301355|T191|PM|D054437|MSH|Disease, Myelodysplastic-Myeloproliferative|9975/3
C1301355|T191|PM|D054437|MSH|Disease, Myeloproliferative-Myelodisplastic|9975/3
C1301355|T191|PM|D054437|MSH|Diseases, Myelodysplastic-Myeloproliferative|9975/3
C1301355|T191|PM|D054437|MSH|Diseases, Myeloproliferative-Myelodisplastic|9975/3
C1301355|T191|PM|D054437|MSH|Myelodysplastic Myeloproliferative Diseases|9975/3
C1301355|T191|PM|D054437|MSH|Myelodysplastic-Myeloproliferative Disease|9975/3
C1301355|T191|MH|D054437|MSH|Myelodysplastic-Myeloproliferative Diseases|9975/3
C1301355|T191|PM|D054437|MSH|Myeloproliferative Myelodisplastic Diseases|9975/3
C1301355|T191|PM|D054437|MSH|Myeloproliferative-Myelodisplastic Disease|9975/3
C1301355|T191|ET|D054437|MSH|Myeloproliferative-Myelodisplastic Diseases|9975/3
C1301355|T191|PN|NOCODE|MTH|Myelodysplastic-Myeloproliferative Diseases|9975/3
C1328061|T191|PN|NOCODE|MTH|Myelodysplastic/myeloproliferative neoplasm, unclassifiable|9975/3
C1333046|T191|PN|NOCODE|MTH|Myeloproliferative Neoplasm, Unclassifiable|9975/3
C1333046|T191|SY|C27350|NCI|Chronic Myeloproliferative Disease, Unclassifiable|9975/3
C1333046|T191|SY|C27350|NCI|Chronic Myeloproliferative Disorder, Unclassifiable|9975/3
C1333046|T191|AB|C27350|NCI|CMPD-U|9975/3
C1333046|T191|AB|C27350|NCI|CMPD, U|9975/3
C1301355|T191|AB|C27262|NCI|MDS-MPD|9975/3
C1301355|T191|AB|C27262|NCI|MDS/MPD|9975/3
C1328061|T191|AB|C27780|NCI|MDS/MPD-U|9975/3
C1328061|T191|AB|C27780|NCI|MDS/MPD, U|9975/3
C1301355|T191|AB|C27262|NCI|MDS/MPN|9975/3
C1328061|T191|AB|C27780|NCI|MDS/MPN-U|9975/3
C1328061|T191|AB|C27780|NCI|MDS/MPN, U|9975/3
C1328061|T191|SY|C27780|NCI|Mixed Myelodysplastic/Myeloproliferative Disease, Unclassifiable|9975/3
C1328061|T191|SY|C27780|NCI|Mixed Myeloproliferative/Myelodysplastic Syndrome, Unclassifiable|9975/3
C1301355|T191|AB|C27262|NCI|MPD-MDS|9975/3
C1301355|T191|AB|C27262|NCI|MPD/MDS|9975/3
C1333046|T191|AB|C27350|NCI|MPN-U|9975/3
C1333046|T191|AB|C27350|NCI|MPN, U|9975/3
C1301355|T191|SY|C27262|NCI|Myelodysplastic/Myeloproliferative Disease|9975/3
C1328061|T191|SY|C27780|NCI|Myelodysplastic/Myeloproliferative Disease, Unclassifiable|9975/3
C1301355|T191|SY|C27262|NCI|Myelodysplastic/Myeloproliferative Diseases|9975/3
C1301355|T191|SY|C27262|NCI|Myelodysplastic/Myeloproliferative Disorder|9975/3
C1301355|T191|SY|C27262|NCI|Myelodysplastic/Myeloproliferative Disorders|9975/3
C1301355|T191|PT|C27262|NCI|Myelodysplastic/Myeloproliferative Neoplasm|9975/3
C1328061|T191|PT|C27780|NCI|Myelodysplastic/Myeloproliferative Neoplasm, Unclassifiable|9975/3
C1328061|T191|SY|TCGA|NCI|Myelodysplastic/Myeloproliferative Neoplasm, Unclassifiable|9975/3
C1333046|T191|PT|C27350|NCI|Myeloproliferative Neoplasm, Unclassifiable|9975/3
C1301355|T191|SY|C27262|NCI|Myeloproliferative/Myelodysplastic Disorders|9975/3
C1301355|T191|SY|C27262|NCI|Myeloproliferative/Myelodysplastic Syndromes|9975/3
C1333046|T191|SY|C27350|NCI|Unclassifiable Chronic Myeloproliferative Disease|9975/3
C1333046|T191|SY|C27350|NCI|Unclassifiable Chronic Myeloproliferative Disorder|9975/3
C1328061|T191|SY|C27780|NCI|Unclassifiable Myelodysplastic/Myeloproliferative Disease|9975/3
C1328061|T191|SY|C27780|NCI|Unclassifiable Myeloproliferative/Myelodysplastic Syndrome|9975/3
C1301355|T191|PT|C27262|NCI_CPTAC|Myelodysplastic/Myeloproliferative Neoplasm|9975/3
C1301355|T191|DN|C27262|NCI_CTRP|Myelodysplastic/Myeloproliferative Disease|9975/3
C1328061|T191|DN|C27780|NCI_CTRP|Myelodysplastic/Myeloproliferative Neoplasm, Unclassifiable|9975/3
C1328061|T191|SY|CDR0000335177|PDQ|Mixed Myeloproliferative/Myelodysplastic Syndrome, Unclassifiable|9975/3
C1301355|T191|ET|CDR0000335173|PDQ|Myelodysplastic/myeloproliferative diseases|9975/3
C1328061|T191|PT|CDR0000335177|PDQ|myelodysplastic/myeloproliferative neoplasm, unclassifiable|9975/3
C1301355|T191|PT|CDR0000335173|PDQ|myelodysplastic/myeloproliferative neoplasms|9975/3
C1328061|T191|SY|CDR0000335177|PDQ|Unclassifiable Myeloproliferative/Myelodysplastic Syndrome|9975/3
C1301355|T191|PT|445738007|SNOMEDCT_US|Myelodysplastic/myeloproliferative disease|9975/3
C1301355|T191|PT|397336008|SNOMEDCT_US|Myelodysplastic/myeloproliferative disease|9975/3
C1328061|T191|PT|447596005|SNOMEDCT_US|Myelodysplastic/myeloproliferative neoplasm, unclassifiable|9975/3
C1328061|T191|SY|447240002|SNOMEDCT_US|Myelodysplastic/myeloproliferative neoplasm, unclassifiable|9975/3
C1328061|T191|PT|447240002|SNOMEDCT_US|Myeloproliferative neoplasm, unclassifiable|9975/3
C0002893|T047|PT|0042076|CCPSS|ANEMIA REFRACTORY|9980/3
C0002893|T047|SY|0000001133|CHV|anemia refractory|9980/3
C0002893|T047|SY|0000058157|CHV|refractory anaemia|9980/3
C0002893|T047|SY|0000001133|CHV|refractory anaemia|9980/3
C0002893|T047|PT|0000001133|CHV|refractory anemia|9980/3
C0002893|T047|PT|0000058157|CHV|refractory anemia|9980/3
C0002893|T047|SY|0000001133|CHV|refractory anemias|9980/3
C0002893|T047|GT|ANEMIA REFRACT|CST|ANEMIA REFRACTORY|9980/3
C0002893|T047|PT|ANEMIA REFRACT|CST|REFRACTORY ANEMIA|9980/3
C0002893|T047|SY|NOCODE|DXP|ANEMIA, REFRACTORY|9980/3
C0002893|T047|PT|HP:0005505|HPO|Refractory anemia|9980/3
C0002893|T047|PT|MTHU006001|ICPC2ICD10ENG|anemia; refractory|9980/3
C0002893|T047|PT|MTHU064005|ICPC2ICD10ENG|refractory; anemia|9980/3
C0002893|T047|LLT|10055722|MDR|Anaemia refractory|9980/3
C0002893|T047|LLT|10002311|MDR|Anemia refractory|9980/3
C0002893|T047|LLT|10038269|MDR|Refractory anaemia|9980/3
C0002893|T047|LLT|10038273|MDR|Refractory anemia|9980/3
C0002893|T047|SY|30368|MEDCIN|anemia refractory|9980/3
C0002893|T047|PT|30368|MEDCIN|refractory anemia|9980/3
C0002893|T047|MH|D000753|MSH|Anemia, Refractory|9980/3
C0002893|T047|PM|D000753|MSH|Anemias, Refractory|9980/3
C0002893|T047|ET|D000753|MSH|Refractory Anemia|9980/3
C0002893|T047|PM|D000753|MSH|Refractory Anemias|9980/3
C0002893|T047|PN|NOCODE|MTH|Refractory anemias|9980/3
C0002893|T047|SY|C2872|NCI|Aregenerative Anemia|9980/3
C0002893|T047|AB|C2872|NCI|RA|9980/3
C0002893|T047|PT|C2872|NCI|Refractory Anemia|9980/3
C0002893|T047|SY|TCGA|NCI|Refractory Anemia|9980/3
C0002893|T047|PT|C2872|NCI_CPTAC|Refractory Anemia|9980/3
C0002893|T047|DN|C2872|NCI_CTRP|Refractory Anemia|9980/3
C0002893|T047|PT|CDR0000040357|PDQ|refractory anemia|9980/3
C0002893|T047|SY|X20CK|RCD|Erythrodysplasia|9980/3
C0002893|T047|SY|X20CK|RCD|RA - Refractory anaemia|9980/3
C0002893|T047|PT|X20CK|RCD|Refractory anaemia|9980/3
C0002893|T047|SY|X20CK|RCDAE|RA - Refractory anemia|9980/3
C0002893|T047|PT|X20CK|RCDAE|Refractory anemia|9980/3
C0002893|T047|PTGB|128845005|SNOMEDCT_US|Refractory anaemia|9980/3
C0002893|T047|OAP|123306007|SNOMEDCT_US|Refractory anaemia|9980/3
C0002893|T047|OAP|191267001|SNOMEDCT_US|Refractory anaemia|9980/3
C0002893|T047|OAP|77704005|SNOMEDCT_US|Refractory anaemia|9980/3
C0002893|T047|OF|191267001|SNOMEDCT_US|Refractory anaemia|9980/3
C0002893|T047|IS|77704005|SNOMEDCT_US|Refractory anaemia -RETIRED-|9980/3
C0002893|T047|IS|123306007|SNOMEDCT_US|Refractory anaemia -RETIRED-|9980/3
C0002893|T047|OAP|77704005|SNOMEDCT_US|Refractory anemia|9980/3
C0002893|T047|PT|128845005|SNOMEDCT_US|Refractory anemia|9980/3
C0002893|T047|OAP|123306007|SNOMEDCT_US|Refractory anemia|9980/3
C0002893|T047|OAP|191267001|SNOMEDCT_US|Refractory anemia|9980/3
C0002893|T047|IS|123306007|SNOMEDCT_US|Refractory anemia -RETIRED-|9980/3
C0002893|T047|IS|77704005|SNOMEDCT_US|Refractory anemia -RETIRED-|9980/3
C0002893|T047|OF|77704005|SNOMEDCT_US|Refractory anemia -RETIRED-|9980/3
C0002893|T047|OF|123306007|SNOMEDCT_US|Refractory anemia -RETIRED-|9980/3
C0002893|T047|IS|77704005|SNOMEDCT_US|Refractory anemia, NOS|9980/3
C1264195|T191|SY|HP:0004828|HPO|Myelodysplasia with sideroblastosis|9982/3
C1264195|T191|PT|HP:0004828|HPO|Refractory anemia with ringed sideroblasts|9982/3
C0334679|T191|PT|D46.1|ICD10|Refractory anaemia with sideroblasts|9982/3
C0334679|T191|PT|D46.1|ICD10AE|Refractory anemia with sideroblasts|9982/3
C1264195|T191|ET|D46.1|ICD10CM|RARS|9982/3
C1264195|T191|AB|D46.1|ICD10CM|Refractory anemia with ring sideroblasts|9982/3
C1264195|T191|PT|D46.1|ICD10CM|Refractory anemia with ring sideroblasts|9982/3
C0334679|T191|PT|MTHU006005|ICPC2ICD10ENG|anemia; refractory, with sideroblasts|9982/3
C0334679|T191|PT|MTHU064009|ICPC2ICD10ENG|refractory; anemia, with sideroblasts|9982/3
C1264195|T191|LLT|10038272|MDR|Refractory anaemia with ringed sideroblasts|9982/3
C1264195|T191|PT|10038272|MDR|Refractory anaemia with ringed sideroblasts|9982/3
C1264195|T191|LLT|10054594|MDR|Refractory anemia with ringed sideroblasts|9982/3
C1264195|T191|MTH_PT|10038272|MDR|Refractory anemia with ringed sideroblasts|9982/3
C1264195|T191|PT|333430|MEDCIN|Refractory anemia with ring sideroblasts|9982/3
C2826330|T191|PT|366673|MEDCIN|Refractory anemia with ring sideroblasts associated with marked thrombocytosis|9982/3
C1264195|T191|PN|NOCODE|MTH|Refractory anemia with ringed sideroblasts|9982/3
C0334679|T191|PN|NOCODE|MTH|Refractory anemia with sideroblasts|9982/3
C2826330|T191|SY|C82616|NCI|Essential Thrombocythemia with Ring Sideroblasts|9982/3
C1264195|T191|AB|C4036|NCI|MDS-RS|9982/3
C2826330|T191|SY|C82616|NCI|MDS/MPN with Ring Sideroblasts and Thrombocytosis|9982/3
C2826330|T191|AB|C82616|NCI|MDS/MPN-RS-T|9982/3
C1264195|T191|PT|C4036|NCI|Myelodysplastic Syndrome with Ring Sideroblasts|9982/3
C2826330|T191|PT|C82616|NCI|Myelodysplastic/Myeloproliferative Neoplasm with Ring Sideroblasts and Thrombocytosis|9982/3
C1264195|T191|SY|C4036|NCI|Pure Sideroblastic Anemia|9982/3
C1264195|T191|AB|C4036|NCI|RARS|9982/3
C2826330|T191|AB|C82616|NCI|RARS-T|9982/3
C1264195|T191|SY|C4036|NCI|Refractory Anemia with Ring Sideroblasts|9982/3
C2826330|T191|SY|C82616|NCI|Refractory Anemia with Ring Sideroblasts Associated with Marked Thrombocytosis|9982/3
C1264195|T191|SY|TCGA|NCI|Refractory Anemia with Ringed Sideroblasts|9982/3
C1264195|T191|DN|C4036|NCI_CTRP|Myelodysplastic Syndrome with Ring Sideroblasts|9982/3
C1264195|T191|SY|CDR0000040358|PDQ|pure sideroblastic anemia|9982/3
C1264195|T191|AB|CDR0000040358|PDQ|RARS|9982/3
C1264195|T191|PT|CDR0000040358|PDQ|refractory anemia with ringed sideroblasts|9982/3
C1264195|T191|SY|Xa0Se|RCD|RARS - Refractory anaemia with ringed sideroblasts|9982/3
C1264195|T191|AB|Xa0Se|RCD|RARS-Ref anaem+ring sideroblst|9982/3
C1264195|T191|AB|Xa0Se|RCD|Ref anaem+ringed sideroblasts|9982/3
C0334679|T191|OA|B9371|RCD|Refr anaemia with sideroblasts|9982/3
C1264195|T191|PT|Xa0Se|RCD|Refractory anaemia with ringed sideroblasts|9982/3
C0334679|T191|OP|B9371|RCD|Refractory anaemia with sideroblasts|9982/3
C1264195|T191|SY|Xa0Se|RCDAE|RARS - Refractory anemia with ringed sideroblasts|9982/3
C0334679|T191|OA|B9371|RCDAE|Refr anemia with sideroblasts|9982/3
C1264195|T191|PT|Xa0Se|RCDAE|Refractory anemia with ringed sideroblasts|9982/3
C0334679|T191|OP|B9371|RCDAE|Refractory anemia with sideroblasts|9982/3
C0334679|T191|OA|BBmA.|RCDSA|Refract anemia+sideroblast|9982/3
C0334679|T191|OP|BBmA.|RCDSA|Refractory anemia with sideroblasts|9982/3
C0334679|T191|OA|BBmA.|RCDSY|Refract anaemia+sideroblast|9982/3
C0334679|T191|OP|BBmA.|RCDSY|Refractory anaemia with sideroblasts|9982/3
C1264195|T191|SY|128846006|SNOMEDCT_US|RARS|9982/3
C1264195|T191|OAS|277595002|SNOMEDCT_US|RARS - Refractory anaemia with ringed sideroblasts|9982/3
C1264195|T191|OAS|277595002|SNOMEDCT_US|RARS - Refractory anemia with ringed sideroblasts|9982/3
C2826330|T191|SY|703817002|SNOMEDCT_US|RARS-T|9982/3
C2826330|T191|PTGB|703817002|SNOMEDCT_US|Refractory anaemia with ring sideroblasts associated with marked thrombocytosis|9982/3
C1264195|T191|OAP|56837009|SNOMEDCT_US|Refractory anaemia with ringed sideroblasts|9982/3
C1264195|T191|OAP|277595002|SNOMEDCT_US|Refractory anaemia with ringed sideroblasts|9982/3
C1264195|T191|SYGB|109998009|SNOMEDCT_US|Refractory anaemia with ringed sideroblasts|9982/3
C1264195|T191|SYGB|128846006|SNOMEDCT_US|Refractory anaemia with ringed sideroblasts|9982/3
C1264195|T191|IS|56837009|SNOMEDCT_US|Refractory anaemia with ringed sideroblasts -RETIRED-|9982/3
C0334679|T191|SYGB|109998009|SNOMEDCT_US|Refractory anaemia with sideroblasts|9982/3
C0334679|T191|OAP|189510008|SNOMEDCT_US|Refractory anaemia with sideroblasts|9982/3
C0334679|T191|PTGB|128846006|SNOMEDCT_US|Refractory anaemia with sideroblasts|9982/3
C2826330|T191|PT|703817002|SNOMEDCT_US|Refractory anemia with ring sideroblasts associated with marked thrombocytosis|9982/3
C1264195|T191|OAP|277595002|SNOMEDCT_US|Refractory anemia with ringed sideroblasts|9982/3
C1264195|T191|SY|109998009|SNOMEDCT_US|Refractory anemia with ringed sideroblasts|9982/3
C1264195|T191|SY|128846006|SNOMEDCT_US|Refractory anemia with ringed sideroblasts|9982/3
C1264195|T191|IS|56837009|SNOMEDCT_US|Refractory anemia with ringed sideroblasts -RETIRED-|9982/3
C1264195|T191|OF|56837009|SNOMEDCT_US|Refractory anemia with ringed sideroblasts -RETIRED-|9982/3
C0334679|T191|OAP|189510008|SNOMEDCT_US|Refractory anemia with sideroblasts|9982/3
C0334679|T191|OAP|56837009|SNOMEDCT_US|Refractory anemia with sideroblasts|9982/3
C0334679|T191|SY|109998009|SNOMEDCT_US|Refractory anemia with sideroblasts|9982/3
C0334679|T191|PT|128846006|SNOMEDCT_US|Refractory anemia with sideroblasts|9982/3
C0002894|T191|SY|0000001134|CHV|raeb|9983/3
C0002894|T191|SY|0000001134|CHV|smoldering leukemia|9983/3
C0002894|T191|PT|D46.2|ICD10|Refractory anaemia with excess of blasts|9983/3
C0002894|T191|PT|D46.2|ICD10AE|Refractory anemia with excess of blasts|9983/3
C1318550|T191|ET|D46.21|ICD10CM|RAEB 1|9983/3
C1318551|T191|ET|D46.22|ICD10CM|RAEB 2|9983/3
C0002894|T191|ET|D46.20|ICD10CM|RAEB NOS|9983/3
C1318550|T191|AB|D46.21|ICD10CM|Refractory anemia with excess of blasts 1|9983/3
C1318550|T191|PT|D46.21|ICD10CM|Refractory anemia with excess of blasts 1|9983/3
C1318551|T191|AB|D46.22|ICD10CM|Refractory anemia with excess of blasts 2|9983/3
C1318551|T191|PT|D46.22|ICD10CM|Refractory anemia with excess of blasts 2|9983/3
C0002894|T191|AB|D46.20|ICD10CM|Refractory anemia with excess of blasts, unspecified|9983/3
C0002894|T191|PT|D46.20|ICD10CM|Refractory anemia with excess of blasts, unspecified|9983/3
C0002894|T191|PT|MTHU063670|ICPC2ICD10ENG|RAEB|9983/3
C0002894|T191|LLT|10037803|MDR|RAEB|9983/3
C0002894|T191|LLT|10038270|MDR|Refractory anaemia with an excess of blasts|9983/3
C0002894|T191|PT|10038270|MDR|Refractory anaemia with an excess of blasts|9983/3
C0002894|T191|LLT|10054592|MDR|Refractory anemia with an excess of blasts|9983/3
C0002894|T191|MTH_PT|10038270|MDR|Refractory anemia with an excess of blasts|9983/3
C0002894|T191|SY|35940|MEDCIN|anemia refractory with excess blasts|9983/3
C0002894|T191|PT|35940|MEDCIN|refractory anemia with excess blasts|9983/3
C1318550|T191|PT|311868|MEDCIN|refractory anemia with excess blasts-1|9983/3
C1318551|T191|PT|311869|MEDCIN|refractory anemia with excess blasts-2|9983/3
C0002894|T191|MH|D000754|MSH|Anemia, Refractory, with Excess of Blasts|9983/3
C0002894|T191|ET|D000754|MSH|Leukemia, Smoldering|9983/3
C0002894|T191|ET|D000754|MSH|Leukemia, Smouldering|9983/3
C0002894|T191|PM|D000754|MSH|Leukemias, Smoldering|9983/3
C0002894|T191|ET|D000754|MSH|RAEB|9983/3
C0002894|T191|ET|D000754|MSH|RAEM|9983/3
C0002894|T191|ET|D000754|MSH|Refractory Anemia with Excess of Blasts|9983/3
C0002894|T191|PM|D000754|MSH|Smoldering Leukemia|9983/3
C0002894|T191|PM|D000754|MSH|Smoldering Leukemias|9983/3
C0002894|T191|PM|D000754|MSH|Smouldering Leukemia|9983/3
C0002894|T191|PN|NOCODE|MTH|Refractory anaemia with excess blasts|9983/3
C0002894|T191|AB|C7506|NCI|MDS-EB|9983/3
C1318550|T191|AB|C7167|NCI|MDS-EB-1|9983/3
C1318551|T191|AB|C7168|NCI|MDS-EB-2|9983/3
C0002894|T191|PT|C7506|NCI|Myelodysplastic Syndrome with Excess Blasts|9983/3
C1318550|T191|PT|C7167|NCI|Myelodysplastic Syndrome with Excess Blasts-1|9983/3
C1318551|T191|PT|C7168|NCI|Myelodysplastic Syndrome with Excess Blasts-2|9983/3
C0002894|T191|AB|C7506|NCI|RAEB|9983/3
C1318550|T191|AB|C7167|NCI|RAEB-1|9983/3
C1318551|T191|AB|C7168|NCI|RAEB-2|9983/3
C1318550|T191|AB|C7167|NCI|RAEB-I|9983/3
C1318551|T191|AB|C7168|NCI|RAEB-II|9983/3
C0002894|T191|SY|C7506|NCI|Refractory Anemia with an Excess of Blasts|9983/3
C0002894|T191|SY|C7506|NCI|Refractory Anemia with Excess Blasts|9983/3
C0002894|T191|PT|C7506|NCI_CPTAC|Myelodysplastic Syndrome with Excess Blasts|9983/3
C1318551|T191|PT|C7168|NCI_CPTAC|Myelodysplastic Syndrome with Excess Blasts-2|9983/3
C0002894|T191|DN|C7506|NCI_CTRP|Myelodysplastic Syndrome with Excess Blasts|9983/3
C0002894|T191|PT|CDR0000040359|PDQ|refractory anemia with excess blasts|9983/3
C0002894|T191|SY|Xa0Sf|RCD|RAEB - Refractory anaemia with excess blasts|9983/3
C0002894|T191|IS|B9372|RCD|RAEB - Refractory anaemia with excess of blasts|9983/3
C0002894|T191|OA|B9372|RCD|RAEB-Refrac anaem+exces blasts|9983/3
C0002894|T191|AB|Xa0Sf|RCD|RAEB-Refrac anaem+excess blast|9983/3
C0002894|T191|OA|B9372|RCD|Refr anaem with excess blasts|9983/3
C0002894|T191|AB|Xa0Sf|RCD|Refrac anaem with excess blast|9983/3
C0002894|T191|PT|Xa0Sf|RCD|Refractory anaemia with excess blasts|9983/3
C0002894|T191|OP|B9372|RCD|Refractory anaemia with excess of blasts|9983/3
C0002894|T191|SY|Xa0Sf|RCD|Smouldering leukaemia|9983/3
C0002894|T191|SY|Xa0Sf|RCDAE|RAEB - Refractory anemia with excess blasts|9983/3
C0002894|T191|IS|B9372|RCDAE|RAEB - Refractory anemia with excess of blasts|9983/3
C0002894|T191|PT|Xa0Sf|RCDAE|Refractory anemia with excess blasts|9983/3
C0002894|T191|OP|B9372|RCDAE|Refractory anemia with excess of blasts|9983/3
C0002894|T191|SY|Xa0Sf|RCDAE|Smouldering leukemia|9983/3
C0002894|T191|PT|XaBC5|RCDSA|Refractory anemia with excess of blasts|9983/3
C0002894|T191|AB|XaBC5|RCDSY|Refract anaem+excess blasts|9983/3
C0002894|T191|PT|XaBC5|RCDSY|Refractory anaemia with excess of blasts|9983/3
C0002894|T191|SY|128847002|SNOMEDCT_US|RAEB|9983/3
C0002894|T191|OAS|109999001|SNOMEDCT_US|RAEB - Refractory anaemia with excess blasts|9983/3
C0002894|T191|SYGB|398623004|SNOMEDCT_US|RAEB - Refractory anaemia with excess blasts|9983/3
C0002894|T191|OAS|189511007|SNOMEDCT_US|RAEB - Refractory anaemia with excess of blasts|9983/3
C0002894|T191|OAS|109999001|SNOMEDCT_US|RAEB - Refractory anemia with excess blasts|9983/3
C0002894|T191|SY|398623004|SNOMEDCT_US|RAEB - Refractory anemia with excess blasts|9983/3
C0002894|T191|OAS|189511007|SNOMEDCT_US|RAEB - Refractory anemia with excess of blasts|9983/3
C1318550|T191|IS|128847002|SNOMEDCT_US|RAEB I|9983/3
C1318550|T191|SY|397338009|SNOMEDCT_US|RAEB I|9983/3
C1318551|T191|IS|128847002|SNOMEDCT_US|RAEB II|9983/3
C1318551|T191|SY|397339001|SNOMEDCT_US|RAEB II|9983/3
C0002894|T191|PTGB|128847002|SNOMEDCT_US|Refractory anaemia with excess blasts|9983/3
C0002894|T191|SYGB|398623004|SNOMEDCT_US|Refractory anaemia with excess blasts|9983/3
C1318550|T191|PTGB|397338009|SNOMEDCT_US|Refractory anaemia with excess blasts I|9983/3
C1318551|T191|PTGB|397339001|SNOMEDCT_US|Refractory anaemia with excess blasts II|9983/3
C1318550|T191|PTGB|415283002|SNOMEDCT_US|Refractory anaemia with excess blasts-1|9983/3
C1318551|T191|PTGB|415284008|SNOMEDCT_US|Refractory anaemia with excess blasts-2|9983/3
C0002894|T191|OAP|189511007|SNOMEDCT_US|Refractory anaemia with excess of blasts|9983/3
C0002894|T191|OAP|16956001|SNOMEDCT_US|Refractory anaemia with excess of blasts|9983/3
C0002894|T191|IS|16956001|SNOMEDCT_US|Refractory anaemia with excess of blasts -RETIRED-|9983/3
C0002894|T191|PT|128847002|SNOMEDCT_US|Refractory anemia with excess blasts|9983/3
C0002894|T191|SY|398623004|SNOMEDCT_US|Refractory anemia with excess blasts|9983/3
C1318550|T191|PT|397338009|SNOMEDCT_US|Refractory anemia with excess blasts I|9983/3
C1318551|T191|PT|397339001|SNOMEDCT_US|Refractory anemia with excess blasts II|9983/3
C1318550|T191|PT|415283002|SNOMEDCT_US|Refractory anemia with excess blasts-1|9983/3
C1318551|T191|PT|415284008|SNOMEDCT_US|Refractory anemia with excess blasts-2|9983/3
C0002894|T191|OAP|189511007|SNOMEDCT_US|Refractory anemia with excess of blasts|9983/3
C0002894|T191|OAP|16956001|SNOMEDCT_US|Refractory anemia with excess of blasts|9983/3
C0002894|T191|IS|16956001|SNOMEDCT_US|Refractory anemia with excess of blasts -RETIRED-|9983/3
C0002894|T191|OF|16956001|SNOMEDCT_US|Refractory anemia with excess of blasts -RETIRED-|9983/3
C0280028|T047|PT|D46.3|ICD10|Refractory anaemia with excess of blasts with transformation|9984/3
C0280028|T047|PT|D46.3|ICD10AE|Refractory anemia with excess of blasts with transformation|9984/3
C0280028|T047|LLT|10038271|MDR|Refractory anaemia with excess blasts in transformation|9984/3
C0280028|T047|LLT|10054593|MDR|Refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|AB|C27080|NCI|RAEB-T|9984/3
C0280028|T047|PT|C27080|NCI|Refractory Anemia with Excess Blasts in Transformation|9984/3
C0280028|T047|OP|C27080|NCI|Refractory Anemia with Excess Blasts in Transformation|9984/3
C0280028|T047|DN|C27080|NCI_CTRP|Refractory Anemia with Excess Blasts in Transformation|9984/3
C0280028|T047|PT|CDR0000040360|PDQ|refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|SY|Xa0Sg|RCD|RAEB-T - Refractory anaemia with excess blasts in transformation|9984/3
C0280028|T047|AB|Xa0Sg|RCD|RAEB-T - Refractory anaemia+excess blasts in transformation|9984/3
C0280028|T047|AB|Xa0Sg|RCD|RAEBT-Refr anaem+exc bl trans|9984/3
C0280028|T047|OA|B9373|RCD|Ref anaem+exc blast with trnsf|9984/3
C0280028|T047|AB|Xa0Sg|RCD|Refr anaem+exc blasts in trans|9984/3
C0280028|T047|PT|Xa0Sg|RCD|Refractory anaemia with excess blasts in transformation|9984/3
C0280028|T047|OP|B9373|RCD|Refractory anaemia with excess of blasts with transformation|9984/3
C0280028|T047|SY|Xa0Sg|RCDAE|RAEB-T - Refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|AB|Xa0Sg|RCDAE|RAEB-T - Refractory anemia+excess blasts in transformation|9984/3
C0280028|T047|PT|Xa0Sg|RCDAE|Refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|OP|B9373|RCDAE|Refractory anemia with excess of blasts with transformation|9984/3
C0280028|T047|OP|BBmB.|RCDSA|Refractory anemia with excess of blasts with transformation|9984/3
C0280028|T047|OA|BBmB.|RCDSA|Refractory anemia+excess of blasts with transformation|9984/3
C0280028|T047|OA|BBmB.|RCDSY|Refr anam+xs blst+transform|9984/3
C0280028|T047|OP|BBmB.|RCDSY|Refractory anaemia with excess of blasts with transformation|9984/3
C0280028|T047|OA|BBmB.|RCDSY|Refractory anaemia+excess of blasts with transformation|9984/3
C0280028|T047|SY|128848007|SNOMEDCT_US|RAEB-T|9984/3
C0280028|T047|OAS|277596001|SNOMEDCT_US|RAEB-T - Refractory anaemia with excess blasts in transformation|9984/3
C0280028|T047|SYGB|110000005|SNOMEDCT_US|RAEB-T - Refractory anaemia with excess blasts in transformation|9984/3
C0280028|T047|OAS|277596001|SNOMEDCT_US|RAEB-T - Refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|SY|110000005|SNOMEDCT_US|RAEB-T - Refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|SYGB|110000005|SNOMEDCT_US|Refractory anaemia with excess blasts in transformation|9984/3
C0280028|T047|OAP|277596001|SNOMEDCT_US|Refractory anaemia with excess blasts in transformation|9984/3
C0280028|T047|PTGB|128848007|SNOMEDCT_US|Refractory anaemia with excess blasts in transformation|9984/3
C0280028|T047|OAP|64839007|SNOMEDCT_US|Refractory anaemia with excess of blasts with transformation|9984/3
C0280028|T047|OAP|189512000|SNOMEDCT_US|Refractory anaemia with excess of blasts with transformation|9984/3
C0280028|T047|IS|64839007|SNOMEDCT_US|Refractory anaemia with excess of blasts with transformation -RETIRED-|9984/3
C0280028|T047|SY|110000005|SNOMEDCT_US|Refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|OAP|277596001|SNOMEDCT_US|Refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|PT|128848007|SNOMEDCT_US|Refractory anemia with excess blasts in transformation|9984/3
C0280028|T047|OAP|64839007|SNOMEDCT_US|Refractory anemia with excess of blasts with transformation|9984/3
C0280028|T047|OAP|189512000|SNOMEDCT_US|Refractory anemia with excess of blasts with transformation|9984/3
C0280028|T047|IS|64839007|SNOMEDCT_US|Refractory anemia with excess of blasts with transformation -RETIRED-|9984/3
C0280028|T047|OF|64839007|SNOMEDCT_US|Refractory anemia with excess of blasts with transformation -RETIRED-|9984/3
C0796466|T191|PT|D46.A|ICD10CM|Refractory cytopenia with multilineage dysplasia|9985/3
C0796466|T191|AB|D46.A|ICD10CM|Refractory cytopenia with multilineage dysplasia|9985/3
C0796466|T191|LLT|10067959|MDR|Refractory cytopenia with multilineage dysplasia|9985/3
C0796466|T191|PT|10067959|MDR|Refractory cytopenia with multilineage dysplasia|9985/3
C0796466|T191|PT|230932|MEDCIN|refractory cytopenia with multilineage dysplasia|9985/3
C2826323|T191|PN|NOCODE|MTH|Refractory Cytopenia of Childhood|9985/3
C0796466|T191|AB|C8574|NCI|MDS-MLD|9985/3
C0796466|T191|PT|C8574|NCI|Myelodysplastic Syndrome with Multilineage Dysplasia|9985/3
C2826323|T191|AB|C82596|NCI|RCC|9985/3
C0796466|T191|AB|C8574|NCI|RCMD|9985/3
C2826323|T191|PT|C82596|NCI|Refractory Cytopenia of Childhood|9985/3
C0796466|T191|SY|C8574|NCI|Refractory Cytopenia with Multilineage Dysplasia|9985/3
C0796466|T191|DN|C8574|NCI_CTRP|Myelodysplastic Syndrome with Multilineage Dysplasia|9985/3
C2826323|T191|AB|C82596|NCI_NICHD|RCC|9985/3
C2826323|T191|PT|C82596|NCI_NICHD|Refractory Cytopenia of Childhood|9985/3
C0796466|T191|AB|CDR0000043315|PDQ|RCMD|9985/3
C0796466|T191|PT|CDR0000043315|PDQ|refractory cytopenia with multilineage dysplasia|9985/3
C0796466|T191|PTGB|415285009|SNOMEDCT_US|Refractory cytopaenia with multilineage dysplasia|9985/3
C2826323|T191|SY|128836009|SNOMEDCT_US|Refractory cytopenia of childhood|9985/3
C0796466|T191|PT|415285009|SNOMEDCT_US|Refractory cytopenia with multilineage dysplasia|9985/3
C0796466|T191|PT|128836009|SNOMEDCT_US|Refractory cytopenia with multilineage dysplasia|9985/3
C1292779|T191|ET|D46.C|ICD10CM|5q minus syndrome NOS|9986/3
C1292779|T191|ET|D46.C|ICD10CM|Myelodysplastic syndrome with 5q deletion|9986/3
C1292779|T191|PT|238.74|ICD9CM|Myelodysplastic syndrome with 5q deletion|9986/3
C1292779|T191|AB|238.74|ICD9CM|Myelodyspls syn w 5q del|9986/3
C1292779|T191|PT|230933|MEDCIN|myelodysplastic syndrome with 5q deletion syndrome|9986/3
C1292779|T191|ET|238.74|MTHICD9|5q minus syndrome NOS|9986/3
C1292779|T191|SY|C6867|NCI|5q- Syndrome|9986/3
C1292779|T191|SY|C6867|NCI|Myelodysplastic Syndrome with 5q Deletion|9986/3
C1292779|T191|PT|CDR0000531047|NCI_NCI-GLOSS|5Q minus syndrome|9986/3
C1292779|T191|PT|CDR0000044810|NCI_NCI-GLOSS|5Q- syndrome|9986/3
C1292779|T191|PT|Xa0Sh|RCD|5Q minus syndrome|9986/3
C1292779|T191|IS|277597005|SNOMEDCT_US|5Q minus syndrome|9986/3
C1292779|T191|SY|277597005|SNOMEDCT_US|5q minus syndrome|9986/3
C1292779|T191|SY|277597005|SNOMEDCT_US|Myelodysplastic syndrome with 5Q deletion|9986/3
C1292779|T191|IS|128837000|SNOMEDCT_US|Myelodysplastic syndrome with 5q- syndrome|9986/3
C1292779|T191|PT|128837000|SNOMEDCT_US|Myelodysplastic syndrome with 5q- syndrome|9986/3
C1292780|T191|PT|230934|MEDCIN|therapy-related myelodysplastic syndrome|9987/3
C1292780|T191|AB|C27722|NCI|t-MDS|9987/3
C1292780|T191|SY|C27722|NCI|Therapy Related Myelodysplastic Syndrome|9987/3
C1292780|T191|SY|C27722|NCI|Therapy-Related MDS|9987/3
C1292780|T191|PT|C27722|NCI|Therapy-Related Myelodysplastic Syndrome|9987/3
C1292780|T191|PT|702476004|SNOMEDCT_US|Therapy-related myelodysplastic syndrome|9987/3
C1292780|T191|PT|128838005|SNOMEDCT_US|Therapy-related myelodysplastic syndrome|9987/3
C1292780|T191|SY|128838005|SNOMEDCT_US|Therapy-related myelodysplastic syndrome, alkylating agent related|9987/3
C1292780|T191|SY|128838005|SNOMEDCT_US|Therapy-related myelodysplastic syndrome, epidopophyllotoxin-related|9987/3
C3463824|T191|PT|0045936|CCPSS|MYELODYSPLASTIC SYNDROME|9989/3
C3463824|T191|SY|0000010081|CHV|myelodysplasia|9989/3
C3463824|T191|PT|0000008407|CHV|myelodysplasia|9989/3
C3463824|T191|SY|0000010081|CHV|myelodysplastic syndrome|9989/3
C3463824|T191|SY|0000008407|CHV|myelodysplastic syndrome|9989/3
C3463824|T191|SY|0000008407|CHV|myelodysplastic syndromes|9989/3
C3463824|T191|SY|0000010081|CHV|myeloid dysplasia|9989/3
C3463824|T191|PT|0000010081|CHV|preleukemia|9989/3
C3463824|T191|PT|U000455|COSTAR|MYELODYSPLASTIC SYNDROME|9989/3
C3463824|T191|DI|U001579|DXP|PRELEUKEMIC SYNDROME|9989/3
C3463824|T191|PT|HP:0002863|HPO|Myelodysplasia|9989/3
C3463824|T191|SY|HP:0002863|HPO|Myelodysplastic syndrome|9989/3
C3463824|T191|PT|D46.9|ICD10|Myelodysplastic syndrome, unspecified|9989/3
C3463824|T191|HT|D46|ICD10|Myelodysplastic syndromes|9989/3
C3463824|T191|PT|D46.9|ICD10CM|Myelodysplastic syndrome, unspecified|9989/3
C3463824|T191|AB|D46.9|ICD10CM|Myelodysplastic syndrome, unspecified|9989/3
C3463824|T191|AB|D46|ICD10CM|Myelodysplastic syndromes|9989/3
C3463824|T191|HT|D46|ICD10CM|Myelodysplastic syndromes|9989/3
C3463824|T191|AB|238.75|ICD9CM|Myelodysplastic synd NOS|9989/3
C3463824|T191|PT|238.75|ICD9CM|Myelodysplastic syndrome, unspecified|9989/3
C3463824|T191|PT|MTHU050844|ICPC2ICD10ENG|myelodysplasia|9989/3
C3463824|T191|PT|MTHU050847|ICPC2ICD10ENG|myelodysplastic; syndrome|9989/3
C3463824|T191|PT|MTHU061498|ICPC2ICD10ENG|preleukemia|9989/3
C3463824|T191|PT|MTHU061499|ICPC2ICD10ENG|preleukemic; syndrome|9989/3
C3463824|T191|PT|MTHU072863|ICPC2ICD10ENG|syndrome; myelodysplastic|9989/3
C3463824|T191|PT|MTHU072947|ICPC2ICD10ENG|syndrome; preleukemic|9989/3
C3463824|T191|PT|B75008|ICPC2P|Myelodysplastic Syndrome|9989/3
C3463824|T191|PTN|B75008|ICPC2P|myelodysplastic syndrome|9989/3
C3463824|T191|PT|U003813|LCH|Preleukemia|9989/3
C3463824|T191|PT|sh88001636|LCH_NW|Myelodysplastic syndromes|9989/3
C3463824|T191|PT|sh85106315|LCH_NW|Preleukemia|9989/3
C3463824|T191|LA|LA26796-5|LNC|Myelodysplastic syndrome|9989/3
C3463824|T191|LLT|10028533|MDR|Myelodysplastic syndrome|9989/3
C3463824|T191|PT|10028533|MDR|Myelodysplastic syndrome|9989/3
C3463824|T191|LLT|10028534|MDR|Myelodysplastic syndrome NOS|9989/3
C1268964|T191|LLT|10028535|MDR|Myelodysplastic syndrome unclassifiable|9989/3
C1268964|T191|PT|10028535|MDR|Myelodysplastic syndrome unclassifiable|9989/3
C3463824|T191|HT|10028536|MDR|Myelodysplastic syndromes|9989/3
C3463824|T191|LLT|10028548|MDR|Myeloid dysplasia|9989/3
C3463824|T191|LLT|10036587|MDR|Preleukaemia|9989/3
C3463824|T191|LLT|10054577|MDR|Preleukemia|9989/3
C3463824|T191|PT|98952|MEDCIN|myelodysplasia|9989/3
C3463824|T191|PT|35938|MEDCIN|myelodysplastic syndrome|9989/3
C3463824|T191|ET|5550|MEDLINEPLUS|MDS|9989/3
C3463824|T191|SY|5550|MEDLINEPLUS|MDS|9989/3
C3463824|T191|PT|5550|MEDLINEPLUS|Myelodysplastic Syndromes|9989/3
C3463824|T191|PM|D009190|MSH|Dysmyelopoietic Syndrome|9989/3
C3463824|T191|ET|D009190|MSH|Dysmyelopoietic Syndromes|9989/3
C3463824|T191|PM|D009190|MSH|Myelodysplastic Syndrome|9989/3
C3463824|T191|MH|D009190|MSH|Myelodysplastic Syndromes|9989/3
C3463824|T191|PM|D009190|MSH|Syndrome, Dysmyelopoietic|9989/3
C3463824|T191|PM|D009190|MSH|Syndrome, Myelodysplastic|9989/3
C3463824|T191|PM|D009190|MSH|Syndromes, Dysmyelopoietic|9989/3
C3463824|T191|PM|D009190|MSH|Syndromes, Myelodysplastic|9989/3
C3463824|T191|PN|NOCODE|MTH|MYELODYSPLASTIC SYNDROME|9989/3
C3463824|T191|SY|C3247|NCI|Dysmyelopoietic Syndrome|9989/3
C3463824|T191|AB|C3247|NCI|MDS|9989/3
C1268964|T191|AB|C8648|NCI|MDS-U|9989/3
C1268964|T191|AB|C8648|NCI|MDS, U|9989/3
C3463824|T191|SY|C3247|NCI|Myelodysplasia|9989/3
C3463824|T191|SY|C3247|NCI|Myelodysplastic Neoplasm|9989/3
C3463824|T191|SY|TCGA|NCI|Myelodysplastic Syndrome|9989/3
C3463824|T191|PT|C3247|NCI|Myelodysplastic Syndrome|9989/3
C1268964|T191|PT|C8648|NCI|Myelodysplastic Syndrome, Unclassifiable|9989/3
C1268964|T191|SY|TCGA|NCI|Myelodysplastic Syndrome, Unclassifiable|9989/3
C3463824|T191|SY|C3247|NCI|Myelodysplastic Syndrome/Neoplasm|9989/3
C3463824|T191|SY|C3247|NCI|Oligoblastic Leukemia|9989/3
C3463824|T191|OP|C3247|NCI|Preleukemia|9989/3
C3463824|T191|SY|C3247|NCI|Smoldering Leukemia|9989/3
C1268964|T191|SY|C8648|NCI|Unclassifiable MDS|9989/3
C1268964|T191|SY|C8648|NCI|Unclassifiable Myelodysplastic Syndrome|9989/3
C3463824|T191|PT|C3247|NCI_CPTAC|Myelodysplastic Syndrome|9989/3
C3463824|T191|PT|E12552|NCI_CTCAE|Myelodysplastic syndrome|9989/3
C3463824|T191|PT|10028534|NCI_CTEP-SDC|Myelodysplastic syndrome, NOS|9989/3
C3463824|T191|DN|C3247|NCI_CTRP|Myelodysplastic Syndrome|9989/3
C3463824|T191|PT|C3247|NCI_CTRP|Myelodysplastic Syndrome|9989/3
C3463824|T191|PT|CDR0000045953|NCI_NCI-GLOSS|myelodysplasia|9989/3
C3463824|T191|PT|CDR0000045266|NCI_NCI-GLOSS|myelodysplastic syndromes|9989/3
C3463824|T191|PT|CDR0000045480|NCI_NCI-GLOSS|preleukemia|9989/3
C3463824|T191|PT|CDR0000046583|NCI_NCI-GLOSS|smoldering leukemia|9989/3
C3463824|T191|PT|C3247|NCI_NICHD|Myelodysplastic Syndrome|9989/3
C3463824|T191|SY|CDR0000039817|PDQ|dysmyelopoiesis|9989/3
C3463824|T191|SY|CDR0000039817|PDQ|Dysmyelopoietic Syndrome|9989/3
C3463824|T191|AB|CDR0000039817|PDQ|MDS|9989/3
C3463824|T191|SY|CDR0000039817|PDQ|myelodysplasia|9989/3
C3463824|T191|SY|CDR0000039817|PDQ|Myelodysplastic Syndrome|9989/3
C3463824|T191|PT|CDR0000039817|PDQ|myelodysplastic syndromes|9989/3
C3463824|T191|ET|CDR0000039817|PDQ|Myelodysplastic syndromes|9989/3
C3463824|T191|SY|CDR0000039817|PDQ|Oligoblastic Leukemia|9989/3
C3463824|T191|SY|CDR0000039817|PDQ|preleukemia|9989/3
C3463824|T191|SY|CDR0000039817|PDQ|Smoldering Leukemia|9989/3
C3463824|T191|SY|Xa0SY|RCD|MDS - Myelodysplastic syndrome|9989/3
C3463824|T191|SY|Xa0SY|RCD|Myelodysplasia|9989/3
C3463824|T191|PT|Xa0SY|RCD|Myelodysplastic syndrome|9989/3
C3463824|T191|OA|ByuHD|RCDSY|Myelodysplastic synd,unspec|9989/3
C3463824|T191|OP|BBv..|RCDSY|Myelodysplastic syndrome|9989/3
C3463824|T191|OP|ByuHD|RCDSY|Myelodysplastic syndrome, unspecified|9989/3
C3463824|T191|OAS|4227006|SNOMEDCT_US|Dysmyelopoietic syndrome|9989/3
C3463824|T191|SY|128623006|SNOMEDCT_US|Dysmyelopoietic syndrome|9989/3
C3463824|T191|SY|109995007|SNOMEDCT_US|MDS - Myelodysplastic syndrome|9989/3
C3463824|T191|OAS|189508006|SNOMEDCT_US|Myelodysplasia|9989/3
C3463824|T191|OAS|189515003|SNOMEDCT_US|Myelodysplasia|9989/3
C3463824|T191|OF|25707000|SNOMEDCT_US|Myelodysplasia|9989/3
C3463824|T191|OAP|25707000|SNOMEDCT_US|Myelodysplasia|9989/3
C3463824|T191|SY|109995007|SNOMEDCT_US|Myelodysplastic syndrome|9989/3
C3463824|T191|OAP|393565000|SNOMEDCT_US|Myelodysplastic syndrome|9989/3
C3463824|T191|PT|128623006|SNOMEDCT_US|Myelodysplastic syndrome|9989/3
C3463824|T191|OAS|4227006|SNOMEDCT_US|Myelodysplastic syndrome|9989/3
C3463824|T191|OF|393565000|SNOMEDCT_US|Myelodysplastic syndrome|9989/3
C1268964|T191|PT|373381004|SNOMEDCT_US|Myelodysplastic syndrome, no ICD-O subtype|9989/3
C1268964|T191|SY|373381004|SNOMEDCT_US|Myelodysplastic syndrome, no International Classification of Diseases for Oncology subtype|9989/3
C3463824|T191|IS|4227006|SNOMEDCT_US|Myelodysplastic syndrome, NOS|9989/3
C1268964|T191|SY|373381004|SNOMEDCT_US|Myelodysplastic syndrome, unclassifiable|9989/3
C3463824|T191|OAS|189515003|SNOMEDCT_US|Myelodysplastic syndrome, unspecified|9989/3
C3463824|T191|IS|128623006|SNOMEDCT_US|Preleukaemia|9989/3
C3463824|T191|OAS|4227006|SNOMEDCT_US|Preleukaemia|9989/3
C3463824|T191|OAS|4227006|SNOMEDCT_US|Preleukaemic syndrome|9989/3
C3463824|T191|IS|128623006|SNOMEDCT_US|Preleukaemic syndrome|9989/3
C3463824|T191|IS|128623006|SNOMEDCT_US|Preleukemia|9989/3
C3463824|T191|OAS|4227006|SNOMEDCT_US|Preleukemia|9989/3
C3463824|T191|IS|128623006|SNOMEDCT_US|Preleukemic syndrome|9989/3
C3463824|T191|OAS|4227006|SNOMEDCT_US|Preleukemic syndrome|9989/3
C3463824|T191|SY|188736006|SNOMEDCT_US|Smoldering leukemia|9989/3
C3463824|T191|OAS|109999001|SNOMEDCT_US|Smoldering leukemia|9989/3
C3463824|T191|OAS|109999001|SNOMEDCT_US|Smouldering leukaemia|9989/3
C3463824|T191|SYGB|188736006|SNOMEDCT_US|Smouldering leukaemia|9989/3
C3463824|T191|IT|0565|WHO|MYELODYSPLASTIC SYNDROME|9989/3
C3463824|T191|PT|1498|WHO|MYELOID DYSPLASIA|9989/3
C2826320|T191|SY|366674|MEDCIN|neutropenia refractory|9991/3
C2826320|T191|PT|366674|MEDCIN|Refractory neutropenia|9991/3
C2826320|T191|PN|NOCODE|MTH|Refractory Neutropenia|9991/3
C2826320|T191|PT|C82593|NCI|Refractory Neutropenia|9991/3
C2826320|T191|AB|C82593|NCI|RN|9991/3
C2826320|T191|PTGB|721303001|SNOMEDCT_US|Refractory neutropaenia|9991/3
C2826320|T191|PTGB|450946009|SNOMEDCT_US|Refractory neutropaenia|9991/3
C2826320|T191|PT|450946009|SNOMEDCT_US|Refractory neutropenia|9991/3
C2826320|T191|PT|721303001|SNOMEDCT_US|Refractory neutropenia|9991/3
C2826321|T191|PT|366675|MEDCIN|Refractory thrombocytopenia|9992/3
C2826321|T191|SY|366675|MEDCIN|thrombocytopenia refractory|9992/3
C2826321|T191|PN|NOCODE|MTH|Refractory Thrombocytopenia|9992/3
C2826321|T191|PT|C82594|NCI|Refractory Thrombocytopenia|9992/3
C2826321|T191|AB|C82594|NCI|RT|9992/3
C2826321|T191|PTGB|721304007|SNOMEDCT_US|Refractory thrombocytopaenia|9992/3
C2826321|T191|PTGB|450947000|SNOMEDCT_US|Refractory thrombocytopaenia|9992/3
C2826321|T191|PT|721304007|SNOMEDCT_US|Refractory thrombocytopenia|9992/3
C2826321|T191|PT|450947000|SNOMEDCT_US|Refractory thrombocytopenia|9992/3
C0555198|T191|PM|D005910|MSH|Glioma|9380/3
C0262584|T191|SY|Xa989|RCD|SCC|9380/3
C1266002|T191|SY|0000056675|CHV|NSCLC|8046/3
C1266002|T191|SY|0000056675|CHV|non-small-cell carcinoma|8046/3
C1266002|T191|SY|0000056675|CHV|nonsmall cell carcinoma|8046/3
C1266002|T191|SY|0000056675|CHV|nonsmall-cell carcinoma|8046/3
C0334247|T191|SY|TCGA|NCI|Keratinizing Squamous Carcinoma|8071/3
C1266005|T191|SY|TCGA|NCI|squamous cell carcinoma, basaloid type|8083/3
C0206692|T191|SY|0000021024|CHV|infiltrating mammary carcinoma with lobular|8520/3
